// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ItApMrz7cFd1AZrsw2H6lwRbpaFwwD8lfByFWS/FvK9AUMIrrwrO6yVtcKfcApLp
0TjSHoW0O/X2w3D2JkSSt4QuARVVshku5c7eLoy3HrO83ZfVqWvrDYwQG0X/oMqT
uLyATszaFxBo7Z1l/lq67WmaYD7CYpntUHki3bBUGZw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12064)
K4sSgGgFttQ9GKNiCAC3Qpz/LR/jGKDFYXHvGwWB3odn2XxS+NDtdIUCDNpnBTOY
CjQCzOCn8W1dWkRwFFEtBjrqW7eEqwAgdQ1hxM4phqYjMb2nTYLnSrxOYokyfRph
QZHTfE104yBrovIBlxFSJuZkTLG0F6/PT6zis67n5/C6zD6tSmXYF+1q1d6wQ8dG
7PU+xOaJmZHc7RxpHGL4yt4GirmS3TJs5RRGCler/rZ72k0N87UF62qpjKIRiU7g
gyjLtXsLKOvWyxusSdWWK1W+1ffOPRVH1b6mdcP71MS8elS6DYbYOwPWz7Oh6XSB
gEDcgivd5XPKr3GSHWegBL6kg0L22sBuAofFlDbAM/S4GSAEpzq75O/eXAhn4/ca
PyrA2oFD53Ik6i4aj7pNLG/uKWm5sIw1I/QLuGcS1gU9ThqrKfNCYkPBu8LMwiEy
Yf0G5G3NF0kxrT/UjH9C6sL1kk4aaclqLnM2hHNksrv2+CxCDZGV6bwg5m4CwmEs
NIVCjrHgc0IiXveY1z5gAYLbwtCa6yZiFsdSAYPXI289dYP7Gw4YJ+3oSFjO4Qw6
8o4mZH6+Fs0kQ1/iZurhr9fcLLF9joSIdOapIkUfipCxmd9OzxBgNTlxrfoDd+EM
P6i1Z9+7nePr2h1gduAz5JWH7lQPypJmF+uyM4ui02Gm3oZqQFCLH6I7ALld5ngM
foYfCIlc27bmgXN2F2DPjVbTbw1Wsn0XxbWpyfxlSxz8FXDkOT8Qna8To4h2AWgP
t97pr1Pxo9yD+OWlbFPRyHfGU1jOgM5gBBZDNqqoR9VxkBb+U46l5gEIqs+3zkrk
T56BafEDZuZB3aJUHMtHLS/dULClRQlS1VW1cVDj3dK7m2uwrdMgNT4ymrVu5p+z
WStF3UQDOMcLS4MbrMnecO7Z9aKHhYxEQbzr8w7O1FLWjno6bepvwCpHi42mnS4+
XT0RtW35t2FW6o6rf8tCtxOvunMOMg10+T5/uAQhLt+Ozfie7pskpnZLO6NfUQb7
Kz1KLZBKwAPjtue0ymOlDY/kKu32wuahSykUhuXH5BrpNtfFNy/yWeDg/QDGvU3e
AnJ8Hf8WY0uc8iIvjzQ2OFVF7zQGSUIpKviV5reUXZPa6Iy0NPrDEuPLlJhQV/8E
fVSsQR7TZ5guxPMizJeR/owErshVNSQDjLL0WrNHIOcBfhYvVWtmjzet9YcMuYm7
zQ+RfZuH5pq+ACCJyaCk52vVdg51C2X2kiQQB8IZdfnoh1Eg6XHpjxWDWL5NHsZn
6zkE2OTnSgPMjbiIshOGzs3aNqV8Qi7UamxHg4gSVlaMw/ZELs6gl47bSNHjsTfF
TXiTe1+pGkBPh0Ky5Q2Otvteun9r6IUnd4+yqG+k5L+vFydn59/R1UVzhlIwc8+Q
BJ3raJ2VVxjgNX1Hz2KOwADhqA6pEnalok16H6vgAF1jBr/+08OjHxjCibc2uK0W
+SRFqCwDarfi3KpaFmIJkW1VJEAoTwKmq7i9t9ThoK8Togv6bw9U0ojVyaOnqWs/
lZd6Iccfmnvnh6E5E4Ft7p6tfeaTZ4Z/PfFxShrCYDTThEr468+yiTUyvHMAFNF6
8BmMY7hspFjq/3uy72DHR8bxsxhY9ThVPZjyAdLJmek7xOsh1lUis1I6NFxTIDfQ
rfnxagiE8SIK2uW/eMvHdXVOn3UHClFjb61oO4LBhqkcUAHirj9soJKI90qcpMRs
sv5C+4o+MqP1/UM+I/l9gRQOtSzuRw/7bLFrcG+dXPMOk0HsxvVP1z+HLxdtkma5
wRE8mCGH3v0U6tRaidov6asWkYcsWR1h7SSKg1L/Yr7UYN5mjX3uukB2rDVfP5YY
qX2KIbfsOQRQcDxqE5I8sS3YhQuE/lV95zRCFKYMzM+/Q7PY9Bjie76a1nZ2yVaA
FIsXgU7fza9pEIEqeLFtPuCtg6Mf+uk2APilMsu1gJtERZT5R9YNE5XTkAUInKB0
WNhwt97pNTzUVFuUX6OimUF1UNCHiyGYcu+l2x2WUToRcL1VWfYxEll4wlCH8/BX
WscpzR4pxB0kR60sx6hw9lPt+5nW8griFyPnwUcCqdcdh0hoQdWxTjV2Qk8rLibx
hvgLgMQHEGs7xJ2lZDmaK0bRMVJuhKK1r/+jaQC9ei25vGbFIhSexggYZW9P6kO5
9YLTf25H0KeVhUFVbncJLlNNs6c11L+52XTj55c1edU9HnIB/mCtcazZcpjtAIEU
V7iYvFT8Mu/In5QILZXx08BJwZZILxkROBkHchPHn/LOuMXTY11DCMKWHSUq3caF
+rRVjCiEhaQ7tE+DV86MaKrh30mQVzKNlAvCd2qgMA+z5ik9Vqc/Q2sG33efYZyX
3KnMVHh9X9Oz29iET6t7g1NkOYqLalAZC+45dJj0tg/v3QrtKaimM3w0LqUIBf3Z
SbnktIvX6CULXEjwH13Gi6Py3lbqSy8aLV3in9R9LmhrS87kTXpbUsQvQg67nkTL
rneiXdgzaoRBAKSbRXWOOfAxRYzkuszDfzP6FXFhPfhn5STdR5wwNl57PA8lxtvb
3in/meuFTkF9qUCsdWZ8tDjYA/O/uZp6k337KhSimY0AHCCI0YRgNM3w36lvjlgI
1KljpVbNaBmRVVcwdYvAdkFiJkhbPUEja50VZ+oIFoWA+ecoDoLNkjGo+YCFlMZ4
gJVdjnXXseTqvx0Mh6nTzE4bhutjpOBQAgJyYQnyqyP4doCWk3OEtZSdRTNH8n7k
PAD3hjWEizWv1rRcRI2BpCgiys9BHLUD00SefsFQcsCBn8xvn36DFuI4mzxxQmDv
knQo03D8u4DdJDcFnthHe5wi+BsDgMRQ0j/1wOL7C8p5bnnN0zNpAFqAlsAeKsXa
cnIuZVroUY31ml/t7AshX3upxf2VYazaGlG8PN9MIYg2DertkCAyPU+9mU6OqNqJ
6FArxB8r2SxKzmZAcC6Aygiy1ReY3ETPzx37k/bIyGXR0wkCz1Zh1auJ9RA7C6o3
/fTF4KOcObRTVo2RwSeONZSXMHoPs7hCP7P+/ALMGKy6sMasb+MHWbJHvqT9Zfdk
/lRgMJVfcnUtac2Ss9cwFq8lFoWF963ZrRyvNvHi8DtfLYCxEbOUqd6o4z9OyxfZ
cOUgvMZ5ghVCR8piJ0RzJSKFBO+oOXXgv+YN/Z9gc3bPXo7V68jKY1o9COzKWYZy
5cJQk1uxy74gMTBT59c3Jt5eb7dnjPIT8MS52xKtKJM1qXHVDX/srjeF+SSbdXNY
+V/6YDekevstZoRq214yVHsMhQG7XWSMddXm+hOYwhbs0lwWFlJESB5hzhEJksx/
nSoaXjmL6agE/6QNC/eVBtXUU8De9OhWayU4/vun0sXwaPKsackEj4PWgRY1KsIT
dRuwjfQPv4tOYEItkBDoylvZMqdP+Le3rsea7sMHdTKHEqSh86KFnZp7c6RA0u06
9yaSMVNecl7iTl5+fvdjr/UqwR74W874BEm2sX/VwS/Ik9utmSfqvKhkBfFu/LIH
14/p8iZ6WVinbm85PjHyIPX3B9jEPihEMrIsHKg8+kMVaJDm9a0wacaSxEf27TTK
1Cy/8v9OtCY7evpqbD3LifyPZdNa36Q6/OIXsXRW5dmbrxIXgzeYE2FpQD1jnqgr
/mV/SUu11maNj5lIlc1TJxqwy64Pzmjk5I5sMhe9pHCxZf8IDrnrUyn8qegKO1T7
5lAABN6dlLLGg2NceNRb+PQGsjTiX9OnypU4ioh/IbKu2SUErtu965Jv689ejzFH
ysL+2tGQEkzPnqYH7kF3FqnBopD6Y07ed+cJoSrPOi1A/lm/pxhCO/Nl0wVdKUuV
zAXWR3lmKx4VcPaIWaYL21wlp+sefq7KxbokcrLgRB9dhs8J7pudz2R6Uj9zU0dK
w0cuvT5tl29P1J6wyCZaiyzupYWIexCxCae+tVpaVXRd2jbLqx8MoZ6G9vBjBWwb
3ISotKm3JxaEjutUdqVT7q+iqgXnTFdhvGj1sSEbWAABWzv7g050+5cN3GasUl+7
2vwtCiS0tq++81u7yIbRQZwYtTj9uuBaa7Q69lms9ewP8BJo3c20dWusM04FoItc
e47rTV4zJHjQME/CRelmKGr/0zxlxRArb+fqpBNcbv2s4xershGmcaLO1W6iOdKD
ftBpABpXltF6jYfsS/xGKp70gyKowSK44sE+n5QBm7KFIl+TDkpAfDShjwql7gHJ
rLvZmJ+GTkT3rB0cOXUuTjhH8SrvjVrzg3XEYnLO4oyfQgC0Tf6q0AxfX68rdvqY
MAMxMLAiyIF73USfCJV7YQKWkOVdIKkHui0Y+4OOsd1mz05Z0WGabGgUVme5iQ6i
S9/DzW9XvwNZwRUFn/+74ejuENeN6QVLvAp4/5ZhYljvk6+VvdHVMUBVZxQJtIAK
ehU9G3vYq9qt3ZRLlVWFxcOa6c1LZxb/3a17jPq/XEuEM+V16rxBmbLWrPLmgEmY
SS9KlCU5HT+WN/pysEuaJXJ5zmhaLZ3fDHNDIZyOEFvoKZ0Rdt85hvfynZO4QppF
NlKupef6c8l3ogeNbLVNGkcnWX/oXur0kyhXvhVnHqoDj0M+oP/6svImzROISkN9
keSlJDS5p/Z17LvbrKh2JuaL73cPfEunN+/DCnbArXCYeJC6WVkxf5K6V6/9kqLT
6p8FuUUe9EIX87UoJr3frp3wwcN1mwE2ieU/K/v8Vd2YSLSuaogJm7fE8nM2J2ZC
2RqLAvd/VYDf1KI7UEZhbl1DePRtCFH7tDIsJzLFxyemKP7sQl0qlv9s1XF5wNBA
BTTOKaH2/VbD4abe2UpdIq4xTJAXaoqbbzyLw4iL6TM/r1q3jQ9WS6vyOAgp9ztB
F2TG3ArBSbmttky9U3TTnRXcmNrcTudNPJfM0nAqipihRD/m5qgMldfm830fupoS
vZoxPe+1/2BAsY7xlDL5R7JWhOBzNHTPz50Ni7fe4p0qAi0c88XOzoMh1VZ3atwz
uvo9SwvCdF50M6ZohqHd/gUhRVgmEQ1ImusiQ4oe3yMdTb1f7AdkPGxV9xJOyluB
HoHRKdq+k+bYRIifULvW6FWuOOEPenm4Ct+NJSOi0aivwwF6AdZqSGGguy7HGnZx
WBnYaOB+G2xdBmAlmgZa381jTPuNnpajTdi1zO9+o2ERQJBjelykpn21axf32+pd
ZaPKdAdD0OaUfYmp30vfXyKnSCwKIZWYKb+zBohZwMhLZQHInF1HlPxP+pfBRnTA
TPyvkhgtKicvI/1uJScZfgKhnzgGvWEiRRVsxrWnAhIxl0TTmxPX+eDNjt1K11jE
R+aef0a8zMgZPAZXX6zUnh26RCvB0KfpkDK8MSDYb916AgvWnwfAl5Vldc4Z7trC
Zhemb0NPIEmQiZnGQqXdnbxff6PdiLCkDrFBPc7UKl2B/L6i+qvuIrSIVGi9gX1j
O43FQLu171Ua6sfhdVGvLf4O/K+OeJBI+Jo4a1pXi2eTbZfR6a10NHQuanwd0Poq
P33VkD8efkJCQuhZEvt2KnuL6852qnquTpr0UkKPfrT+xW990Fnd+Ta9FB/zQBhD
v89WzpPDi9E62/IFriOc4OXCxwm6C1NCk8BiQx2l1YG1NaQkiM35kN2LswwQbUM/
S41ruEz1sRocHfGFu43nV3C/uwoL5pC0OzxlupqrsbncJgSMBT2vDV58odYNW20r
lPWzFBJfuOgiCCxP7yV/ml3EYW2E++2JGBUo+V5NLUbRWyNHdCYT4ayJH32Skfqt
wbf9gCFokhXtdnYt2vzbpNk/8UtHjCca5tMCrkcl9K5/adnGfBiKZsgina+rfQ/P
u73yKMiRs4agCkSV45EjR8cOdlcUYARG1SEqb3bm9iFj8FXcabxj5cnNk1MjF5IQ
Z8XZSD1p2a+g953SGmoOiEHpJ4cfriLEwmss85snA7SphKhMloLkVwVxYOf4du9t
gz9XOUXW07dguP3fgIGG97BQEZPIgCIfnR05wzuoYrb0G5oxzBEN/0A2Lax3Z+fL
rlHf6i2st8whXMHtURr0JES14wvz2IEqyP0HISmgwwJQxUOehI94dHRMfDXOsAWK
kNbdLMGRgxBHnXIoNLMxklqctjKXxjpSeLeyUDYMDTpiesHlEI5Zlh9fNZ3XLIYp
e7p6dYnVZs1Ibwq1MYhY3EjTAW0P+h+rf4l9OaoHWCQwp4WwCS5jXtfBCbjSecnz
dlItmQQs7AcYGj4krgZJNu+0mDon4vAzrdugEYjJheNPIs6LBlqxhXlflxejrRcM
dfj4x10B9Y3OuloWLebmNfPNdcvVA81H8QXE1w789IygM/K0vfU1SnsK/3Vnea+C
fFmadh7TvDDaN5aaCAFWXLG2UR9IZMhQqvW7M/nNSJMwbHXws3gEb0vT81AT9Y6E
PqdQ6StiD73gX4Igt5A6/Y3m0yHvgYlvAjXy2Dpz9NG6ed+ZFUknnTdOSxXAVcCM
B21sH/UWWupSAX1KYTDx7KHsKcKDxRwineaj1qonZDX2T3WA582hHGZbneihKNxW
hb779xnTN/iaXBDALHDSgQ6VIrZh6pzpFJc9g4yqi/FZsgDsR3ql/l1+Q/bDH2Q+
hBS5ZOxPpmzPXzZj44Sst7uZMZaAhHPg2lHNPeMXkUPFndYDmVwP/U8FqI5YY8Vz
pEcweWd2A7I61l32OiVEib8MAPSEKfiv4HvVVj/9haFNTqeF4fuCYCsq1+WDlnmz
mHeRpB17kl2ueku66vr9dINkzLeTmGYa/MlfKZP3p70PzPO2ESFYlxwJtl6C84+X
e61+7NG0GCdDasykxqUTPNg8ynN/dc+CEnhzALY4zWf0O3nkxR5dkfPQLXVOE2Ju
nPz3anihPKBuZsPQHevdOEWgJHONEH+erEpSSwzAyNz7e1CMknamWxrcpqcyVz1P
93tKTAT3IixThL88ZWzRIfxB9ZTUe02Kvj0BGsHQ0oHKoWJ3yxHgZ8y2pFhvS1nY
451udPH5Rz9n5l1amIiiHuNLE/lVWKroCJ8/7KSxRC1HMv/l6pxu1zXeDIkFUlqD
VtCfWqhaRX9vqrHyB6I2pcJb4uSQYpogKgGXyzRo5dQsDcEi/X6pGj16D/FJuXIN
e3mr1c9S1bI5eOdRafIV2iHtU8HoXy6G8m792j4o5Vid0VA/7bCjfQiazlhxf40h
1p2adMgNGBj0DtlIZgY1kyOSM1I2PIe/1cpz3i8Fzm8yba/D8zn8dLbaUqbj9ZHg
AqVPQHtWsEEEQdjWXRGhPIpvi2HLfV+Lo1OaeFxGVvBorL8VLs8zAh30ZxEw7PMs
Pcwi0sHQAo3vD6WJFatiVTeKSaPA31VEJprznRaCViM4ZxfxwDCBTNFwcLH+JcUE
PeFEFWO68xifRj0PkQp3XX5hbigmvxjzLOhLIhzcLXolXm7MySwIMHkTfqY77d+z
NsBZrMCNONMheq53bNVslq9IOqa57cG1MbyM4AcEyAAWOQbuSfsJR+vOJ5AdIQjR
Iy3VqoVnh00d5rVeBAgLm9se8WUI/KWbb8nZSv6EgFxUOTUcC7Y7uCbh2+efIldB
lC0fXzBNWnnx2Sq44b/aZyMxUmPl4ELyR/KbWYO7QkTq4JYFZS8cpVIQZIr29RRR
TaFqbkpOi7YBCxtODFqvjKyoo23HhiFnGKFtjxrTI1NYSOmT1iZuIo/h+FRXSqTA
1qud2dq04uleF4/ZXNKa62hcQSEUt2BNGVevbnn34Y2OYT8wE8wqMY0FQOK2VzJC
PTkjDkmCvhWMYQSiqLMQTAPF73oIxTqsyTTSBfIuWew9abcHsR5uRH60dwzqx3rI
Vupm1QAIsTmy3+Lz2lTc51cHowqWJL+et4yCsvanrPxJHWjBwmHYV6cPgDyDsiLQ
9bb3wQk6tPZX2+7+wnD8Qa+nBEgFQWfuvpjCufNtuBz7IF7UpbqHa4Zd2OhO2k63
WoARXFoB0pAMrzBF57wTO5Vwm01uuP627qj5JvuChGjxyCtC/vv/Qns2nn8sgu69
elkgyKSvqyNVTaSOh7d0llN1M7C9ktioGbKJ/U54OnzueH+CjkSv2yUhVvJ4g84A
jAo1RXpnHtgQtJejEjqSZ55Mpa5XO80QAFcxM+/RLxlT21zQWE7aLn9GzfDZn6DG
ZEmOOXSfQioX01SjQvnYMIfyoFp+ePSGuhiFva5eie9yEmGpAe4BBC7dcybpMlwY
Z9HfNa+DFh6DRC81rXYsdDJ2Ip8NrZxKpsRFZFIE3pASIf/cQudOV+3WkzTZxTd4
0JI1Jw3+lUfpe0obbL9SoyStgNj0Dx9AMv0gfTDt8GSJhrXvRUEB1j5ygr+xarcr
iLc6C3JnLr+MSDg/AIQkX2GxJBWkot5sZg/9O+/0Dl8R63MdU9NV/O6MZ3u2xgpx
Fg/C1qM2+mB5AnVT9o3IwF23/ochVNoT8xe8ZsPPniAETSwqTFavQEzwnA0iDKPv
Ol30p3gmxnz4WztoUBJWf9/Li5QdYwfZagrDbMQWVVu6/bPQo/2VQl8Vv/9FjRNn
3jVq228Mdjm7BjOM1CobcxaHiK6laW7g6QoQ/apxyDA2NkL1HEp2RLf21gpWODKJ
NoaD/MOOje1pxRJWFxcyYIvrOF0fTB8p4urdnpt/asYfHiHfDkzsMV8tY15PmrcR
mG706PA5zM3pxmYnfynRcYOBLbE/GK0yCo+Dsasp39WN7CGvTyPQ2F150GdW4lwx
D3ifcnTluqD/mRvvKHgNZ/9pe7SJ7zhwfajVda1x4SDzJ+MxBPxm00dO98dh495f
VszIng6yDgMvl1rqM1BNG/9AUlpkgv9lqNokp8yNfiJBPTtwKWHqcJ1hzEKsrQ27
Smy3ClsxEYrPlxYWLIw3A0miOqPldPjpyuJbARnJfGZRn531zRPT+TMTdG49NiWH
fKhPU5NPdBpdkZdgK5hyY2+N0d8thwGituNP2z5MOME6u7hS9Xa1b5/xxqBv7dt1
q8U8fbaRc1m7Njpe9dzDj6QgNWfpmmozVuAmIZUsgSzXW1dDmfb4sn4YLnT7lDZ2
VF+1wkCIP0op7NOyknQRmT7xGnYljhxorWY9KGzTlV/9MOq7Xd0DNiEYlCIZG/7W
Eu2WhhPx3D2KKoVX83PwJ5k3sAYGbPztgiqa0m8EPhh0MPZnV5LFaNm26Zm05Sfx
c1JwZj913CRhVCZLMoFP8PtFyjjD1Kw7CZeQ0PIa+jhqE7/UuxJfl4hvWYAuWjgm
/GnwpzsKCWSQ1k4MM3qvVgq3lgpAih/+vktGhwXZemBtWiQm265UcpPB9VvFxquP
UELWTQWo+4qtgFRi7iP0beIBqCnIWOIwfmv8marBNLqCDNeS0u31m4IXelxLTd/a
kx/tEJ18vE6fvUARRTpYy1Er/MI+P+8f/N9G+7pVWUaKey7ShG+DHzEthCKmFi+Q
tM/dthPSWMjZIX7DJrDFV83T6D2ICkbk7O/lyo5bV4RJslgVap8D9QjBAVpdSWpg
GFOSwEkn+6Da27yyJpq+ZQL3mOcsuTolsZDKcKiiiWms/fmz0TTvGCVJygErG0kp
/Y5cinT+xXGWva/GI/TpljArn082xYDQuAPt4Xd9QdWkonzTABLFo1Ghn6ILqx3M
AJonhTbjNwTZ4h9thd0t3qTG6KAgcXtF9W0sraPlRYaf1v8b2rvnjY1EWyp+/tZL
BfFN78CY5te6LhHAhmkF56gbYnxqhthDTpj6azSLeIO36AbbwWOcRqJbCxmm1wYc
cQs/ErGPE3TDHEIaJF7U/8boz47TmUVe84UomeQD0DFuNZX0g/qTjTVG50d9lozL
ZoFJZ4DJ2SBw+p8NLr80T9DNi9p1VOayEyCIJCHwoehEfEfS4q/fiQksr40nRHTz
PPqT/IEkd27l2eOzOQDeEGKNRJu1DwbdRq1lwwXTtt/iaK1pMRqC4WISbwhlw20K
9ecskGz5GHqOThbhxtnYOF27BoLrk6c/JWj+CCwGGYmes7Ovn5LeB3/3xp+Ei7WH
UltwCW7000wuAUyW4Hbc3j8KSz/8uxjTw6JLeHX4f7vuk4ws8jO8YRqAHTR09de3
mTW7cnQFC+UwkcnOAddX6aAAAOmfuBq8m/6nLRrrbvvty3LbcKRlKxbtxBMndSdm
e9+kJvGqKnoguk0lBUHD2tRE2NaoKqEsepiXyMHOJANquwiULTGQyvFJyshT8+eV
zTLQzAoMlNZ4q5QxspUZrr+a8vTrcFgRAANZpxymndhSmwwXYd+xHj3cr2dT90Uq
NyGmd1nf3tM0dne9dzjtcruZzNQH+38ws3ww5nkkVBRVSmW25e1zoaNSSe59h9wd
vrvW91UZJwiWH0TftFXvTbTJBejO+zjKFkWJv6a7XGE0tHH3D4s7VD09Gl7UbVmK
dE5lUIOXbEGWc7k9bgGGbDkvxuZNBpnqvj05EHxwTIdG7Dy86hEQh+G+RCm0tJeC
r+8/FF1pRgtfLziF7O2RDiWg2mhma6GRYR/7FS7pV+PyTqtv7HbwrnZDzhR+v+8h
iGqgztJnZqjFGxQDNIgGeP0CLLx3mXAIaDLNxe6wcpVZa/jyhW6Nbree1qcSVgyg
QKSVxmEQcaR7gf65ICOfqK3cfdgHEMZdd/k5fMr96gZ9Alj77pn5E+ai3nn0v4be
EsjHgzkwx0EnYNIz4HhNW+SrYvNK94dz6n2fCSrSqL0uR+w1yQNSGnAVI0KMByzR
S38cmXgHwsZ03g7QtW8KXt4EeXFjnlEEhl1pxbCuvguPBdisAl0uqQYd8cawSA96
ulxQCYXmyJO8WfeiUmUOQ+IyiO8m1Djm5739SPYqwNDFe/SxvW9SrgaMCs/ksNCr
B6HUOKVGnIxkTuNn96vhyUexnmvuirQKbozrWGzmmH5pvzhtt72MvV0v1cW2b8Ls
BRVDmm7909DajYaqAmKtWYJi5JVhQbPH5jDTv0ZrZAYX0WGqpLVmcvuKfmZjDat2
2Ks1DANuAmKekK/NGEwXCM1RPbPWlBsqado2e8vr9F9gwSD1LYTnaqtkZcIKMM41
h2lzl2U213FshsAOeDZl6eTYA8DJPCjCKvmDwsjYvHuWyKqYLtQDQ7fVOUkP7G7b
OQ+trHcuyXGWKje/BdLO1muxbEt96m9HYdDkkeiBkTBsVwM/SdVSfYUjEzrXpo/F
Mf91L3c5Q+UJlZT39xxSoMC7apQ74/QeVX6QHsjPKWYj5FHpx1s46MpSUeKUssCo
YajsiPjsmYjqQSTBe8QU5dkQDmbeUR3Kae16X0+c+1Zu7o+MAqAxJ/ExfSdNfCol
w9xey9KCPvrJwymziXkVKZk90V2uClgSBgU4nS6wl7UmUFpkTqhh6RvF5JN14LzN
NteJpFB3nUEAJMFJN2DdLiC5oXAfRdQRhDjsjX0FUrGSD0sfEifb8FYvCDbPbgdB
i21GaXrD6lcDIvVx4dX0CqjJ0XhQE4bOa52cSCb2IX0Q3dOEnVPqRJ+aFFT3LsGF
WeBtKkcTOfP5RCx4fnCvAKAXepbpksJWLLv6i/Npo5CWFSmLxvlg9EjpAwHv2Bhm
2oka84IHckcVuMccvT7UvNANtG39SNnVXCMOX2+WvX1LFm37UVbZKOzsqC2nehb4
3WZiDbzffUIKEEy3qx0n6ay0APUDpAp0rdYzW7DZdEBrEKzWX8o3u1DM4qZRb/Jv
osFMW/K/P8X56XO+XI98nl6UZvlxLLeact8TM0vKq8RK/USPBVTFItUcAXv6yLrD
Hi2lpUJygqEclZ/6L1jNA1QOtIIWZqRRjRcYHdKv/8jNgzzgiWzYLoVEOu7hNL5W
QLGeaZWFJZjE7R0p6jNSgm+gx/yXHriK6EaUAhZqd5EMESwKPVCa8zN8wF8pWxya
jID+cCO/NnfwCYZj7nnH+DrLgPMy+mSwVu9uAs68t/16srOsSxBu+YY1L3eQVCsc
TZvybPY3/Au6zSnMgk47oOkXRNoAl1wdRsA4TNbcUH65JXrDLc2viDMTuIuBkVW9
5ZZwIviJeRLkmPAaN6StkdiBoN6h0ggacwnY0H9AfNkucNp16ZmfQ4BK3uxk9TOY
hJvT2eKkKmt5zUMXvDEa7bR1IB9Fy8K9MX1BTzs7DRgpLbMg1d61LYUDIn3QpCAm
KuAqkW3lAk+cKieX++foKsrMYtDgyWPLjpt/bo2uj3kGfrzdskho1ze57cuhevwx
S9MPbi75QKiKNJSXLojgeQeVQNMfmlflT5j8cBxpYLeXiS4R0rWXvWo9XtoSAuH/
TksqYbLaAapCga72ztpmAQyUZuDzarSn5lLsjZXZ9zF8TO58SkMgfwo2aE5kB5jd
V08/evuKm9z8RiwmfcU9OOJbD81nodWDKUmXKYEOjieWECS8tVz7V8CQ0h+5NdMv
rAgKa53wJx0wZgD2esuj7JZgNgzrY2ZS6l0WAory+uo/MoZhpo6mjEpSLxyD+ASn
TyWXyZIx7wlf9pxlSaYij+c4X0CXGLrP9AWA7iDnRkrLSJ+J2ibfLr4qG7gKZhfw
9DFjctYVZYBs9TMjs/gA8P5WE3+8W43LmESxDRGCnV73eSC7eBLqHTGBv+OWtWKx
r5o++ArngjzrtIYuug7oE+4e7bDsUw6Gr/KnXXN9XvvLpsx/bwEPj4z2Arg7Xdrj
xHDvFZpRymSTBKSpyKd3IOYwaYYSd2vtl86G4INtYGurxc0zSxjMpkuRFxhnGo2r
5n2ruqEwueeSyighmivuf5jubWZT8VXXOKyeIBDSMvHHFiCttVVaBZgxXFfQg3m5
7AXl67Cc28AGYKPWL1GWd033FCNk/9TNieSN3Ovot7MZtxFRk/LD6d3Orowu1G7F
Pj1GIk8wKc0lO3GQLdi69Ne0czVQAvi5rYjdzDots6AJOnLxFspC4/wKnHaKct8Y
HISihYZ0WsWy5mv1YSvL01DiT07qbcl3gGvT9//MOCQZHpH25HThTUF2a3aYW4Zp
bfRFhXJXDHJlM2xlyxwRhxoh9j5ql9MNonhhvebdVUpIKWCogq1d/yAPiHBW/KN8
nyWT84OoBPbgtOzjg2dlEbU/5oGTCiA/wYoUqROfymk90exE2SBkCLjLsoi8rcl7
9wt9DeiqOt7SdH4tMc7BrGfxBjSM4KBViuBSGprshvcShYFCNLeGY00Id8W29xfE
9OSVMxICVaz/cKnpJCl6n8TYDwiJAl/l27hioGAWGLBvp8ldzj+xOLRW145Ec1k/
XXYM8bMbuDyKRbX1Bpnhah25tqsgHD5TEl6hPdcLAgMK4h/KFcQn13Cae11mNauo
pYK0PRI46TH8K3n4PsY2JAEMGqZPKAi2R/xqGZnDPg8D2UKjN48rSXiK8+H1Hoz8
8/DNmO9U2SiWrXhJ5CCm7/Jp0VBwXsR5tp6FjfMD76pkkbeyzR5WUTLwy/RZ6pK6
NH6bLhA74F/nzUeHVbEfDC+O+peVVYs2KPAHhls3lSdP32w/CUxo2JzShwL24RN9
OFJDsOSNduKBArdGTrwXDIyeOzmQJeDNHxqrIseR44dggUUcuxtDvrV+MLpZFasg
l0nCLqK+TVICcYwl7k/sbDctnUJ/qwVEbjg26it3ci22xuw+8wg1098wT5atnebT
9zhowGQorJ9fSivkOghnYbKtCiagYbBYxadMMpuSG7zZIpwxkkNZbhO4C5JN+Ful
0m2TK5uurBayFUYk709o59jZRHqHjsuplYBPq4ph5Mb4ijVs17xQlpBYoHVM7dT3
SacpdotOA16cXfr/K7oOXXt10nTQA2+PpsIY3Z50IfpDxWjAdFDVL2P9LzFH62UP
YKfIfMb9UtQHgX5TYN6ZEK4Ayc9OrNE9zg37mCTSrh7WFzAzZ7Mch+TL24a1L6Wc
TnWZw5QmsjxHfovXXgG+j1Yw31+CA2O8o/lr5Zs+Hwr/5KTd9lnA+RWeEwX3HDCJ
7q8FIOu7AQAIIsteS9BQ2kEZpQrpYlBa/rBwPpUP6zeUbIACdePcziDJoRd6mIIH
k6HG+KvO3H6o/x+VUp8ITHkfiKepzt5VRng0tf2V1iDVru7Y3tz8bsKNltEhzAqW
SJFyIMpx0pggof25wXr6pt2CkXNOoJY/euiuvysBwRqqulWIQ3zgGMGq2y4tQNPJ
pspvIv99NjAXw5B8fnqV50h01yC02HysRqNnqQe8K3bfazZs/BeBVG+7CHEt+xdd
shR99u2RcrBLJf8xo4ETbA+PV2dS8hpmew7eAhuNXGIAN7iIiFq8sJ7D2PsHG8Lc
iInlKCxKbBUnqbmT5PqedATMbs+cFOqWfZEn0Hs49UteI7Al+uAscquJMA8AfXs6
jxQ2yZLDZH5Aq9tS+dVvwkqLEV+MmkTsPsU0ngpKQLtskG4VZ4dgPDXeAdLlFtjL
MwSeR+Uzji+UXKOt6ahcjRwVprcAIz8L3iN6RtEP0zOSm96SKliPtrEtL46BToHH
Yo8sCFd+rEZu/+Bu2TBJpa9gBC+uATbsYGT8S0I//bW0RQ9jsXpudj32hNAdlbix
Nh1tjRoEOIRuqQO3cvJoi1DfKkBqoKAeXpTcpNPQzw0q0y7Oc5rJx9uBI8qQlJBr
IjmjqmUuK4aYlcLng/Tj9fZd0VtwB/+tAvT0hw+4+17TNQYdSW+85vhDopxwVKP5
ddVdIme247YLDC2AOxf11pg7uPcDlEo4y9bYH4b/Ja4w+qMlJAl5UPn0o0n0TJnj
8DB5uGouFIcbG6gk/wcn1ajMZ8bKgWWlXf4R8Rh0maHMH+tH5l1tZAyDZM9uNQZo
Y+irXLXif5DFabxIKHID2aJQxvOzWQYrpE2m9+N3NNlgoXBzOYBSGVpg9mvvqB+K
bla88sPqOdW9lIvX+ajreU/fS8tXXwMNRebopOOdFyDUgdmMlTOQyo3XcIM5DH5F
zbjfsKqAStE5zoU/HjaWHDbf5CCUhG8Pw3/ebENskiUeHAfRCkzZLMzlSP9mw1AT
IG01LZQ0mjwRMxuujuGJ3ZjwbWAZHHt8RmWxw/EU9s7heK8R/G7zjGxXcy3okS56
lbKm8oftAcMYXCndNaorPAfeSTSWsV6/xt7fqbTcmSOLymuU22lEBEp4l7rW/SmU
dylh9h5NqU/QkMqd69PUDqNY1PwZw41VBzDYvem5fpnAcm0v4CopSocC34BfI9w7
TLQse2RsQJq5bkV16XF/nkc91wK7tWzxc+sDJms7/KqLQUEHvPwPqnx4X2SN2v+U
wYw2/9WMxWzJx5Fk/YkKhyKRLfjECDqLDU5lbFWxqdgIuwFnO7/WtfT3wyWJziBC
1KoUbs1o+Gre+UG7AGHV206WZJwmL7QT8osJnSQBUB/IhRvGLcdKxqNtH5oNEASu
xebMT3UMRK/IuyFgVRtaBZoXcBzg8QHcHR4LrZLnwe9o5L0llL5JQle/OMgg5USd
ZAzOAtdmZK+mxK8NWcpZErumaPUdfEhmU/10d/7CPERm8/Ise6thgva/tu2kyXDR
XqbMgqrB2tvKo7d6wmmUvuXsVDbmUxrjBeQGFWLKFjUIplv945lwp8BsXbbTSqPo
eMY91OsxdUbHXbnhiZLzzU+/GtK7SUoOl+2TH3R5K2zTTEuqyUdH0s7fzPQ0miQ7
AUtD/6Z9ImYcdFLWWnW8eUVxGxCmrAsNKdNE7n4nZAwez09S8OAAOjX89SCgbbaI
LGEslchbZ967tfPaWjjMkuYtHVaBc3ARJnKTpFqZybP0Yoz17sUpoObyD26p6Pya
17Y76Axnceo1aWMPcYiVqXDnVkNYiVwRCQp/u8pt5aSwgEQilxeBJF85PYdmAAZ3
AbDnSsvoI3ys3FPtWzyorOmMW6TnJ/oMzzVxj6j9s0hnmmZ1MhhdDfD1oVykwYqH
NSG5I9X58g40TTQFFlpSalOu8ida0gelK4jBnxE8dAvWvomJWlN0Sl67+kw+DOk5
D4CzJhjWakaOlwT4YQsCQTQ0Mtrqt5CAcs/bLlpMUjZ3PnjanHev49AN5yCgbu+T
cAy6EzgFcLU0A+MhIuUr5KfcK3zumiFlbrQpZnwSDDHcvXdb2ezVsfNqqe8Qq68A
1H2Qnl6PNR4zNqJCsNqK/1c7KY0AvjB2+BSA2U8yOOSa3Q0Sda7H+NexWIst7L3d
IsAW/u0/SYw++XMZGt0lMA==
`pragma protect end_protected
