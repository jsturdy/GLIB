// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ABMrON4d7zhRI+FX0lRLs7IxSNzvOCCtjFa6qAFW9CyxYey2gnolF4i/5szQ+Zs7
my8/adRoiJw1SWC6OdGcX4xGIzE86lBEG6hoQyWs8BzKRNdusiFw3mMAJUkAXvb7
BbT//kVh5ig6A4CH+O5l+9OZ6fOVAy3H+9w06khTn/o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18944)
rzTkx+lAr6wRCc8vfal+EIbUdUpcUJd7mCR2RAkmP1ETbG0MFc9FVy0JBcxEAAYX
N4/soWc1RD2cbYaUhM8IgXW51kJc8XX9BQ/mqAHm3+YoFh6KsOJWujBtZcPbDQk8
6hOEpIaWmRsx9+nBD6NlfziNLODnInjPJDsJdw5ICVUjp989KnY4vHUfbtFVjbHw
5gQdo2YFkarlnKrS553XwEZ0jeCtNlnWLD0X3klGjWqxcJ9UtTXLTJzXRhYx0p5E
JUoecOCGg4Qkr9q228UmOpqJHl5rTZHcBbby8plGjXqUF4yoNRHV85kBhNEdMBL0
LbYOmgfGND/bEgPO6e448KNZxy/6I5DYJ1Vj5n3ct7qnDeu6ucex5kwduk33hvVs
FaPw7De2mafc9bnfBmaTtoYzRdDD6xEjkJWEOFhbFdD3qDBRlVMexXTbvHr6deks
VobWODOKD53WQstNv8pfiteCFewRpCqwn+/eCMafI6OHbBEdQ2RYDV64BiJKHxuQ
eUNkQ5PqP012W1jQH7oa6YJnlZUDBwaAwz6zsqDf/08tQw0a/GL7229yxTGGxaM0
bCvEK6neicnZ6pX9FcM9sWFzbmGRhKtpD2V/5brVwsLCF2DhITImGuoprf8b8ndM
Hkzxv+nHhaBXx1xOfzbOph/Wag+61VPGxMH+Ap8mKgpBksKx39PPMwHcL9M/tnkY
qy6ratdxCGhm6+aWpzs5zZbvwqSc19MK/ww6d2q7vYmH8TGjakp4yaAHtAe3a7le
1v7MvT9C8W4WHJFZ9uCXu6tr7zTnwOL4jOTXr4X3Q8Ly6pecienn/zl1sdzU3L6a
M5HfOivuIjqBZ4M6jxbozsuXEvPgesYtjuUs0Ksf6Qz7VB83btp+2yp/01yhd6Le
kj4X+F8Enj85eOASo43D9XpCx45PWuYrDDCBFciQD5qTTafuP04kcrLSeL4gJRSc
/5CMXMrG7ZVVVmGkq/H9AR5wcaO1wNYm/WqPVzRvsR6/gwWrnDgzd3CqArKVHkrL
NFKvLp9kh+66ZmRgITlJO9e4QEA4+ujPoEQYwurVp2XdSuSt30XG7Iytj5K6VnHH
yzsz9uuGfA4UdNqZUKsDdlXKPnji2T7roYlvF7IVvntH554Sd5mPVQJg0O2rYKwm
rL9h1YZA3LalBBHAVysVobn3gf8yFnYnj08X/5VnkcmGCYIHh85NCxfaBx6y/Wth
Gp5QQsWmqljrjmBXZ5H1MZMIAXEPfNsrweajiWqMHeClsBUoOZbT6s3u43YGsNQ2
yT4e+iTW0tSEHIcQEdHNIrpX/DcrZgkscQK92rDBvwsJKd5D6f/BTRNeKbF6WKpv
tVxL1unmRp6wnQQTGzT47GtFwd8pIwMDsctioB3y88W0Pj9h6FOEH9l26phbWN4/
wVMYhWDhp0QDcwgYuhqN4TAwHwMo6MEJNGkjcXRjDYUBUfmXv9GlHsiKmWleK4yE
HIUdVN7wTAv+kgPYZFuYz5I/Z5y6uu0zx20quAPX65hw7ETJQG0b04pa5W5F+6Bo
ImOVeH4tyOgjBIrv7bZ5etYwqwzKLvchJL7kJUN+tauqT+FFtykQHhCOjJYdNHlK
YuKHzKLQgHa2OrbE/Hul+krqN5wBcnbd8QnoDK9gdfjZYvpfjXdLda1XHxjcNB9C
AL6tFwyqW9Js2NdiwJH5d8TdDsRaBPIlyW92sGmoH9X7ZlefVU3S3v2hxTJt66wu
d2QAsY6QBNhOmtS2owC/g7QeNEFSZgzZDngxoHBeDhW4QznRi6/1JrM9JbyaNOZp
uGRRGxpLPolig9HiqXd26weFU1eCgc4lvgwVqFEQVec+UPdgPy3ekz32m/goT35E
Vihd1ZJZPKHbvdFq3bllWTNGhT8Dp0AP8nraavfGJUvKlbgJ5AJEAKB50I8T/brf
iihZRwN255Akh6PokNF0T1Wwrs8r2QRoMoHE2qVPmC0zm82P9sITMfqhWlZfwPVh
DWQ3znRvMRgCAnv2KIqvatKrluiEMuHt76G3N4Fp6VLo0vXGjdDQS4xpBHMjS+Se
kaPJ8LUjoQOL4bnKIVRLLFmmnjpNgn3PUKTXU2sEkffaQ+yL5M4VmtenK49PFlU0
X+4+fsBYOCoeXnWINhyWSjZd+7L7HEJdLEtjaw+Aq701vK1rrclkphHuM5tRR163
h4AVX0tDvDGCH81WDERAl0OHK9lBOuZBsfA7wvumOhGIae9JuxWDC2T8ZS3fV8PB
Vh3AcWJc0OIUKQIcZIRPCFMR+JwePjwTQunPur858vF7N2slaX3YGKXICgF5+/Xt
W53RfB4NKcxzyaQb4RUMqb37K54CHbu/mvpwfhz1ZnkfHCkjq0M1yL23DWee7X9p
2f4uLQJPM0lRhAuF3LsGZkmRfIL6qZfYAAUaCaXSpCwZXGfEvM2UPsyO4kZxRpNu
ygxIjEhPmBxW53XrUDjW4QHMTBaV7N+5dbuZWnri7IbaAVMrVX/fpvPzNwOcD+JQ
85qS23xuD2EvViUKwlAWGz2UzVmEP7YNEka0yD5ww7jR+mnB24j/3Fq/VTzOPFUI
G+I+2ixc5QMsNuMhYY4WzVmGZEfuJjlOYMbTLjglZ1yFzLzrauNzEynZh4QbXFKi
M7GyLU+Cn/urR3XigGBybQYmuA/i7vkKlg2YI2OE+JckV9CeeRhTf+akCeswMlTj
RLbU2tajHKqyJ76T7e0Fx0pkvX5tlA0erlZJrz5gGYak+CnFtvqv4DaXdM1PRH09
1jS3SFVrTbHuqA6i8lss78kGP8wUMsAyd9B5LEnNbpS8j/g6K2Qhx2GF0K9CVRty
YtbHB6A4S7rZwFEf9FBpEzsiZ4EzLJ9sY7jxLXncPQ1qE0cWvoNVsJOG9fFNifQM
UPd0We4gJXic5DrrSKM/6GtyqsnWnoJT5yGajtjovGALWHtss3KoCkgsbyuBugbc
fqHceFm2EisEWco7OdInszgScjSmdtJoNjH6UMjZxDb3LpYt49Rw0NyYWbuCghCr
4WZdTEYmd3G0i/N1JB+eZpCe/eNJnMkOH3UpKdoQOrkgU9bn0LGuDfR5MEn5jhgu
/DNrtnWccnFlHffdVHUg9KT59bj5+HlwDZcqU7kMQQ+qlhdV3tg5WoHRU9g8TkqT
6iK1FR9Jbq43DkLqaNNCieRmZ7ZqQI4eUvIWNOycY/HHwOypVnQ84v4vrqJWpHha
vxgT6acObL+PNfm5jR+vgDZjRd7gdaNbETe/gwk+AQABDwxzB5xICu8sVvha+KZe
TxawSkCd+4H48qOin5a3KJ0VYDVLX6bJCTQ4rmwEwnYyZTJAoOdPSvJX9PR+iPtr
9BZ8H0ihMN8TDPXCtMPbFsebWI0S0XOzzudkyUPSgGMsZAOeZb9KJycNWzDHhDyY
10VDvxu9JCNvvxi18rBIcKdFfincsHjgK+UG/KlvdvazZUZ1i2cUePkNTkXRTxQx
0uUNoD0f92Nm4uQSybLMn+5wYl7Az+SrIcwUi0q9kRpt5DLzJRIVT2JXHzcyQQSo
X+VQ4EFNMNOBegdowBgvrx63R8nsUFuqQbD8g8hd1hL820x9SfRp/13nruxsSDyn
EO39fZxvN75lEpENhvqFFrzJt3zGMJf/GwpR7agXd+s7iqFtKxicrXH1SHXY687i
nJZNFdrms6UCPcMlEbBiMNuDrQ61e3/HLm6em83x6nl9OV6y8G3JrY+eqTLY6P5l
PAKKo+7+vg2WoUH6AFvXMXtLjAc6Eiw+dl8Y7Qux2WPVIGtcwulRY68/D3z/sxf0
3wq4VApiCR5VjZA0rHFBYgjoN9KYzq1FfITLjiMgNM3L3qR4P3xokk5JxZgFQTVb
K859Q4V37rYgywcdxbcYckL+qP3ryzUiH6gHIaAanxwzK17bVt96S3S8JLWm4q/l
ZZBxeRQn07uZaXC2hFGFLEal0uEXcxkIdVYS5Mg7m31RsjNK8Amd28L6giLtfZNu
2nGA6ZnIwjXeGh8Z6/shl60VSFPc1q3Ng5HttekevWMfsU0VKGL9guiGjV4Tbyl3
Oc/DB0Qcw03QIoLFL1sCxrbHQrRar48RUzMZv604MuleUcJVv4VqFZjWDlIIuX+v
ops+zJ7HPLnr56GyHrbkwWU+sL87G4VjoP272FbOioqX8QBl17u7LsXCmF1cPep+
5f85SbRnl+/qUu/JjEeNFXslulw1bv7bOFzqKeRKvCQIP6VT0L9EGNUGo1HpcOMt
GTYbJA4mz+0e/SLqG6CSUzRDZDFxQU7gBSuGmm10GM0JBpT7bwTD2LtFA+x0NggP
HFgSnZDsPZdHgjEIwYx5b0lQNg5Kw0OIG0RaJuUms3Bbpflef2UoMbewvr2o9wT3
91sKrCTGjpzcZ7sECEQg3sqrNqB0N1DriYJTfG66PF0VzMw7DAHfZgHJrlH+3IPY
E6a+Mfjk+4q758bi24rdSUdqMujhMDrQy1ENovBYnYpRI9vQdypu9/2SlmJBeh9J
Qgc3asi6+Aj2JFiEuhyR1JnKZfSS35LKpzW1+zx/5jmxC5ufVANYTg17+jZQEKO9
aBqbcwFpYfxbUOdBGQK1be7uPNGzpMPzmtmh8o69v+3zXlwE3DbxhbDF9v33PFQB
yc9jMNnJtRTZimLEktchj4c/YUgS/ZR5f9ThgFsQ/dM7DwoU4Eb44ms9phkTRL35
dWHMqNU0iD+rHfKMNVVfLTpwmaTNV8uUfWDLSbBOaXKH+YvmaFlj9UTEKlKMlYZp
GwuHebUMwF1r741nyVPU3iYpmGUkr2MDBtwgZtGRx4CRvGZOh5MZiei0wBDxmOIs
tiqfyIvsN40SYAtVkU9lDGNwv0vFiZIWR/vQcr1uHj90q3kPocf2ny0IVnh1bn99
yGE69m+fokYrR5CGFXvbIOa2HRxA0KPq6s9EgJZFoGfr6VjZME0sm+A4i20/ZD21
N0/bA3+PldI41r6pfl1/q9VNC0QRT3RnjimTCO3FWIptY5Wu/IQ/BkzpQhZtr4w1
7THyR9Zvc2C0pQC0Uuqg37owwts7v6JSn2RxKXa7BRKNwjCg5D52dzZGe9FZdQG5
CEhCNtNxEZvCSwT+SSgMGU4k7B9qowgmqYYXzcG/GUiCsQyP4VibwOf+qa4sgEfs
oPSDdf207JxqKrP0BeXIQkRMxEZAGhXmTVsCdIxiCkeVSAByFFUf0NwVvLteAsRP
GfXf8PKy3+ZbhpGWchNflhNARhyyCyNKdM0qKayio9vQdpPRHZp8hQVDdklIHm5A
J4l7uVWe+ejSgry3blmNRDjj4cb6XKOaAXkXU3IVyPiYr9NpXXG8uv+XxC/wMPaM
mLlt4gpDiRoK1NnkakYa7HceBGwR3WIOw3NBNEQpPxippJulsLgCgnG/8huSdF/N
AstEfpWSdzpk+1spAU7rpgurE3hHIHqFMq3sW+cShy99RIg0O9HT1Q3xNZB1XLpi
sAwiMU3dfNHdM8IryqyuuUOM9rGkqeXYYIFVjdczy/L/dCz95hpRqHpNeSVCW6iY
Zg0g3XEBUw+hsIVaFn4PaNTHlrIidZMmVQlwz0i4nSCz2TBsOaGw6awrTK0xz5UL
8lzHMkF9nmo0vU1H3zqUKoTTN1mwfftc4UtKPjvMsZYn/G7BNveMm1T0AHJkS5io
reeBzM+te8SXbEhgFvFiySXD/4JbgWCrNjt03vvHt/7+QbB65cCQ5Rfx/lyMOT7M
2IrcCQHCVrU636+SAL6g5chMlL/ymgV6plnXu3C/eWIi2PRBpf/u4W0GYzTz5T6j
EHmZ+XxtptkrZ3MQSqHfP1lYYxmq64Qjk+PCY/inT4KeAx/55aUj4QV2Astri23u
850rs58i3S6pZNJc1blRzR+hH31scD5pqmWp5uj9sXM819QfyNxTvQQHjjNVSxxX
JH3721f9rd5pqTsQnPDdIGWyPK+DJCSo/9jgZUpjvZMBv/d/bO5wXYO0wjelo7RD
/L0rPNRrTFWrlp6kMO5H9k23YgnxOoL9koPbD0dDvGoIQo93Fb9TOpqZKCuFMMyT
DXebx6VHjADQrXDyXkqcQrIWT0j3ajaqpYyWsdqNbWEa6MifHnKRCHIbX15WmvJO
pOz2y3EOpThR1r0bLAa8+rzj9MfYqxlt9RE+UgQ+64LqBere5mjEhyi5P6AXdYJC
+I0nEsEZdlSYzxwg9Tzv7nwwqDTpkewE/ZypWmHwAsBRUFPUwBZ0ESPZlJ8iGgqv
EAW8I0MBM+P64wA48uF3QgHqCPWt4TXiRUdl9EPCAcjvz/ftK7BxiZxDZE8Y8pgT
QXxy/raZiZNem/xBKRMyFOT3AEIonKPe9Nh2bdYx3H2adi9mPyGDTlZ+MbFXZnSb
jR8RmMmSbMpCox1S08KUM5pBxiw9PnXGKx4qJNumkFK5z1l2+uo2+ieUXh2QQxIV
9U0PzpE6LwilWuPNC+GrUCuaFXMVyDfV8FbzoAEJOuGbjfXv8m5eZIZGFLLKcNho
rYuiLfOnMF8BtlgZQ/xgQYxv4hzYIi77UDFOZdklSBsNTMgAXxvvQ5pY0n98LGwo
fPg7H64T2J+rTD9eW8Wq692vfAabkfw1S8CLnbELoqaT8Foxbx60WRqAGAvSpYF7
tf3COYNvag3vrHYYvFEXPGRSZfs9TrMPX6zeq8l9JpemyTihFunP8riQnggZS63o
FR1hfTDBiCKeWnBOceQZfN+3S4WBmuHM4tbKkTpTMM9UfSTI28N5TXI9fadIA75z
I1jMtLbGjDGhpsPFji0/AzEN0gPbBObjUAbwoiw/iZpi1r9m8/gcTPi8rCwlR87A
Go9mFM32MVa7m02jGdQp3fswtV/A1jSmlFp2kybleLWO8R3njN8LyyKIksuvwXIc
UBT+ETejnRvATOss+lKT/xwofKRTcgRK2vSctRdLK3a3mYMVY/HNLZbvRZ3quOoi
IFZCtsRXIvdHl2Ym12hdaDcGnHaMOpLXTxjPh3YRPadoZJ81OpOgKlVyRxTpewRJ
+E+gg3VW9/Wv/psYZV42ZniYBaSkPh4emClA+7QLy/H79e1JcMvEwBM65ybWQhlx
mcDU8/0Et0A1ZCT97VoXXfdfZkKJvdlCqLSoOHKtdoZzNUB5oLqEozUTRQcNGBef
+ahbLM4z5YvBFaVHwYlUuJL7J4ejTSQhpA6qsKFlgRfhjt9CfeXHHnEN7mbHC7sT
vcxxE2hgvRDceGc6o5Ke/7KRePg+NmF8+rV2Sdkqb9Wx4b47coMxrJWbciV2tPb5
fgxI7qbU529vKQkLgHdWKLDza1LKEh+lIYsjA34fXcJ98FeTS+hzh+jjTu7K6MWE
2tBcD/2fFzZ5TBReLh4dP+QlV2pCdjbOWPGNhWheWN2tfcTcY/+c9ZeVur3O5iPT
p3h2T0i49Hv0/gK1eJSG53+BRlcrAkqPlNogU08QxdsCObXbQEKzapMViNWAiRjZ
SyBhDzR8fSbWUzhEstJCwEdb7TQqSMk2+r9XgmKqEir/jMThBac5nd7T3371k/sQ
uaoRcenBOPqWz9G1oAN//0qtLoXoLdlopSdR3JAhCZC5ely8aFt/IOgr1udg7HWI
bur3KyLiwfll2KHc6y5Qemark4cJlNlzJMr5yGcw6ZlfnjeYHWlUc5IqMFa4rT4B
tKWCAmjbAubA/GAbdRu36DiVo8Zqe/1ltjX22sdlvTjluYxkZjHGfS68o3ZbWSV/
m8c3lpB9uz78KwSFH7lbNjhb8qIZVSjDWKarLe04SFsv0awQrk8x04Ebgjmy81Xj
le0I/6XSoVe1Ki0F5lnjYJTzOxFvW9sDW4DBkbaK0J7laKDb7ixRgWMQoVQWXh19
uV5ddiSMeF9eQKa4Kq81rS0dsbFQsjBS+N0zlGNTpXIJgNBI5wDFWAt7sQ7ESSgJ
jV+hF6lEdLUdavuPEZjB5klLuq8z9SR35Hq5/xTLkGw9s1jzNuXixtUhraTy9ofI
p/6AmKRorcPntd28yDKEq/RzWQ4jIUBoPdkY01lEHoII324Ra66wV2qhQoQ8bRD1
up2gtKsXqWOEJaHGP2aHqIaOZLYbwylkkjvBtLC0Z1zuqSLwKzwreNHYcnqWCgUk
7Vk0WWI25LpTjqNrlRObgF1b9RoCw6mkatu9gmN8/NshSf924BVcfWqGu1Bg6q+S
rnf1CYJ8MGtymxrX1VMNBC6AoBxIoUoAXX9aPCj5ptXDEqScXa1RDlsR7feWw8HE
U2h0LvZv8z3jVHJF5asvMdT3o/l6r0KJIcnHHhwUdrCmzOu+O126j44q/BhsqFsb
ui7aJWfsY/vvL2tMaLLhHIiZA8Cy+t3DS849fNbF2Ko+8uECiqhQHXu7x/qSZS8h
IA89RRSBPRkIBV8YPvRGQQ/SGwlsqFAPSVpQCYaASvnbvz0unFZM629NFYyQqvzE
uo2/UpwEUtFqehpweo3a+o2Qiw1GZGmfSGd/tgxnfUSxlvipXvwNqRXj1rdKtm4r
Xj6TU7sKqz5UAdCGf1vUy3rmNNbDEVUY2EnYB75Os3x5nr47TbAuZRfEc8EX2fix
6Zhi2Tm/WR11tJFWTiUglWgsrQUYjfCqK8q6Jya000jhuvcG/YfrlZtjItksdsRf
dDmfnVbCQwWHzLkISGHDW/ZkqZ3Hv6uoi98T9oR8ZjC2B/2L0w7lAl3yMs3gcEyD
2Y+96EjENFLYH8jfLbfgJceKtMSh46E8DJk6jxA1X+4Np5kW+modHkub9zzcU7t0
5yaHn+37JM69fhmPEFggWKrWpb852/J47JFq6LUF8vYAeS8U3VSw3SMGI9ir6JGt
L1CmaFulJy3qm9U6Pp7/eya8iDIyUsv/J/6agG2fOF+OerhWmq3k9/ayNmkyWHj9
RlvH3QCUwprTq09O0SbtluIFVscX5pJKrGSfph+zmFKmptHc0Hs8h0ruwPvdlf1r
aEepMaHk3LnVQCYNUHMajnstLEOKdr+Ncydn0SajsN2NDH2ZpHvOD9Jn8QoWhEKq
DkbTYdF4AtCV8l218ujhhBopdltLzVvtjsbYeeT5p6s+IoE18K3kBXhPQOxdB1xR
8GketHO8bKoiApN3EOiCTUvPe7cxZd6rOQMGQdzshgEQWlUe8dmhB1vlM3v7mXDU
qtNR45hMIuPS6E1SLbU4fSa2t8DrpwjYHVsUKlvkYVnxPjkOWawK6N1lmShYQhQv
gQBVGaqL1pr0xoh+LWGJUc5QcbWYbAquCY0HwDqekarOsMTPM60xVNMxDzMl/kki
GWnZBE6/ZYY2P66EbICnkBEF7FsFLuN36MVP6tqFtLJqj7P4cGb+puzLAGGuAKyY
eJRKhV7F57Gk2qCm1YEOlocwhsI4djz0i7R2YFGTvQTvB8yRWCdQ3jwdTe3OZVkj
G8Y06+2GlJtPlPMTSLNUos5xq5DmKeO3cP4GIZ5VOh8vDdSax01H55VE8zbKsPtJ
B2pDWLn7rbLIuCMKLfQ7j2IQxeQgvi8lF6xff9hW0bqkR837IgaMVJsx0+90gDKf
gwuvc5BV6CmB1gn27QozYw2mfAwUBQ+ZCS3hqTRmI+INswkXOASWHDjrSgvIQ3tf
vpgq5uM6oj7SAk4ixXUtKvgfa4f00sQO0NXVibOW7IEwu7PVU4rb2kN436O2bQAw
iRF2v2hEo6qdkiKNR3I+ApcMz6LyKJVjC5uwWlQEuvLjsQZZ/6LK4U7NvvEAzhSt
mxkGZQSCyM3/xrn2+Td0SHIn76zgLZXFAXq6vSg1EaPWS1WiekzcovKVgkNU+u3M
gawpGsGRlVyj+bD072pi8MlQDemNRFBbAC7RoPEnOYtz46+sY+ZYxObJ7DfFpYcY
M+yx0aRYXIi1op86S+mE1e0hP3QqYJFM72+vckeU2o6orRlZEaka/UTJkio1B2NQ
Q1j7/JkLmOezKe4qWirjBlgaKQsbzrGbFjOySOS9QKR5iJGUlNwqRZmOoloPGZ53
VvpZfr4a/SrDb6Iu9NKNFHRFNCW/po26Ce/6j4y4EBVakeyXHHZuBBVLSxw4kJrU
pmQPQqGe4EUsT4UeMEUrC6dLEzawOu9O/tyMtj18pwo3uppBaG2u8a2jw1Tku8GY
mNqke7FQbivtsbxU7S9MnuspcHS+Y6O5pb4QSKFYD+ylMS2L9QQoiwVzCblxTaBx
n93P+l7uA5SEm18mH+n9MuYG9XD4fC4oz3oA2j/JdQyY3UAwlRWDhwNyICN+55a5
CabTjbf8RMnJBaxDfiF2ayxNix3/fyCCe9Fef4QWrNpmdELWIlvVhoVyhXfTDCOx
DDS2vjLDPv3KgAaFbY1QJyvGDSuczU1RLRFP6aqEma4OyS64tK9jSBBr0lRfaod0
ih8tk3sQo90BBxMBwzq161va/yktXpzjAM6WwMppKEVsJD7TxAu0fvDmdNbPbZyx
ViIt6Xtj9MKzjzjPPsmt7ue6NNVJsoptJb2M/ldiA9uLEfoUoXLuE7gb8HR/qWaI
R6g0cx1wjNot11sQu1QfP6Cv73P9eh5WPNhQRvIEzo8ewRRr9xqlSXJ4Wd3JrtqO
W2jEYWN6yBKaqCPDvxTZ2ty1mvSD0/yT9YG+rmXu9WeXsTAhO0tRlK9kZugmdxJ2
L6p5rE20OrFg8IQBmNAKNpixsxGIbcERjTEju/7jf7ITje95YXM/yA+cknTxMif6
j7O8/5gYrx1P0eXPsaJCygpNW38TuzKW79UihRYEXn7eIs2kbnxc+QwSeLtd5PAd
vZ/FEmHrnhRVA/FNXKKXBNJ5mtahP811UsfhCJL0LvZVD9AGcEEPgWUg87ZNE0HO
lhvIHmodrrJ6s8UC5FOImDPsV5obAflcjIyl7+6rdpYIujmcQfDdi6aHkmmqvzFR
Y+klBBW/3fyApNIrCNWl/ogkcJOOvVRQ4SW1RHDpZOpm/WT+D08sNmyzLIljs4Ot
xSjsvp/CqbpRIKUnP8XwboeF3d8ztqEntqEbWDrvZcuXIuT7088qHmcRJXZDK5Il
0zZOLi6VpJLiAAUo8IBntMTBI8JiXOydlI6/bWnNNW5KfZ2WtlBt5mYNr5rurYIS
oPS9LqkDvouqFTyU9EpxzPCMQoddR8dwA60c2t5+Yya7ABwAa2N6NWP52zizV2xB
N6bERNM8IFONoVUBBuR+g3wKdSSJtUOs5S76NnHVZTs6+2MixEi0IIjAO4pNEkdy
wF9lhTx3Dejau7682Gq/T+pU1X9k97LwuxvYV3t/64wuO8QPRxgScDdcOaAOA2x5
8o3VGuz0PzoSdJaxq9IoBVBgUL84+QRKXD5/GnMltM0pmQZDkxVNjjmr9viBgb4n
wvJ3WC6zGyqhGWWW0rE5Mzyx8vMo8100P/xcmlC35YHsCg3ay1tpxqQM97YeYCuF
xCtPFseBTDwQAUYb++vFaFIwsFDrrBdqK0G8JVhOlVSr3LjB4PkBeXC7KBGTH1So
58KXuilHpu+kTL8AU6aN1HXxYKowVk9+5oIRoAMN6P7yeIE90uFMBoF16+IQ/rD8
cmwgj4Wz5fSoCuiEhdsa5QEentO1/KEBlFe159eLKVgcFn+mSOiUecvZrX1V5xO9
rXu12HPjb6C9ZICrnbuKLTetpG6f0e7dLqIhLB9OMG1dvgLipDtKc0X2/11a+e0f
+6lcmv/QzUjxnnJsXRraNFMM4YM0458Wn8akiNyQeLR3gEmzCPmUnycFtGIfMNap
GVef3jzUgnyQl1nwH3zjzPh6xTifQ12OzpQBKJaSb08xyi+r0Vik61GZZtP1CkWW
F3ixZu97+sp3B+R9WD29C4695kQGM2vvI2SJF93m67J812jIUkIDVZSb7vlvlxsG
N+O4nS74D5yriaHN10QX+fAwoKyGCZOuZmeVo2D9EOTq5sUQZdkIEiOLXmRPid+e
2YEZAN2z4WP2QtKx3eivFf00stR0C10/yo1xp4Q/aChC12cRUWDw9h6yEPPnjOVb
4uNEa9mvKxh2+UE4CBg88K17hWmbOoKkWU5dLEAJpA5uKLelqZpEkaUhg/RgdAgM
zYzEeJZ8a5ldwx+KiISUkcHP64rebnQ8Av9IrU1MnQ4HNgH/0XirTp/eXzmfkXP2
luXz2wPBnzRz2AyxOdrm+1Luhj2LRG7zfNrrT95S/dWuLcCsbIuxzCmeDmbqSvzp
4xywrN4+hkKyrIveMcH20EVyyNEOZ70WasBbnFLfryUAlHyl/xrwZq+TSIx0SxPA
SP1FZ+f6uXH+ormMp+9cmkgxEwHygkKuNXWhnxOCNBvDzPmBHgR3D0aEBhKNCipK
OQDRv6LERIlqycKpV7wlS+ZkzzSIzfbgVlTcyJ7z1RCQuMy+KM0v6fY/vY3Jo9N/
sp+Z+dnMnUu4UTVpqmxTb7LDdlY8jehRdDJRbQAK7B2iCzrwCCfQ0Y/K4tZ+Qz0/
SV6/LmfzbaRiDxeYQo/UT95DZTPaamM2+FT9TGJ9KhWMZqhdOECIAZkDl2z7RuH4
cE8Pw4rNkJsDkoACphvxQOs/h4FKUheUhIlxWzqEmsqTq5JmFNgKo/CfuYbGc2h4
bxOY+0wyTOupFstmmHXP3dW5vlK62RjS3HiVxPkewZFlz86cRRbjl0YNsc8UeMuk
rHKFWU8LIFBS0Awme0TDQQOy6z3lR8rzmZwGYF6YWnJdEHXtTNKxhkQAoq2AN+Vh
2XXgGaiqpQtdz8OCe72/9FKpX102fa8Rl7dU3No+A5ZTiNadqzkPOXTP/8U5WMAx
FwCrfyegadnaDnRDkN6oteIFMX/aJHcAZRY7qxFq4xGPCm1CifNpaCMNrPaUC+nv
oCd85rtPVcwdRJkdkKGpQlhASmZLHs7MXTBYQlYE0QkmgtU7qR935+FVocHNv5Fa
tJFinIw2uHDr5F+0ZyZXso5BqaXxzwsJ5HXVSjfE055A+fDbIjkHh7rHW5ZbjSya
4DmOcvSr3Nlnlr5PSvKzYLZMr+ZnnKQgk04FCy9DKTLCDRyK2m4mPXtFmDi65PcC
75TRswLRAKZEN5YYR/Xfl8e4fEBxsxN8Un7L1fRy3JzIWPQwU0s0RukJTr287oJJ
YWaZ3bu/5KvWAR+NQ4ik1imdnwrPm232SrVW1RKZfSwygy3MGsLxxZmxtPrMw9mt
ejO+Avxz+g2VATp/FNsw9zNmzBfj1b57oGfOixHGwSzJs1IQAI1X06crhhVpvFcR
5J069KzAoc2/SslJxuKzTZPgBi7eNtRy6UOLce+Ex1kqMWlpHxGdSrsRahG3mPnS
M/sc+D2osp67TUztgDo2YHrQNQXNMWyd+mLZN04g1lEbPWnnjvxIaHvjU/tABNRI
Lymw96AXIfPCliZxNAeDZiayRGog3q5O1NrY3NItMLEVsH1hFLU06Eo5GNUgBAk8
FrrlAbnny7edfJqo82VtBcJEd8p+PTNEYMoDV1ObFiWvenWBEtrbxJo89DyOkkwr
xXF9tSdM+7UmNC/nl1DsHbxCm5aEfBm2di2tVUiLeVweoOe0omL9GS5sjKFZMMeu
mfTJyXooo2Q/jIzP7MSjTVw/HdBtxhnJ1kpN7MItqRA/gX3InVGj7Z/lfeBHnwRD
DNkorEgTNJsgjYk+sEfbfQU7O6bMaLqIHL1aIsl/LYfjfqx5IZaksgxg84ZVnSy0
te4kDzfHcoy/gF3p7WIkuIlXObGbGyKxKgx1Nu/Mdwwb5QpNjTxVW8Mw0oVH9cxa
4ZM8OFkpBuEjJ4btL3KaMDsTj2ZMdQuk4jCQR3m7B6zacxXVD9n+5LEFbu9RhldO
hKsjoFF1Uhw+OidVYyI9OtpIPInoX1koOFVYw+Wbn8DNMsnjMaZMfb7v16Wte0YN
+bIPN5eC8SgJ2DWB5wQz7Zk4k5ID4zosfau0QVgdnljeCl5L+8RwHZm/Xr9NEvwR
+mxx7g7l1AWMqbkdtXt9HKvdrTIYjEhIZ7DWdeJrGu01DtLw4muRhWVxm+ImwcUT
q4LpjHpq8CJvP/jrzso0BUMVAOQOL8K+mE28Gvqgb/lfRBxn2aQG5YOsP5yHlxJW
cQ2/MVfErGOHobzwkR0OWDt2r1z5/JTTcSA97+CSty9xNnUFXLWA4nYNVqNIl+aK
SoLhfhAx4/p3BieBCLr8sqR55X657oQUj250ZRsTTG4gq/T+x9/O/QK7giz/wT8E
mByZEzhl/LOkBIPD5COkIFvEoTYjfvR1J8y9Pl4b6Xor5AuwmxpvrnvkgirfhOru
804+6lD3LFwA2yVPVfzjLTP5KOdB//7hs5UoR7L3uJjkbjieJD0xF9lfTk44vBjt
dTrdf5TngOSTE4wTT/wa8VJrPDY7Aa1aphTe9Cnz0qN2FSYutVgxnVXI39fjDMnS
dgEMgy1CF84tBr7p2YMCl+VnUiFgRzWShZAb1L7gV5h8Pgn1MdCzyrH+PVm8ktMv
rO7lQr7wp4GUSPEE4ttplwE7aLjnbSKi5JTMx9yvvVsyGNFfobJtnyOXCva0Xp39
66XUhSMzCaz0BQkGeWmbO4GhTqM3UUI+WwI3Mq9ISKlJZnXMoG+Cr9xffdv8rV6I
k9Ll2BxPkEPBpkrw6eFq5OuQ2RWDWzCNdu3IfOi5qmbYH9vOclzvisv4YBU4vHAD
N5nBLzyTabThXfhUErhfV0scUhgC0UlJRAXFPSBC1lgXFd2tpkotgSjEUrpNciIn
wzXvnhWphsBhIrxQbg1wGmA/F8Q/gPrMPZMhLAuV/gwamZBRpOfHNKcDAoK9cn4W
GIMdtkSnRqvcWa805lNF3r8XaTll2ChW0xJccN+CermuC3IiqrtbAWLgxPOtHUdq
VRbgP50nCv7/AIc5n+RemrQ7QqonMyTlql9Q4+Ln90M74SeY63XdAkEhEboR7gGR
/bFmyVmnUvnSfGuQ68cPt72kq1t1zjue9vQKvQ9Fq2Nu+Oc1KFI9gfZ9jdjniMng
RB3Y1DE+bqWBAe+Rk+ORKK1QJv5alhkh2ywHYaW8xk0KKz38h5rxH1enDgRc6DV6
wAXrBfJqUqGKvyphP2lFfh//2RMu6jemkE08yVb5jcfMyCaC88DJI4HyWS9bO9YR
tDBSGPRA6eV8D2rN5cNNTSDmwyVRbP6FUto8ObcXzGb30qAm1BRc+fJT5GsXxf2c
/0yFoMlwvCKFwqSgOGU53vRhVswyXuv2fiCIEdQlu4uBkENPzqwB8Uq2XHSag3Yc
gTZQaFgwRVlIJK/QFQDQKq8RCZC03kujcdlEORrSMzQ/mghcf7X+LgL99oJI5jnX
heWf8JqN3TT87yYBGVDYZCzLPl6kMjXiyGOncrKbYNYSNXkggQN8Pkt0/gsImqsJ
v90XY/KZfxeNqkQwobmlvS/Y0IYOgIXXTxdRGh/0uX3tD21WQmv6Akxzg9ETstVd
1ixE9lOMxezbx9awB7aHNv7Bsulo+RDEhVxI8tQ6NHnF43eDWeOhgBdV/d58KdJ+
0340aHmOOoa93+S2xmor4ZwEhEmp25VoJGpsmqtApFfXtIOlZOfqHjeSFQd2+JSr
JGVXL1XnQtcja4EoZZf+RQFZYlsbwjeUt6AUud6+bUKGH5mHBIn0+70rq+g1Xtss
biqDw9xdSEoEeAL+X8O/qJPVk7GOdPcj43tlkpKrBUOvTNxZ/vaDOdo2+CuwlkfU
5IIuwssp1WpTTCZSTrSNlRs2tGKOZJt0O0xyTUWJD0ok+YSIgBEZdXDD8FtlgD4Y
DAkVZIAu7qIQJRok3uYVe7SgonPyLKjlItwGu3vn701fXJt1yN12rvq23lI5+Az+
/ocnkmHy8Er4BK5YzMDg1SJ5EBqpfEo2tCOX3Cvcv3TMVlT2HUjWGbKbUWOYaXJf
7mEq6urr+BQaAKYGN+a3U56qAR7ZqgSgNqzN/wvRn/qNt5VNVoAaoUslepmCZihl
a2ikzgbP0plQwg3HSDTpY4BFuco4nF2y1JnAy+tbGZACBXHULAXuW/RCas59Wrro
fRHggHFKNAUUmXTJilh9QGj4+46sFkg0DZGTH80qUwNFIt/tHUWGgFMH1TYkC2Ji
kB4RoXUpnmvjgz+GLwV5VT6xYiEIqYRsV9ZxWdu39FKenjZxbno7EwQmF1YAtSja
/LgQhDZcZAvm6lfda2tTBwGCWvb9yikcYUO9WDOpuebKbPRmJnD1kb7B9BhpRoSW
N2o4Yr0PWbalAWZrJbuq0Prtu7m7YvzIE0MWIpxVFHxbr8G4F5vTX7CLKBMKM2So
XSpSxu+vTFma3vXVRDsL1H2YBDaNHo1e5vAMPqGZXSCMSVdXSVqTrGr1pG81CQ+Y
inhUby8cF40RzRMlM8G5KFPoVzS4MpAL80KhL78DXj0IRp2ueb/f9EB9dYLpkFOh
dHEsWZz46bwJUPBGzEL0H9Kgch8817eDIeCRPzW7eNnk4FrwaXGrtcpkc8WybSmc
fZU/jiZ8HSgmS1/LZF5rIZXnD+U/CDZqfNXn9hC5qARWMaBt/abmkLxg1vkVOm/a
84fSXpb0epPvC/0DbdLUaY3fhyGN/E+UIfZVJOT3BNV9sQy5pTTiDZ/chyL1mChd
iMt266JE6DuY8+TmLTHzsMn2ypi2tErXBta/7JASkuhYVq7rEjHTFuixSEudBnQt
Ie212Q/39m/IYLVUoD67CBu2Dq3/Rczf8L0AV12RDnbXr4lhzZuzcfVcuIoTR+Q/
3Or/jW5DjCzWj29AXDy79MDXw94/IhGJ+K04hpQ1Uwf/AtEDAq3sZGSvi4rv93TR
xDqFbYySKwtjbrOAq0kyCYMPoHbjYlEAL/VNMYcwi2r9b4vSAsDY3UZSYUbwpQeI
6VRmGrqTlFrVEeIPXJ8I48j8DD0U69QqyyQ5L7bIuTbHDhvOpiRY2vpbKVkel8I3
xWFbPufwNTOXxcVFg2zFShMLdKUAuNSZISIUp1eZWWRU/eQeB961TXfIOoxICNYV
Z9w86rrqERcqs2XV+gOVqssBmSqhexKVAb74EJpJJXpjFMf1QnjIRMEbOvZ1ppNL
eb+gGZ58AfyaJCaMBTuTxrQwTpTKe1SmNcFevqC73/EErgudoBmOHZPPIdxLcaeu
2rGHboUhR+4StOauUk0UDLbeWiYpUxTt8zySyEc1EKa3NHa+7vFEjGpkLsJodmZ0
Xekm+JQBby396+wo9kGRZOFxLBwrBXLrLxl50Nw+BXnovSyqchCx0M9V1wnmM5Ws
Q4lUYKScYoFk7T+HuXDrYlDA/4IXti5jExlOOCAer/Q3Mn2RekcafDUxUGv+f//B
gm3t73GE+UswqrPE+IP2JohPyoeWZNWUi0fLJBUU1vMvnRBnfz9oirh2on0YxJvq
9eD07Tka9ZXBflqByYM9rUo0aY6YPo8ptG/Yp+BGFwA9WkVeSm6zbNajminby/Yc
zu0yABcZ4LhlGAyIaKvXOEhqAWpCycIA4Jt7v5P7vjiW48dtEJ7sps+9qZsE5qCd
L4eUpf7ulFjylH+7HuVdR5vHc4S3xE797kSVHtfkYndTFoVw+jV6uUy+ypeWMDd6
ZF8HNqF45qZQd2wZccflxB8M1X8MEHlG6Q78id/AbTEVKd5aonL9aOYszd07zChM
TQgfP85SDO4oNgyBAzdpamezCe2X6ifZyFDw9Qb2sx3sTiHlE7pHcwLY3pRPm1od
29fYyyv8RsAk+pc1CvfQHWwJAVs9aW4/jVi0UkWTOYO3eCyJd/hS7CG5K9FAMD86
QrF2QUJDs4Y5cznSCvzwxs/Wzje9ESrLFIqczIUm9BDV4H31OD5F5pLhvPgesUAi
IMeW7Ba3aTYurcTCKzM+W1baiKgyHmHohE4TF5FrnbK4Vj2wpPy53G/VpDcONFFT
JQFlJtJuoBet0plTosluBaw+p8ABRoR6Eebs79400PWWltesPQm6tJRtCQO9NEYT
k83ZcZaKeuzRyZL8gOg/smP9cv2vrVaOJw3VTlPgqNgfbGdN1duPdrGaILYA3s14
7OZa+4vLqwmluPRIupiSmfoKyEm+cPsrod6Em81PecUM6MrPrWvmEhMUb1/A+WTv
LhgkixLDLNQwwiW5XjoKG2k1ztoLb+n3boMZ+ZalOJ/UqUeozdGgNVgs+OuY83J/
hlfzvdMVCszOrazpBN8S8rYpdun2bi92sbwaKfZcDBICjLly4iYx8Nrjmm5JLNB1
KhwjOK5LszFWjTCGREfP83Vb5vA+rGz/bHTUsVi4Tvg8nC6ifsD1UmbzKOwNS/x6
3J1H3O5A1ajwelYiU2TluLF1bV30ZGe6bdYHSaOcsDyjfzqsEj6ODZsbeVCQVDA8
yqgnF3rPzDz99ux+8TLzC385v6T7GY/vwuAgeGIKLmxouLKZx+mMFwatsXHAzqd/
SEwJvcd1N+Cf90IKrSo6io1AC7QzSXB/Fkhvx+SbUAmuDBXWeKIsQc0t3ijrNBTQ
fVS/TIxCNN9S321PWVojIsmV9qBTBh/TggNSDZufeRUioKuPS4ctrj4zA9fm8L20
qqUukQWYyFCckIm//0RmYXCQoT2zs6BHY58r1AmWC0huAaWhYWTv4N1VCAQiB9+A
M5oxnGikzVArGHztSVVJ9IxChugHYxfNm3opWUwLyFTix5wbkgizXwRyovIL97NT
mOkTO/o0jj5b/A0l36735kphpyOIZBEE6dvIUF1f/zO9koVv78VxPq4moqlNozDG
uadxE2mYvcEOWx9nuwpm+lS69e4Z+Cu0jxXBlwzU1NTHohTACdSXIwRkgMOGPhFB
XHClg8lhd07YLKIAHp+f8E+JWu0yTwKjq2++5/8rrYbRbqxPOnCjYrm4t79MUbZm
1BBfWDv+Rcxtk+nSTG6iIAjHbcAinzOUIHPFnvAd3mNeig1gXg+Rya8V0KGD7Eob
/GNL6uv0Fv3VpaX5sDnzMwrx/kvkpz8KI1kf+YerKRCqv6HH+Rp74fFFLOca1i5Q
6O4uPn7lc772u+X8XzKmtA3/VqMWXrTnnAnBNBjpsQPFNHnwkd5k820KZtF+xmoK
5OEx5V5b6HtKo6PQ+qvRTrhkppFkWjy4Mq2w/xKEY9dYLqFhZZOny43edtf2tR7s
GbO4BpmrUe5ojmBjxQRLA00XmuyNUL4qcGql+2Pl5KGv4vVoObaCZi/n+A+B6xbC
Az1NhPxCvf1FkJGwt33N6PznRL16PlYlBTihiSPFr5uaNg+kXJ0YHHQtvjTTt6i5
KaE48sAOTkwSFgB+QMWqzYOcurTV8uhKuWcnTTZt32cdo3juHAO8r7F2MY0DpapU
VcI6zmyZ/wOZHTnE/FgSsDdRQXTny2HqI944AP0gVE5TDWOaDUh5ExDJlQLxa7rB
3pS3xVbFEIFHE7wuSdGlFHdKJDfgBM218Hlp1T1MaqwYgXEtPJ/g0WVZlcu2L934
NPW/Ulu+iyNG9nxoo1mn66wo+dq1tRBGsjhDvzDT8PSim25oLDxXBRZ40kN5YMc0
AyAn1Jyro0u7YQ4HYBAag8zmstSKUv2H5d6qI0atQ0ICmteAORKuyCXNeukQWoF+
CSIIfpU/6rq8+iijT8HhBLyVZXtJcZqfVnqK3OOYkuJbY7R5pqNC89JHuvPd+TbK
+nYsKoi/JhH5xjQc+Esr2ZZMFRIARLSJF3VV69/4oip7Ig0gtl4TdzXhvGgJ96vQ
yzMW35/2hyIbGSWYurlHbHlnE6+sEz8M+jn3fL+tNP41pC+R7fquwtD037sukGiS
i7TOnSm2FJW8Qn/NALE4+uDNk7iu8UeY7k1Dj7/todYQWe+mhzAwVKstIDa0kLk2
xDLgv9h/vgq/f141gbZQzxaWtXyllVXn9d0O/SvTQ8LF/9NuEBoLY9XZFl40PE39
fs7U1KAHL7cYpkpVT8F4JWyA9qz0r+5GeiO9aXuILFmI2XpLp5zLxI7YdYaWxk01
MloOnDbkbENqJOfb8VUpXbjXZQePUgQwk40N6NUj0Vj8nbR37RRo9/+xIgNRYdU4
54+ClcSVED8E9G481Z242GKeYX8OEb7bYnCvfE1FquuSV02eHGWsuPXhRrvRgX6d
SfUvAtQWMMdrAebLO5BaxK9gMhBYFGs7VlFLCpN8w+CuT7En+jChaBMYNhge2Dvr
z1n1L890KyU1INcke2buk68MDdI7Cg54HFnJSkZ6XwD6+FYxAV+FqBTJIxrAiUOl
RCxX/DUMhuFrpdY0Qc/x4ajxllnTf1cljsueACNLAPkuzOxagj35Znc0oFrREOwg
1lUIlVRFJAAp91Pg2NGVsNb2BjQ8HdG3A4Ndcf/TiFpchUe3qao84tKCp9MCutFU
LQEWJC/JefyRDT06S5hp46aE40CAw+xGkC6aPQfUUgrgLHvYIgpRnlxS3wKnsYtm
oqfyg+cqQuitsWCwa1dDgPJ4lHGKzL9fSAcKV0nUflSoqnyHJZkF615JKBRh50xy
F1cWHoJp42rjk09WDC0nr8fyfxPtgbu0I/rMGf7WTav8CJtwNuLGsMjGYwK6TYSV
4TW6wum+rbm+YyZ0aKDJcbYqldf/Nl7CDfH8TxtL+WMg8tivG5TXyC/x98jPhX4J
vdp+9FrluJgigBxL51RR+BEH9dQkE8oYph0c7ygmU326ZZ55tSUAe9pDbO7Fra/j
WZyIGOEEeU0ic/OEqreXcY0ntjyvPs0xeZ8PeJNYgYCijcvM54dS6TVJhcq1lj0s
4G1zxG6QCb5uTLM6R3ZOaQ/sSwIrtCJIhn8/5HD2KEOeerrAh6+haalAmFDF/jWp
Dm1Nb2lqQgrB9tzXB5aRTPfnFwd7XtccBv6CJsxvgrfmySMomyctfuoO6/iHmdFK
YcuURN3wdKqe6iHcXrEIg9WE9CevFfQU6zR/l3il+x1kVdB/VAYXCjvlsyiwtuAo
RgTcYXRLK3v8cYYsnYZVj9KTF8ltGDanO7eIcUXC4WFK1sfeGiSau70WGylRrVrk
5pzCMgrlkLU1qduVPYHawHDG3Esu8Yi1RkOWMyKhRJ+4JNOslgvcSL8/jsxEr7TY
QbeZIhGXwsXk7KSfQ0JVRkkHBnejtuRhQgmMc75zOXk8+WXF0Jm08XswRgl23QGk
ctjfEPc4t9q0Sx1wbVTZ99j9+ZzUfKkxDavA0M3d6CzBCq9LstqtXZ4CElPqFLR6
FMy/vJU7qQ0Z7nA1iXzISmsejHiEp9KN1wPGbWElTUikHJ2QzV16qqEYh5lELPRk
HIxI4LGstdBzyoGokmuH7xaAlHVO4Q2RuyMsccQ4aqgrM+v7Ll2CENQAq5MSgkQ8
IsgyJkb5l2hBO7K5qgaEfI3mNhI3T4Z5eIwGsFpbZnNEAmwqGLTRBB5rxesSJYdJ
K7zuBNZSnoY/Iubwnh6A/KzUm3owVwxjfWYJtdcEZRnpMjLdr/HqNTmgsizKmdJk
jpeFCrpDLdv91QzETw70oyAcZn/x2YIrIegCekv7U5tsQpFTjP21spkSl+a3w1MC
tyvW50+U/kOVwmz3xyfH50WDUYKqenSn2mFw0mOpEgg2iSpVqzQzWEgXiD2D8Fjx
I/NF86gOvUwLls1K9n7Reu2jK8Ug/fO5m93Rlc7fz3Tj9VDhwz3qpCuJ8XuLgwMw
xcFIEukSrxd/d8JlGtUbAO1YLGUQ6FSuzQNAdglgQd5IoO0qwDThuhMTVBZw+tRr
mp3PRBLTaHY0bp6FmWknJtx5/gD/1PZAMVgSgCdgdQqUBLyVg/ggYLSYxWuSRzoi
jHbfScrceqAPqq9WT6+7LdLQDm93GfoEnUoYl9VfzKu36GPnBuq7s3SdXD94tLUi
Oxz7AU9RwY7XfXsQdvtZsxsUA4qYKbtB2Bjy5+qMDnxBnyCnh21oAgYPYepLJpu+
gfzYb3iDjfpHevdo+kU8DK+LK5yGYFtaYVnjJZ8b+zZ9YtEX0m1hpStv8Y+gmCQ4
tcGS2MOjU+QzBgMNqmAqTrB/l+uMxYv8ekXrro+xizoFqXne1WScSY8JBbN1LE3r
KmJMoDqDWG2r/LrxYU8s3RygDrvctjyD8EDoudgkfb5zTuaKQ0sr6TCAGSc4ARSj
s62bCEwYsFSrR0F+DxNxRmPUbuRjs9qjxF42PtWmgjdKGF+NgNV9pBOpRYu0V/wE
gKHrfCoCTjT12OeugdAMjjxSdW6dlmTLjiJ4OZ5FRRe8ZuriF87uZMFTP2Wp7B7n
bErHOhF6mEhikB7UwGNvhwDhdhjCqDNalSMD5P1TJQdZ7aXiCUr7BWqphWtVume+
WNPwDUNLipqZcI3KQlTYgQfu9+adCmV5MffA1kyx8crHAHpEEsofGlZIdBCv6uze
bhcRAxNowHojeR8dE1XsVV/X180xjnSh2w+j4Jc5MvxCpO3mirbz/7HVaLK44Ge0
rInkZdGL1lVWheHKULlZSCh7i5IRBZen07jCAcAW/Ol8aZboUpvElasd7LwZCwh9
oDKDmA6MQD9SWV5peYcqdtVTeCtjjGW2TPTG1vjTPTbXkjeer8lV8RqSubLrNWCN
bnW6RbK3/iMo0zoonenq5D217lPUGNAnGZcx4DzpF3DFHKo3Q+6l3PJnYl7wXsf9
NGK8i0FdA6JtIU9+kkcy7UAy9Teocc2UF0g7lc73hXYS/mmqSNQNVMVUNvUXk4Me
DCbKeWYPyS7Ij0ySGKBIXj9EL/zBnBX7x1ew1z6f3feQdmtj+YY8PIjuJDT2TTya
mt989ITat5ioAk8n9xoh3VArf82EeByEeOCWdyFrjfCfhpOxEpdwRE71bCykmO+G
j+ro0o77cO/dYd++66HV91dEXbZudz22NHzWbwFwuBlZ6ErBshKUXg1uuK/ZlVzU
FbGnlooK5u8hsT5ZjSbFOHsx/o5vGRTquhLwQBXQbeec4EupPHGG+/qVPK6ULHav
AS09RIVcOY7clqp/rEGe9pZ72rcPZxUM2cE6sy2+r/JxH78x7Zomcia3K2w3ltI5
wlsD5Ir5iQy74wRlxv5trA9Gv1cPOuDxX2DnR+i6PrXZ6ksdXCCrbQcnnfG4gZIi
wMK7jytsDBQbT5IZ1DfQX/rqiXjno56d+KdgCSW5eOolMocYoaDAhUVFY4e2j86D
waRB9sskcvoPJW7WoTxmmiiecOMdXJu/78gvJKsWKcEpvX85/4piQg+mFJRgsZwT
fSnKFBIunF1r0D8t5+m1qEmNYuDOiDgPpci36dROQl1yN8sio5ivNmhjxsVYsbjg
2tkiho8USkjChE33OMYoNN6Knz/HS/n4CcZGvLjpTzjRg67GNgAxYDLGHvCDTkkY
jlFEtu743XLSd1Yb0F9OMPLWQi46+kgnFUvLw5Ftke/Viy0FJoZyeDQIUq/0PHe2
vnfyPmKm48s8f1n6hIAsnW6qGvYCzhqFxZjahGgWK5YVa3DEI15wrtSYSyPnsg7G
w9S8bkuqzzdlESG84i6ac81VHm/0+ivcjKdUf5AQ8Zo0Oh5TQ9TIM0uF19PcYJ79
k92uhxK8J6Iqb9yliIsJA3pxrSHlPjDpccVGja5ikNTAbEeVGkGMdWhDPPFSlakw
pNQ0eVjWpMVp4rGx/r2nW6ADCdkZQB7oreVCCC2ZS6kF7BIIAVGF55VepkHF7//i
EdnGMBFVssqGidxsRYHXaR5yNJdIGhrT2U/koMPlbLW3VdEYNMVTHS6lrO4O8UsL
pK5lAbmFhYDP807gKgj8YMuyDPxNLI3JXcTymp/TyhOSe5kL74m58jPqIRuqKuKK
/vjq8/1+khfw48PIIEr7CE38qV0nWzWcP40sj83imDq1pkGxPpHFjIEsxfQDRbEW
ZHOfVgOwofeRSI4J84631yAbHP5TS2wq2fWDAskZQXCHX1jLz4SzAAIMvBIKW11A
MiSud0nxwW84vHORVcDcdjFKblzKnDKRSUJZwSdclzyBvdTjWLqYJraN1xhh1rM4
DOqwmq5oZSC08blxF3b1f+4q9dqjXBBOoasQImUVdV4OcyM0GJkfdOwNCo6hU/4U
tccyCIJOAlEA/5ejy34+2n4HYJCXBje975un7HD40G6tNY1A8J8xtf4DhscMkEjd
mqdpSDdFAvPQSMF6tIDs5iZjK2JbfiARDktznmyVk95rT4WDX9MMgTZuy7MheEQ9
imGtqV/Ni7RoakUNjQt9zSGsUdje7DG1/Sp+R546wX9hJTnjrkKbSUZNNMQHDTv7
ccrImcr17p3+fcguwnjaUaVlY4Nl5KohrWNB2PgNwcv/esbsERbGIHVRNvqGnW/f
YQQJuSrwg2dMvxOWZHEkRewUzLT+WTn30ZSjsHS8KaTnmXt94t4ZheNjSQ/vstD5
DFKg7u6jan+1FyK0Xq86URC1NIskt968kJPeEwDlG2xs5yJtqQLcqyXHeRKz2UQc
WsJm4V27dAJAPbpw8yTQ4Ax2Zj9aaDrjfs+zImriUo3tRGiBiQxDDKPhsiCT7sbt
aycFdx/YnOBxJfzDboKZ3aJKHoUx3eyVcMD5X9lrLuCz406Zi8mhOh30sLG57hd+
lHMwqruA9KH5BP6Asc/IWvllmW+/yVMxyNskNdUlbLZlQc0IpJ1CAvzCNpC7J4zf
dOz95WxwPCD/M5FZG4MMXcmjOgI1dMD4zhheEDKwehuWwzpRP/VePi8+0e0VKAQW
jQKiWWYXBKFn1esuJAP8vuiA37F9YXWWkRiuuItitTcZ8w2f8LyO6GMzcZ9GmCZf
LiBWM2ZBQagh/gPhO1KFqsWd4kSVXhve6b2koHAGG9dfKaAQE12zxN3K3yqXwNAz
btgjewAVSPZijZ0yy+m8JtPWUijdgTiw7XJC6BelJSQmAlxiJDFfXTar3OfOZO1I
G/g3ziMuJVu3qmqpGhsmRO6t2ajXe03GRico4QwWmSevLfKOPvJaoVV8Br62w/7a
THDOEWiyy+zuuniVXB9qPvO7d0qLv2mvhmq4VKWYnfJ3SI74fMQmBPHKFQ9AHHms
CHvry30TwsSgtD63vNKFetw6lMvpnAybwp3PjfWYSp8BQ0e09FpQGAlsGnMonZDL
c1yaMINfkkwW4OQssXGiJXNaF2y7kKKxDD24F50aSam3Rj1UcRW9+DZkBH55NF6i
0LZjIMhBFUADnRrOpsFP63sIOB0HfngZweVdTfqiEbCjAbDNeIemvj4/JR165ewU
YI//nCT16bgp3aSps2VGCnWvIB9U8OtLPgMUu9GzBDA9vWnB97ao08a1ZxDrkEs4
kpk2YAF6/qutWXe/pQvQ98T3mPCCfZkFYjkVF4X+4SKb0nA6FrUO7y7yjkNI8qO8
Sxu4fmku21galIPMvIMe5S1jv95pRJ/TZA3mH70YbcqQUynOhu1nApQ+z9LOlmT/
4xo919usdvgBz/5awY1oyjuBlMpjznPDQWo2/M3+AEcI+s7ftgr++/OUa3x8aIl3
cPeFHRWtti8JceXVApivr9tEBI0g33oGWI6sK3FjGe8=
`pragma protect end_protected
