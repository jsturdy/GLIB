// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h1VYcNFN+wHgYAq35dFeSVs3x/Rb6T7EGa6Qmx4JULHC7jxnhjZ5nyGH93m89g9F
7nI2ViZvg/SwLsezhhvqF+NgDq/fhTfa4DZnyWSUzLe67M7g85XbXUgzfsUh6L95
3atnMKSxmkc2lozGsfPgP+egApgXLDKGyjmR5xV4aeY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 125888)
WWIgrRLjgk2dYFoPcpDmyiPEk1kRaeiznOhDLm9VYlzzcDXnJTYSyQi9g8ZxLpCk
YDlIQm1YNaCyH94U8MIj5N3MHEWxSF0kpNiFMAjK8MBjjMFtZFA1vDtWJLvw+xZH
09gvVSTaCA2/0FivyLPZiTo2YeTGS/gKWI+UjMGVZdYWjH5V2/D+IVSUK0ceBdfr
e4vehe826e0+Cr2eD0n+2RBsQBKT5jigB9pYXPONie766sVqrbsqy4vjRcJpdVhX
FowGgoNAUpFyRvIqK4auV0ixDy2HK3noq7MlEZDOjflM+/fCt055OXEpq+UeF4Yq
OWX1tHCIJ+LyBugQa9ykxs54o/csekY703/H5bctCLyvkqJRD9zCsuwItEaenbQe
oCovpIX3oIlIphFGZ4ES6KEb3yg6PaRd/DjoFTtoVlZiQQiZwaSr9kc3NADSAzi4
Orf9qHQv1M4b3cPdzQyI4k4EQS10i1OimdeWT3KvAuC6s7OLRsI5/n9J8o3muIBx
Mi1syMBrCuP4hyljUIYGkAwQROMePK40zoLTyfd+jWDFDzgWjs9Mb5fCjXMUT+t7
Pp1NsQRY/gzRZxfaMbsQ/0DPRSotPo9KoSf1/0Kqrm27whyw9mOeMRPM7Nxz4i3l
FtzwcoYGG50cAKk7mGpRiaIImoQL0ibPKjt4nYFdoDpPPDEBeeOhQfgQ1ur0WjXq
Xjn1Gog9fVhdoiQhi99UPUJHRdcgLvqmosUXKWEeApLEZoxJthVLIQXS4GWCscEy
JUBVHy6CkXUGd/fprJyu4MZddxtloRhiEV2ljEJs+jCCtBSPEgrsCsECGPNlq71e
tPRcqkz0XjK2U2vurgh6I4yc+0CA2B9kiCUcEqoN5TTepLhSe5SHLSgI3QGnJzeM
13W5VdMa7aY0AmOeIVRSOscU8z5eAxbzOe7W9uSOfAuBusnAkb2gnc0PprrXEqqn
cGvmn1a/BgCTXL67AOty+JPYfUD6jVSp1aWy35pi9vbd/7Rb+6Oj7H+FvpjiLu6m
cQyKLoEGubBcnDxgVn0Dk5o5+PaW4aN+GFHgWndeb4X8RnQ3IVIdT1+4jEJMWRM5
RfkfCwQ2nxgTVgJ7X6FWugRQGSX+S3OdvD1JfC+PpPv7Ic8V0kc5uHsl09JAyDi8
/Rm7fM0UFpq362gLBGQW3lQ+hdreHs1yDyzK6z37wi8onjKnkyhao1XJR5/9GtX1
2MmuFKt3LXlX7MMvGCrx8nmQ7qTAGhpAUBbbu+FDCvFXXfqYp5jnRhDbSWuvxOPr
iJwIJv00Pwn89dbVUUMgUEMMkUdyw8w6JlrTJzd0Y5tRdeB13nzTemXpxx2CWSBd
FCx8wmYfzEwmvSQFx6kg4UBKfeHNO8YKotXy6QtFRazPrBPIM9UaSDVNpRYOjXry
w0GxZX8huNbwTqstluvhjbMHLo5ENwM98TjfG0FGQyLgYT7RQmVBqlk0RAJePFjH
7XXstjdVskEAqY6dDRe61Y56fbYEoBy8r8VNrW3RxNVH2lbJTUMfNKWzf6zXva2c
upFtUGamZuxbKicIaBcNZy+ATD/kJj4sX+42+WkjxVqJD9A06EMiTM8KoQsZUsYk
nzgMKXy5waXHdR1YP+tlFHE6AqBesYC3w4C8RrrKphCUeckFzqQUNZTjfIXbXotx
7+MEtGTx2SIR9SM+CSSEeka3lO1q6K9tCMz65f/zuJcLlwxXH8E6N5PJwGwKg2bv
9dPEbjfeA/FEYfW2BgDtV9r5DxcvLD6rFCxcMq6b1/NweXxrCIgdCBwGsinIrJru
fJr0DXck5es0w+sZ0ozvRpIaUeMdudEtW5Cj7FQ1kVXvrr9DjTW5gAMfbTAF9eOZ
cf+J5BUhC46UtzhEUPasMCDyr3DM0dG6fpAgxUmxCSanD5oPks7UvGSlU9uCQX4w
f4Cp+K3McH18FRTNuMA58gQSoadan4KycMVFPZzt+4x+Ov5eFFUJe1nc1bb0pUoA
56Afvk1P1yXA9V4Qoz+sAuIYB4l+IO9xSCoEAMmgAINstg8kdxBkU/jFOuwaqtuE
D0kjwaGD1L/poF7aXgiVcYZ3RwHs8ia7H2wR8n1NlFF/yX6AocqulrSKY3SC1tuj
oeXdQkJKnzUDX7Cw1SBL75ouII+NSxMjTYfdaXj+X8hGd4KfZ/uwTzWtG6fiPvw2
4BJN6/h31YSRrTcEiW/zGV6o2ohTkBq1jNMUKrUR46FkfBcoPJLPmvmTlAxXLzHh
SdTFNO3v9yLChn/HqQnfruXQuPpxcraCi6bgfdbNShoBYV07bUPvFBbzI0tVyQqN
0l0Rnm2hA+Zv94k0IaKmoZWO4L4fCDPWgwvZit8EwAuTB0gvSKhaO4qxlRMoGRQ8
ISyogHk8FMqAfEBSl8XfsqOQ6akRWW1oTnbNavqniFHHcMnpzFoI2HOO1eFSXqb6
IRb6ytFSz9/1W6vYoZ7Sm5Nyz5NgjpYupLpH9u7AuWsWUW+BdCH8SrrrH+8D9utA
hTF0qmvBtDm8wvq8tVyZlD8DFGN0ipIqNKCl82y9eXjCOrYtJdUFxaLC4WAOY49G
ZyYDStv6Jxh5DnV/cRsDZ3+h9aBJtR07k8vgQfPDp9vbmm6iqHs874JlRjKCQK1I
9In7AVKUPnUcfmUZjN/d8GKhMYvdL/X+x/sKH0rBF6KGIyHNLFAkQYL6o4rdlq37
7xZEPPyP6Lm3DDL5m68Cfs+JUXgvBUwyrbmkGr4aulACGABTqpIEflwqhmrgfLKO
WroWCoOzmBP5ETqyP1Fhc7H3vMK27sRL4CS+PTcZLGYs+4mKEJRvEqbUSzMSKJXB
3pSW0TZH7dlWTLDX535OPojPmE1FCXNTv0F5sE6E8p/Hr7+miSdEQXDf3tfJ+0Np
GdvU+et2nsu6RWigwA+3zECzw6YsNegRBVxZFmLzufcXFI777nLpEzN4LaDAp4VX
h8aOGHWKmYjocUhPEwMtHcJIoQiRGpV3IWH3irw0S3sWX3r/xkUVOT8UC8iNsood
c1vylgeanCkTwkQu3SOJG6qkUMEGEdqkYkA0p+csXMqp4ao/l5/suk7P0OLG6Ssx
Il0rMGNrRDScsLXtyU7MTA20hkIPVmkUKyHPH2+TYpZ492mWDLVBagyaciO5Ckng
OGH7OXZhB6JglQzRbbYa+K052OAR3S2O5nYEbc3CZ1PsBy9w8VfFeiEiHNVO0GeX
RK7Q0S8qsRMopSlnxNy1i8HJYnvBH85/WHc/ITcSS4wGbeXGuuVIt8sO5E9SBF1c
OwPXt5MD685k7xaMf4fCmPGLMj57frj36QmH90a8h867asumQHHi02NnYsdDReL/
GqkYRDWoFKysJzegUpL0Tg0h1IzHK/xGikgGJQlyySw51UEeSjIOMhe0uvU0gnIe
9i/fhjD73cNxXHS1EL3Xm6euZTMx1BrIicdOfOfHPVvSrVs9T2257igV9AWjTPiz
TgnkVnLjs2wHEI2eV+MaVVuAXD2LXu6UHTQfiC9wedLqYg07KW1uSkUSzwAu/DVp
ufqdzQDxW5XI4vhh+xFDYNguXwdMlw/LhHOAsb0YngbrtZUnN/5Ech4tIeX6AkDO
wwu9DlHotOZWVDKoj2xDkilBDGnmig5rJSbasn6v4uLJricQzboW0037v60XCIka
vn/KTzxe2O9p6PsL5Ocj3MZ6FkrHhtj8ZIdru1d2HxUjE+Dx7beq0I5oaYYn+3gA
PxrSZzb7DPJiWT9hu+T7H700VEq038cjdY0oJoBf2suLA7Din5mEfqJjj4MHKy3x
vwo5NIvb/OZ45VGhS81dS0oci7zx+n1mjy7v+KCe3BCy8oO0YMnRLE2qiLn+agsm
5Xn9B0wEF0xoU45iRCuWSUhZG5/6ONpxGYpHUmUyAqiJumYB4bKqm8kltwLQZy1z
myF3ZstDtAKEy9+5WtsNdvFFBnQ6FIN9kfROamTZJ1Pw7SW3rQ21KOEUsMxoBx2W
VUcHT47zjz5GijLGpA+hmH2w/AqEHiqukP/tXsY5qCosY22VfAlep7JwrX1hNL27
z7wI4cXWeAryt2RjpL400aA0cfxYo31gO0dXIUyaN9bvN6OyIPNY2t7vYngL486d
k5tB/PNJX4O4l3nviWPgkmCNwI6Gnh3SjoecNb+mStYeqdfq4cLcgYYmqBhAsI9W
qYABlxW1VlHY1UpgjL3JtMwLzy/JTMi0EsIpmMxcqNLTi8Kn4fOXbCj/5F6sbwHC
O2v7E/Yg1EPruY2tLXBYm4H7WhCOJvI6sx02j+ytLOZZ5Ki8mNiPsMivwQlsHXfM
oNVXXJ2i5ESUXOaHGP14lfwj3V/z1xRZDmW7OE2aGPkWAB3sJY5IyCzdEIl57hmi
zmotIMMCl3IdY8ed5BsZqtN9o4WaTT7hqBSS0BnhfDntsrM0y+2yh1dYE8GPNUcZ
oIjAZ4MiKVufjmrHW+vBoVA15OOfXpdOOPUeYi/BHG0SXzfK3o4wCg65EKiz2MBL
iVbEilwubIkqvKMCE4y/hLEU2uBuG/Kz3YcQYLbBZCXh4xZ52FqVpVtxzh7BbkCj
SMiIHdeAg6M3T+xOHZuwxHt7wTJIgraxshZki22CdbWd1UDCac3O43hrbeX7rJ1U
OdqcZrJMXNM8g1nhuS06CjhPi+R7G1YnHl2hfnjDck3J/ed7r/oa3tt+CvJiekht
1GGc7bEeBIQaeiBZ0cXXx106ARUws6AtpqZEvQm3Arcf16Q7tE6JfbS0ZrJEzGuB
gBGcDzytcLQiENleBumeM/USN50FjqbkQHa1qZsqwpvCX6tzC4xMk00JvaoIT4Xh
jUF499PKM6WMfeHVSnj7ypmte/a+rfYzUFPKdfhczdlV3LN/dW3x9UeAlTTChggy
RN6hSLzx1Akq8yRHovtw8ayjiH/33ganj3BKMUHWeJ8OplCqKB8lnVpJEJM7o3lQ
zVUpBBLoKxbfeQ7YkLCrOr84hVN/I32qIBUzA4In2sv/u+NE86IaSKvz9ts5rENb
63Twdql1Px7sbSEPHM5gMo9TWtEYHG/uCOW8fW1wu84ucudH6LQ+dF14BHCtZFP+
ydcS+wLp0VkQ4q6C3X5AhACI4ugjelYbulkP5GQZHe7k6ILYT6eCz5DgiKQJmi31
fc7UQIhixNt27Mmr+sZJ16qTqnZlyJXAU5WhTm7z8w8l1WimYmUA4EZk2IFhQ9SV
VX3I7NO8fbrUnReQEKPILtdR5iA31t4KrsB6SuyzgWY5PPuvI+9Dk9zDOHv7EtV7
UUoMmBsg4a0Hbts9sL1RfAnrG4yRWgdCSXwTok66Xn+c+FYbd+SaAEqjFUMxRINQ
wuJrte4h6dtzts2F9FJEpwH3xbVXQjHtN8lB85lmfKUxikq41K81ag1SJgrXVW8K
fwEsTIzL6cfNbz29MD3tt2XIP5035YutnYD5z1l2L0edeNJCzuT+c5UTL7nkE7Fn
tIp7vqKlUcRWZNzOte/DFbNCSpQOe6uld0qEIAyRLv822beIbP0FYgto8U9GvzOo
OrIbDYfwySntgGPQNZE2jia0js5LTuCu9rFL0O0Vb93B6vKymf1rsJhbDwrqCzyb
2UvYt4XsgED2PZNPCkBjQuDl5j97dDRoSBQkTMHb06I6hl4NWJ+r6hbLX9cUuXOt
4qac0KqR6Fk5/IAX8k1Stgp35tu5T2MZ9jTdaW8RwM85KYQuJzzpR+hGrciWbhQy
gvhMIv+9enuoN21ZYsdHXV1jn0FRaCnJtT6Y708PBPhAJF8ly7GAXc+Nuqbg5CoK
6N6UhtKTT1bloKIlMdQLpGm2qS4Ed5WcNBaVDv8+tKxU6Dnn2DPf/r4QiQ9lZM+c
17BrTiO+9fKKVY42kwBBXlckOyKeB8Mz4jxpUxyGKJg9Y/QdgETBmxhQopgtoMIn
EmbWChlT0meWcXtffequeDD04biwpKCyW/EZ5xRABsve8ZYQYCMOGmF1DsBTm74r
sPanXIGGmhaz0k4NMPbw0gqox42tafkrs+yiWEJbfk4cx5yN/siw8F2WnXWSz/XV
1ZHXVtNFcq7mG2BUvQJMdnPY8IZIqaIrCh/AwXoxvSs3AacLds0gHprFwzYuBufr
kXP5co3Ck0UUZTeU12KHfv2KnUm697HHOH0CkdO+Vi1HeYYhAby+cIEwtIVTGYMC
iR6n5l/tcm9WmVnlDHpUfTo2H6xdFz+olm62Yp0wrgmJfRA8uAi+G5tena3NShvL
TH9YVXWv2VnOgF2grBndfFaFBk7Zyo+HIoVqiUDajXclHagR9RIwB/+Ire3a+GkM
2+n/2K2sKNp4yketDawQBOG4bP0HEI0LI0XTB8XEdvUKLFrjfddaaoiGHrZNRmV5
C5WHlfla88SQKBx9wPXrPpJ+DRlERpI95TdHT6GO+qaj6AL9J78/7ksLCwJmLeqT
FqhRUjzHzlKTnghtQGMHR9Zu5Lt1Vj0NI7qhdx3wIvCuYTmWAc17J5axBLnVL0q2
pCvDUGHr9jL8ZY4POBk5M14jNrwSl43nc7GL/HrTjHdsz70uHeCQxaUe9NS0KTvP
OGbYPV1cPoFRi8PNxnDguKJayk3q67SJr51wdfGK5TB8ZGnr9BgTP+C0APdU8nHV
PGNiius8I2DTFytpoHKucOarrIHCKtU4E78hcKOo6ORGwoBOD68iUVJSpAIRofsj
EGO0t9teXLjiB5A32DV5z80j9Vxm79ieGMJ0wsrMticW/aAJtNosBhpO+n4WwU8S
va8B1mip0vOoJJSk8I/ogiGsVvxI8r8f+E8XymqDXlHzIL31zKWHY/+iahmJD35J
6O5M2SQ5/WuD7UPjL58BcKMvqg+PkTJWxIa1LrsSJG0U83F2kt4x1XjnzuKuJVP4
ftD3Pdmpys8v6VKRzvtKuJfNRp3c1lhabBXcNKwkjFM1uLDU+ofIDnF4njJ7w/gM
Rw3ROeH/ixKG2SRsqpcWdpzmrXN4PZ3lEzsS/6LUW8rQB6WLEmFuG54Rb5d7H0/r
kSfu7RhFMqUFxuxebz6X7osNdjrxGphvo639qTSve8F1mNEXOTCebf0PzWxDvUi8
nGWyOg02ViSaibOZ4q95GyhYP8RVIesr3QoFVxhFBXhIn30ejU04v/rKqgTgUIpt
WHtDNSrVU3vuAFjFwBpWOUSUXXas2YVJOBw6YYUQUxg2GiZeubzQ2HWi1/TrdOwh
FLmsLNErSQeeHmkQSZd52h2xz6Fli0X+gnEguY64YbR9sD3/sZffyRKxCW4mrnQp
5G3aieBQylcFYB+diS9t6c25tiFs3BbqLwk0xOuII9aeW1dNIRXetwuZPEeOiBSs
aOhv4mOePM9POQBs5ucCksi++Ni189MSVz2DXrla5OAkcfy7OvV3h8PsUUTz68O6
qGuP9dn/2NBL3z6GvLGyIjdXuQ6hDDCj7hTKiuMKqBd1hO1XyccW+tG7RmVErcKX
ncaeLnWisvvqTnQQyDJEIwU/D2VXAN3w+h8HQT6j9990ZOyu5AYtdkg+FPtV80o0
wMHQrpyOJau6rN2XMKsN8fDvovYJOK2QWtg4dERs6W9CsZA1Qh73IuXrapaJ8Cy0
snbnKES6VT0Hhnr0b6UxeFiZ9s//ez9gYKYaJZMsIFFcXQGQ7SzN+dIRIUmMPumW
zWEAmnZriRmIWiEsNhHpsFQAJSwC5UysWVSLFatz16C1SrnW9RfRdrilO0AnkKqc
hMBPJQP92CW5x9yVy6PMudKfC4ZeOpty53qLzznvQRblSjGCor5FmXyd/onCMSIp
CST/mi25oUCDG2cmaYunbLItKzpq57hJpy4L8Jdbn+t0rncDgwF9WO94sXmn/A71
ZWLj4ENwvmTiTcrRGjxqzXyAb82zuuM9XCTE8KHQWJH7SYDC1QD4d959uG4sgUMc
qG/hY6WGy0f91PoghHkYmFm+EOlCL7tD49wwIX4v8UuWw2oRJZ9yNXXYYmztWebt
ihKb9Yvu/GAXgteRysteAvYHoZ9eBZu5Szl9Gj2oa/WL0fBXhkPKIrlYTWBIsOC+
1eTNA4S0I7y+55WGuIQ8VDIzcY1UNtqnuYh3TzXG68VoEDaWNxe1rS0M3QZiOjIx
gPl5DOj+hrvvwI1oke93xwAxlioozOir+Me3U+7reUj3mY8XqbF44gE3YE1DFIuo
uamz1i+T8E2ESv64+GXHV8LItxDAWfgg8TxeXWCwox8Fh8R8z4fI9GpU7jtVYS7u
MHJcBw6etEEJoJtor0YboB/uh0ru5n1tdV7a1kYQZKKLGz575vIovdCfGkO4Uv7m
s7DluhuoIxaxcj7na/447xruDUo/5miGqRgIWuW6hzRyihLKxP+At8CUl7qJXZ6q
eYa1o9bdv2a8nBdRfrooOae6Sje+bL00ixpKnHW+72iOJncOVHg5g7dUvkc4hHEB
lW658nukgP0xJAQEY5ioRhde8icPT71e7eTn3WT0hx7wfCAAyKjVhtGruX0gdjLR
YraZYbfOTu7+/9775fL5h3tQmqaaVyXu7Ch9EE1GQhoNEyu267II0TF5rWRKlwf3
XqVYhmUscWCpMFx6RhS9T0pCeL55uSyJRBlks/5yTeDMzwGJqZxjrp4zLlxDw2w8
cMu3pg4iXycmmkDqzZFTJRnowkX8PB7BLcbqHG81pxfs9s0fnvQzEMaVx5MgASwz
lEI1t1eshTw1yGhhlMzdUNGp8iBJJhqBR2NgsQ28HbRW+b5KSSaO7GqmxStztNMk
KIX0brMTexO7CbGGmcGC3QQkNh3gf3fYwCZozmyXEe3mSUdL8Ly8Qm0BH5/H2J+B
B6PalyeO5Th7kxc8N4yTPB3hLD7Xg4AMH9C0qUzrchc1bewi4176DC5Ksms3Xns4
UqG6n4eJ3BcwMk2CRYzKofGh30SV04ZtqXaIGYNCLZnaZTVGNo684XauOo6JYnp+
/wvLGyT7OTGDwNx/y4uC2tLlXZBTKcZwhCRyulJn+twWNYp8L4sZTN8bgp1FWwRi
NUQo8U+OmQa6ELzgJlFtdHZx//cv8XtwlwnySvQCfNOraP1pm1uOtcGeEuQh7nic
CfQD5dB89Gq7UAiWnO23gqxuF4dvppJMi/3s52L8szONNlSXd5w2RL+BB6mfPYjn
AsMM8xvAWzcG2wLSeL6Fdg2vzxeBk1OD/gRTsWe11yImpnacm6blR4JvHmu7Ptwj
eznLU7U8RGEreifO5SY86eCR6v7/wLEVahOqQS9Kd7SkQr+uicigszwlf+Ps/iH4
5DJYd/HEtzHXSMg8gXKoHCf16IxZtXl97wA8zYzDlYQmlQVif2wA96U+dcG35odo
dc1AavLIFSwz1oizqyQaVvGr9jAgUHJaYdCnLAInMUG7MBr5DO6InBu10aKJRZes
0uHTBsqX98Fts8/Pqyf8djSXJsq/oN7CFL/4c0m60oNVoWcSMvqThbxBQZYhjVia
WWGHD0ox6aXDZCR9kB8ffKguHkBzPkrOhAw6+1nk8vYDTAW41QOlQC7W2qOk1OBO
bQE/bKyESkEtYJa29w2B4z85p3+92W8apRXtXfem0v8Sl4rBGwfCx7B4NFYgkJoL
yRsZAcUTnCiwuPvE58pJJbDFPD0vk5a1Uhx0Dn993ogGNdJOsdJKnnDen2HFb5zi
t6f9cZgyBlHwtb/oO620ijNVYNFEQo+7U/pDHphH8FPUItadbI1n+ydS1IE7KJGD
zlCHG2jxTaK82W/jPDxBbyzWtDGJzd6RcOq5wbW0DX1BiNLnCZ5Q95D2/ATjuEg3
H2Rvr2WC3XYYFotPtAX42Z1F9bcnQZvPT1yobqiHD7GLhhaO4YVX5aZKDLk5N59f
dvdMxWDjCsMmtmb3rp7snPBmR4J7EvBvn89dK9fBsx2SBwH/omM369rWis5fGkJc
yYitybt13igXEw3dlp2qXQEa0r1gJpUkAZ/jeeWU1JoAZWTYDi3DY+BFmzJnttwY
xBl1Z23SR46LD0selbZv6GFStzsGh3BahS7QCXVvKSfVcg8ewGAfaA1hsTxx6IAT
NIJnKNIOFcPyrbYFEYwMNHjE0dLXPgZ0fcPux3n5quQdDSTghk4HEolo4bpNVR+P
ErjUrGpPAhjYAcfD0wQfUmAdc1tkmuhzisZANRg899JVUZPPbE4bM4G2ZrSz5dl4
fZETjHwiBNwcFGY2z9t5ZFN75Wf77YtgZ7zUg/iJvMqi+4oNuahL5GLrropAfcJk
+AuRMdJdMWnGPPbJizTqmyAxCCWBQdx0P4dq0YbnHxG15T1YdSK1rYhZ47kO8Di5
zgX0tnuBTIupGx2ykvVyEZf9HgabX6UPmGE0vNQPlxKfy8IdzNFYYjefPE05LF5i
6mFK8Bg7r8Ky24LEaM2EF9dtQoTHEUNVXjCaRf6iFavPQuWAECY1WbjFu8zes+2V
H49DQn/qb5TE2V2Qgr/8sd4a3YoR3IPfLUPDoEMxPB2eRglI9Ecpg4ednRVuDeNI
ds3vcoiDabMGvVLFLgw076pPO1y5TW5O8u6LOaEiIVLkGoCYo98w3ABko1f1KoiW
l9eDetbF98TOYtu4O2pnJCGgIPXDRXY6PRGC/82AjxmCrxrXkiIrIXdzDLiIFvsr
K+Be8BifJGBWXLQpoaj7v31mqHYotpw4vdWyYExfPzf/PGLBeuWpANcATWU7L4S0
OU4AFKMYSbLiclz2hax/L2gguBugnBOecmQxhSgY+ciShImdp6JXX/1MAQJx3MIe
OVHWEUgwCkD+GTU/QcVIcTQ+G1jinP7nfuBaHHXTQpVykqcpTQoBtgtDnE+2lDJq
0bRR4RfbHGCKNL8dLmM21ls7VLo9NofnRExLVdGsQg2baFrRUwI/IM46bBAfx0iQ
U1gA7hTKLlOwhwtFA+Xe4j7W9rS9SoCrVnJXDCIehGescTQVX3B7ZdvBhB5wW5Z4
DEs3cbiVgA6RaOYRxXE7hVRtQUHpV+RQxODoXjUhcPiHHnsKuTZppxbJazIp5sri
Ntp7q+WACcnQFZVladF/Oo1tkj19B+l0byentkqIhdnIkJcBVSUwzyhXGEPgpVMl
kaXPTE3SlSaiX+8ZPuLeTg8j6p+wwStaDSX+RZ5w5/bhu8jjVV5MUmh2CQf4O5FX
akJ+OZBbiuZuWqoiB4xRA1edASi1GryBhY9MuhuH5181L5gRn7qf4I0ZC567n5gR
8894ypdYfU2gl4qBEfpNSz4G2RbmwvS1x98RXV52zaoNnhZWoxfd5r5ay8sYh+J4
SUUg1UDl8VszwRoMP3xng3X+A646uYSipbBsxZcxuNHQ5O78qYpK2gNDBi4nP7Pl
+aNa+H5LjzJYVtDZjNLZpwX2+D34JxB+jNJ7IJ+8J9FCi8dEdF79vORmnyoujBOt
BHXcbK/WEGnU1VSW4+MnxKlin+uhl/7Y0zCQg/iTrUidGpOtbxBt0vW5GHoOAp8b
EbLUPChfjE2XxrEhGfBwHaUuci/NweqNvu0YVEhdSVQK3JVClVVa3kma8IyzJL+g
aO/6ECLW0VFPdYX7pFDfqJdslajbNm28s3wfT8h+mKWAThDXvt/bAMQMSFKeDqbA
ecrhwNzRmX/nX0RqCIG+uw0vz0v9NlA/C1US/WzRlH5Mzz8TkN3ZpPLHgBue9pFc
x6C8gqU83tB2r/LnDTRZNWDiSAoCjs3MRkmq6mvWQqNxMKgIMMoLyd4lFtyoytxW
T09c68L4GwZApfJbunH4zQ6xWF0UAnq8zT84lqojypnvZKWvQYWFcInt2pHGOh/E
fHTOpVS1CedPEb8LzgWUw8nOTfnUPfOVheTTx/GCeepApBntXuqOT+T/s7OP4ogv
3+VD0mbzvFkuT2SetCZp3Hcl0ObW9D7W78hcI2k0n2aMZZBNa8LHfKC5xsC9AALG
bNlLqgjMDQg5fgxoLQximiFqtowBb9E0PUovQZIljh01rYkPk2PTCwKDFHsyHI5B
IYSoHOth1fKfGh9a0asFSr8qHRrkwkbVKLBRwCJbUh7i13gQsSTQPxew5WEdwr8X
RX6x13Eg1IgDxj1EMN2nFPsSaNfjOpZftIj/9V0slnbfbm8twXPFJ0KbJgkvcwi/
JZ7+RYGQgqHiazH5WygOP3BwXHY2MYTucrk3k+KtvexTR/GYS0ibL0HBTvTqzPSL
ZAlmhH5SDQuQSPMeDw2wplzzcW/kYjlV0Sh8ahVt6xnIv6NOjCAAp9UwN9AGOoAP
oAjsJTcG738KqiyQbLPzwg3PCOLi5ky40vVFuaVMgUNjXPBPaq5Q69wBWVXGsGEY
og7WZrK/60oqGH1Go2ub84TOzGtnHcCMt9FkvdO08fMUaMerXcvCAVV+MK4/BrVQ
MRawcQA8wzf/52UHMzlryvwH3EFSo9osP2oXFPzyc6YcZ6kkaxNB6qyl7+HJRRXe
kL0dNYtTviONpmKG+8Mrx0Yla48meMxEe5LLikrZdKxwK2oiU+SPVa/WSQQzwdgl
FavEQjpjnFnRyAZ1w3AgRHbnSx+vnRdKL5yL5eCCrx7RAK0dzP2vnBH9X58Zv+Do
uDRw2hiXWqAdWXLNxaf2Vu7LnftZL6PxICXZ0NAXl0jPUqMDvFhn6RFU+p74adg7
rHV5zS5uwLO3vLl5Bpjg3NYErHdWtY2joabdKqhFoTCjKL+AJbd3peA+ze77ivPa
/Ednq5vYDQeE5JliEkt806M/hs6dgIHZgfgtu1EDI3MRYbOwBNrgiXAtsobAGfc/
Gm9epiZrPoIuc8VeCVuWVK5CZEodFXqJaN7tTH6ww0Yxwz369EPUvgI7hbopYiIU
YnigLEQ2Wsb/7kt1DQqAJnXJ111Hvh45bTDtL3pL0of5TQvc9wisWoGuRV7ol46x
oDryk+4rZoFBN6HzpGS7eUYtd0uvmPCaZUb1FV74LfX6+6Mv1L6C8f0136LmD4/U
BTaEpaGYfrI4FXcoxvTMeA/Z/pBC2+SrtZ841YG1FV/FA6yq7pp/hodNJzbqNJkn
Vvhj5DYdwWApj/9UHpz4AC1uDvyCe/jdYYos1xeibEhcKiaa4RLupWyO9K8H8CGM
Q8lGprI6G3qnRUwFGiI3KIAWx2JUfHdVh4yf5H3dO3pXnIHL89Rka7ZLWqa6i14r
oIkaBddvoC+T0y16Zf0IV9rFUgDxTv/6xA68HHO7oMLSqFXlNpBwuHTxhnXnO0bj
hKoy94tXkzTiFjUglqUAwGeSTGfnf/4EaWiSnbG1MIACAaaPvwQueDv+xd6NXFQa
0Bc1Gp6Ueh9FcAfGXfrUhCTZgs0L8mUGHIkHO2OZ3YhlQIK8GuduvCRWKCJOKJTk
MMGI8K6DLwcMdopw9Ubz47KUULV9bXlZ0GwULogXzlN+ZjwMQVglk3z15NZymFTL
GzERmwO4YdEveW0UJWoz5Z0udrK/J4pBbyUIrYbvWP4QEsRmw6zMw1omMnNp8xxI
NDDgjAMcs/FmXTabKV9+YpLrLYWweyxwSGH7PFXrCt+OvdntaCxoyvGJXz15VJJw
SDzuz7/CifKLO1KPhKnDmUbmrIS1lcTvUHxkcjD8If+IV+BvR1tKKBCG93OXlyg4
+trCMUOf0S18FNGU8wZ5x20pIOELbG1CrwwQwPwOd3R/qsz4pRXfsYKESJq80SH+
sg/oJSsH86ImAA5eYvpYhdbastwhW480xK6XnP3IhbFCVrX7tiNjKidjA1mqxkAv
nIOCPAulKTCVFd17FqjermTEZydKaYMA7QPrj1c3/LPOgXJU73DC/9xrcuFluPz0
ySze/B3B6WPlzkgPmPBNGXSbuCbAcPq328bUgl18ue4PgsnR+XYM59p36eKOgVIT
C5ARPGFqAWTM8PH/5GpWjfXYYip0u58nggnM2v7DW79pwkMtBqrxGf47XoWYg80v
JSoMxTtuqFSsK67QI4cVYH1efxCF7t2FNJsmdPLP63/oHOq255YrNdwBxmrqU9Ix
iQmEKhwtRgu9Hp7Nc3hRAO8JWTfyTzHPeVxMQdJtC8awU7AHdtQGyNbY9EZNP9JB
v816D5/vKI5u6OpFcGEUotLoW4I+YV4I9CKoJmVGz065raZM3MahOF5E4AKR/lKs
x8n3+/MEjzyivRnmS8/OWkfMyADaGoylNFqCcnBtX4fj+bZ3Y6HpAc7U4FU7kIfb
wArjH4vOlXYu9HFuINHQFP95hRNnSh82uXCDaq+TgrKun4Se9eTKb1aBnjxzPXLv
TCfbVay6ZnMb4+VnJKyRpPUCvXjBBNLQjlT51YlsZYGi01Ru5aMbs5wT86Wm83yw
VfXMp0MSZw735hgjYi3Ktu+RoKiaqnVuZ9xX4FIN5AtllDEbEJlHqkzQtJHSHEPn
mA8ABBAA2xcMZAdciaOpa1CsuiaGAOr4IJ8csTkA/67bEd5DeVj9BKRWSs4eWC7Z
HMix80BsIwT1noSK9f815lXH/DrYJz4O6e7xVyvcqFceqvLd2q2SqECqhQZKn5Cx
tPoeEDsv0+VqlCyEy/QEbt91asFGDYxdFU0mRzEVqecR9YgjhvwDGnGieFXA4mg/
HvHEK/HToHwIFFzgrz8GEAypHvpiuGPLW+G58E3JKfJ9uF7M0NXMU4nxqVfOkG9h
//pvOMDn6XTdxlx7m5cO6LyEV3t8gXVbLHsH+QGXIETQ79grWw5/mcIiKYo+k56H
05UDFk64toCUfQdbP6gnUdpPrJgd3Y7aj3C8DxlRW0aD69HhEciObmTK4A5Psbmj
DBwPA+aqLrPNWMFc7CuEdVhtSxwYSymFZ1knF1lYeLF3zXN8qTL6GjYOtYQOKHzB
uB5abP4od4vUvErwzHAxQ/WD16FBaKJkvwEgeIFQ1gEH94/zujThzUBT7kvUL5V1
beqbOAoeAIuyO/khgPncje2gQkw5xptp+a2A61+sFfEW8Xob6N/w62VmHzTvoSMF
iymN63A+savvXGDYbfITAyT4UK4naTT605b3vN1rQFbDlzL4PUk2xx5uEhsZ01JR
P0cDL5WtPdV0t6WdzMzEPSx97cOkHvPMD+4snF6pL6+xjWbjAqjZjzALyw9pKX4E
m3kcpj5kfjh0ssJ2kYxOFA4zepeWj7KL2xt+pox6gvAjr8+niBWp8q5LHgc6lLfO
Fu0Hp0mYFGvsdhjfE/kXvCDoiDDG2pc4zxxGGophwyQEREAdnc9fwc+sAHs8snFZ
x4D+TQ7YFV0VGuPAXWJ1F0kh5nmKreijCVDJMW6Eshb8v3pgZg+2yvv6yfbNdhLK
WQfpY3UKlaEbmtjVfw7B04JwTAwWS/cOabN2npFC1xW+TmZDH6Z+5/tPuP9JrfnL
rj+T8GRJ1YCqWdJ6AWRIFlu1qBV9J51t9rgcvtK4ah0+0+GecD5j1f1L5PYin+7x
Phji5OpKn5SG+XftOE8jWOrmS47kjOzA0/WlVKLx/Ig7Rt7GXyd7drGorPbFmF6W
RGy2HDSnjcc7nkKfFXKazEFLFUyBkZ9xZIAo3xWGTCgvanVaS4WgEIoPM7RO5Kof
lrDx83CstERB1dddYJBYCEIe0ioECzkcn76R6gBPLMBkHP1ZWim6u4BPARkAiAbF
YjmSldFeNDo2dxNWhwkfsO/DWMAQ66F9lM7tMdMtu7ualZcwIXYDIE+c+WIMtFQ2
HSiU5/TE+UtziWgaLuzLQylAajOjvZ28DxWNw+k8sEPKkRhqfQClyKJOzK+qhpP5
1Ib8eNXmNYpNcSfGzjF9MVQLddv8QskuB6nULxGkdx3nId86VixjY2TvySIlkkNm
BIt2NZOaP+M5Tb4PkOp/x6+NDn2DWdHVel2H1gViPWSVpju51rpvn2yxk6tY11mI
0576okQldl2VbUcDG7Dt+e+O6AMo0GKtwoENoMiSFJ4H6eU2O9DfzMIIz4ck+QxI
gs+WyAz5dFwLQ6XXoXTA5ysYvO3FoTlxem9wlZA2EUS/YwjsJpXLFRcf2kHx6rCS
e+NDl/iuZBuNKW0v8R0yDM+yhZQtOsr8W8gV9oonV+nnBnRECUk9G21gWCxp8OOp
mOpWLvXGXkwj3rPzR+52jeWIg/NHK5CvvQi7yFEjNOZcDxdtdi7FYH1qJRM0/pTA
PllEnTVPPl2Barg0nDYL6lBrgLvdWkaKGlliRTAmRcyC211YbnUPiKGe+2YOcSBX
StX51C++XAk7H16E/N/nL6aeRrKi5XgFmtyumh8NVHzlVZAM8HTQ7Kls4YDNopbj
2cL03FRIpchv+PrjtXRk+7MSXk0JuL2HE4tdg0VwTT+ulk0RddhH1gGj2S3NBK8/
uRaNAA88REHwMg6F6WAJCNnTImUxToWFAhyGNa2HeN+OYCyfNdRadEMwGq1JY0ls
9z5HtJuF1V7msRliUkNthZrDE+E0x2xb6GF/HrzFErDXYLVb1iKHIhe0B4Ohrl1r
zjA1f/51Jnaci05fMdag5t3/34gIvT+67G3ak3zflV+Bcp2EdgAwQcMIX4D/TbRu
+qZ/NtcwEXUPN121hSRyOIooue7CYukpSNHHNK1YheKeeStOi2FR/q91jnd0vO8a
s+Bfg7cyBl88bEUIElOwGcp13Q/m3Z/FHjmDRXHt2Fxt5OgIToCvHAW2Jz2uk22I
Gaae4Xb46M2eug14IS8qOsBooo3rOUvK2LESfAHjnP5be/ALMMyQY69bxQ5N6A/z
wdfhdabfRspuGKcPCOSj1IkCO3UTgt02l0Y/pFLkHMWzJ8ARUjmdkAdc//q1Mt6R
tgx2adeuiPfBGgcc+xfoqDOSnmzVVSxXDRhfhaGrlxDke4yuXBQCkk6XNggf4XeU
daPfIBrqO3n9ltlZAhYOJ2f8mLCKUBFRfoPIKz/Gw1KQgzLU6A8TAYlGLF/As8qo
a5c/grWk21Kv7tSnk1jlyPqU5gQmjQC/1GlGbRHrEMA1EuXlKdfpRf+xvxNd8T7V
NhNb0CCaP5j6B4lbsHbFXBxzqPxu0Ckyif1+5PzDWwwcflfIVTcO5kPWTpdxSQ5j
DET/VAHCGKJwHw86uBAP6FgnC+/nEecLM6ZUkDvaquaLGWrMW/hIUuyjb0feSQkD
xPRCMG9IHl1xvSzvTH1oLMYpj18F9si+JYQoMJuVz7gNsj+DSRh0aFlbtHVpzcV5
U6VC0K8hVbOEIAxFhpcfnzl8OPMRhpqldZDgVRPbQSmkFE8Kn92T+ce3g84t/R3z
mhCcPUY2sLvoipk811k5rxCPna7hr4Jn9DUNCkKZQ9iDc/ByV0i92HnaK+VsssD4
pRIMr8ahd+wFO2AEqxLey4OAriwI0Ku1OFKVzTZd3W9aJJYMWbYeqRrHDdRHAgyT
4VHUHMxYb/1pO7oGRBEV/Ry0pxtWUv4Q8oWP0YfnCi5mJuB8y2fvEQM0fT8XNepj
tj47TINj4vmqJb/ujK09BFPMUKycVnaUm1DsFpUGZ0CvmnTFdA6v/Ac6+2/uqOBC
RjeS1gOf9Pl49OWmbQKXPx3Boyu4qzjPhc1AXylSPoVTlc/BnCgZfj3eYpZdkG5d
q14SsJMq830BM+huMX32MljJyG/GbkM3BTbsE6jNoGON4X7ZWaFf2oboJbQYawI4
aVeNY0iEBo2qNHZIGmr8Azjxx78rf12+tKbdMpxkGSOp7+k7RCr+XWmJXjkcXXMT
AMo0JgwApFvGpfz4m+ouecAzHQNEoFuOXyk3Nx4lKwg5/SQveWrCfM52qmzhR39V
JWLLFtidMxSWQ6f9zWC4ICike65c0SWxDysASsTb9BfSpkg9IH4fNtMmgpRLhXip
DNvQENCMZlPsB/uk4PTZAAtXnqZ3A35IOEccS5Qyk8jjmCayD+xj7/cur5CkD/Fk
zmm0jxVxnfJJ04dJS9a9zFBZKHfHfTWZp9FiZw/cd88gCWq32imxivNihDbF57Hf
hbxoQDbCBbEPKeRGYSngUTrbXh9Djj5v2+GbWDU1Xehtq4CbvJQjvZShCO28F+gV
T94fbjde4cKuDqAaHqDqURa96/FvobMhwooaoGtESKH6zLsaTAnxwG72GIHPmUVz
MShLsEAz9Ki9/6KJv1clxFM8ehrLnUm6BbGinm1V1+TwJJ05GV1ScHcnq3IEHnWt
Uw5HCtKkB3UwdjqgUI6Mq0dcd3MESlNgeHMmfNsbPnEt+UBfs1N4wJAEVLuAk1t7
eePQdJMh2XgBa5Z1gjdcvpygrDtTo3U7MsZk1wgZakEVQYcTYLHvsdhMaftZrOH/
6RH1e1hPgqE0LOpPDf2nERCQYtlOISm7evc3p9w/v9tWUC6rg6+xqyxaeTArRgPN
3ly3ymsXF48rfpbYbqQRvX53bnw6+6UeUH2jrpgpvYINu2w69dTSf4EVQTl2vlsk
0v1ak/3+ek45c9RtUa9GDwmwdqNzPtKRZuCRYshV4F1sRLvpMxIDCFsKKw/FyGdP
CwtQSYJau4D9KaP5nxrRW8j3xpbnPtEihWp7AyJTYtNTugzCQoGrMGX/29twg0pV
AGznyIVH2n73xxM7Rhdglx3JFz+D1hBB+Z6BwlViwKZK3sOnZ8B94fo9COBHXcmk
2TKZo0HtkyqHKXMGbUHjQnXJOE21K5XyXlrcuhKjr8wlvcng1uLy/KlfqzjIXOdI
egouT8z9p8QTVWQE5SoyoxWCEJaDD9Jx7wbaOpATWkfTNRzSY2pYmvQp9w8HMmHf
hxr75TL+GDzH0NVmio/CBhYQyOA+ozYaGYjqnSw745YzdDNzpXb8TPECo2umDOgc
tDBHaOh+s855c2bRvgP6OKKnnJLcU6ZFwnTSWMbD/6DXiuNfbgz7181Lv2/AM5ts
lACgPkjyfgoXA42CZ0YyNjbIu4ldZLfBHexTzf5ysNDReiUXPHwyqvB78qN1YEMH
OWxxwVylTDlKRHPiprdjTca/m9yvsGjPvTD9IN1sdm/UiCUCtARPlYUJHuQF2qDf
eq27fCkPR9rRzoGaWkkBsVzCyzxyWE52pQ9i8ijSAfamoAsoEfBhfvPBgwHbG3vc
QuAX2oWCRBIwucSHHktqrjW3GNBhF7zp8JUli2bNRMWGXz2sDWIqTV5qYPV1/k9n
yfTCkJIQ8RSW5NKipPWn976YHT2msoGaBzgOtYuLfGh1sWIfp7BcdpyJhdyF/m7H
MLBeDxx31pURPLqfEYiQ7BMem9MNFLf5DByh03nP9wqO4QVX57vtkssdYHKN7xxE
vFngOVRRe6X+jHY0a3e91HwbVYUy/e5ZrUXDEM5pG/z/QE0Cezc2ERhppQJbPe2y
fB22XuypedFmu0W4E/QkOiAiX5W2hLlZyeyKeX9Tw9lg+wOaaMPPS9JmezW9WVZ2
PdNsznv8BgXuWIip4wwT27nFfgXtAHMlM9cXlKnBMEdYQ/9zHa1JnGMao1bQCX+K
PUVWGn2/iE0bpcgpzw5c3NyeMcQf3Daps+4Dy75RGhsGdHV8s4eu4NLLGikMYII+
8EzgfA5lE2gnsKDKcWCOMKj8SLLY7oVQTi5KVbj6hKqGuDZL7FTUtIKZXCGuCzr6
Ggpr7+VWrUVmqarXFgTNW+xf2Sc5t+aCpVJG95cjqtDnMYzCqkchOuEbbyaXwIKZ
emH3wO5g8A+qjzHclVx1Z6CrEDX/nr6aMfwWIosyKZ5PHSqPPqOsbCeTldQfNt/h
oGTwTXvJ9+owXEFvy35AgF4+Bei5AuiLdpLLd36BJrHi1Sc33bB+quPecJjojwFu
aTWTCHmAUEtSTJxPgBggrSSwKfQw7vmBrLyajV/yZr+kVX3AaAIPLFtV2umG73/k
C9xFuVv9nGBGIy1Kfe1pT1QCIk700gaLtSGnjCH9pKFEqb++s9fOn67BhtMpdKLi
t+DFx6Bf21mclFjqwMvT+re96o7JED7BrWgTtWgLFbtvUzGWWUpvYwFlHKrO+TOZ
Li4m4LHAsw5VQneuZtGTxVYHJwgn/4dsY1mYW+XeBF3Jzun+0oXNgpmdzOUD1tuH
04dXRWEvDhq+qFs8+DErFkR+rO3hwERjZVH0T2Y9H5gElE6EB8YYNhbnpevS9pEN
7Awx+PGv/xcRJUJSHyU39qstO67HuXEq0zHS4eJXwy3r+15ipbtGA/c8b8jg8io/
42B7MOjdkbAnPCbYG+cJe+rFjK1s2TXUzHmUkvLufsdz0I8DPztBF+INEgYA5Ig3
RA47jX4iejK87q2jf1elBhtB7VnWUp//8mSD9AfOokWxL84j5QwvhWqHGGDmePwk
kxyQJ8vfVKhTw8ZH/0IvTIbM4Cijj95t4PVs1AwxeD0jwn16a6NzHazBDBo6Rn+r
rwQ/SkKiGrITkiBAdSf2w8/mXIeepXhbEGzJEDxGqqZo0jfoHYFRTMY2XkvjBnrm
kf86NBpYYOkN6nf19mYnEnHYpVxImXuEZSU6T9F8osQ6lkBx+3O4Rm0cfzXIc3sG
Q42xegFiKrcaySi9u+Yp4DrN6vOqP7FB7i3Kkbht9BPLzt6byS75ovYK18KXtR+G
jh/EGgS85EbvwZC7lx4RJoM3AK9DU+lYar+igq4ZeYbDD4/dxKQvmx3vEmUok3gM
P3fleYXCcNEjSHPM6nuxzolvxG0i+77ziDyB/CTq/L5Jr/o0/BqIWFlXzCIFugM8
lsdwoxQMlpXZdxWeI1YFOAq+KEkUlL+NoEuklnt/mVBFGxa4ey0iQu8mW0Vdij6x
BoPgzV7IVOh2ueh8XHTjpWfchDKWeOqj6fCIA6TyBfMRmri+rQ8Qb4YUthA+qzGr
I00r6DQIF7IeVO/klXNOlNwX+1kWgUb/oLHv1jl4caKokkzTMECG5BGyiLjxVybc
sqSjUw8AZtVmFAM//ZuqD8eIGPgZY+61/Y05g7kAcuYTsNMrMAY5bSxZJkmJMGAc
5ZXX1kpvjh5LaAyHyyZ9bcqkBhc4v6GZJfMtqU93YLf67F7Ej3jVeDisZQxI3nop
bd9o+Ks8Wf6QYRLeJaFPS/zDO/i5qcLz7e7iBL+kCV6TAocxmoiNFCEWlDdsAqVB
bkNZz8RPgXH4Tn4ZREg4YPbyUznYeKzoedwFaFDl8KO68i3szB5XJCFvkZFqjzW6
YE2s0hb8hSOjTPz6hzau5hRGIrZ8bBJQcMgZyfk2SyiECLjC5KkT8KPIDHpkPeKz
JKs5rWDg3+EOPjOK561kzXEDMMSQR75J5H/Opbk+xexGiK8MOfoX7kM1a87k63Th
I55sGbfhUE3LRCJFjfKeGfrigY54bzNWK8lc4tJU7jZdvOpVDGTFOT1wAX7OjUVP
Jm9p0CrRtjlxwedQR37gRFh5D+SNtwzRKJim39t8nWnH2MkyFtQyFx1pal3429Aw
SU7yyadLjzhSShCZiksZKa8NfZEbBQV9oPCs33yYUO/XkiOz6b/iqyQefj7DCLoH
ZfuaGkJxAWvJ1J18985m7W3qsk5l3Ec1MIZmtHWzmikJp8cK70bkNckDlc7K8MLD
BKAnFqX/b285T+XSW6Pl2BSiVgWqwAwpn6G1gfOiIZ9+isjLM2aoLveA2o7NmJTv
h8E6ZP0izf82XEuZ4CbOI73ZnOEulvl9DQYFSCmCQ9laM9/fr3VDyDcmk5DGxonM
AonrFcc3g2mnONhlV7Hwazu+bpqcsgacga1/RQZimIixS7E1FE/Gz0v2XwzMpgn5
0lTcKsTxCfsgybMYNUjZxXoJo5vDRCz//luHIXR+q6t9tHShe9bJLCmqV//HfaRw
rQ+RtuYgWgSisJr/vK5ZehBVkiKmJQzYI3uXsOCZGQBhhFpWiYGZBAKP5l3bJ/rK
JnGEKYcDXrsHVvvprf1myNwaf84oQ/eyz5bfYx0IuydvEc5c0UzSFoj4tS7vWqty
CIIBCaEYckUI4WI3M+TaVXSHAl6vZ57e6bMyGeFzkf3DrWr7KsWrWc8esdXp4Fzj
QvIngj4DtCljqtMMjV+wjjOP7o+r1tfY5cFp50si0C7MgNI5a/lMTQWGY+uWNEIG
EHhEqw5UX3Ttmfr5e+7fiPDX1FLl8OkAw+F23mFDfI2XjQX1yRWZoJR1oSHpErEb
vvqqfmXXwKhYOVOsvCKiAvkTaaJ4+nt/lOf6m3XBKtCkOV8gYPxw9XbMFunsTv0w
mApu3siqA47UcaCukInfNOHoPcUGjxintnC/5y4iKOBohmZSETqDa2FpynniWW/i
72WrneNuIREEnQaw6EDRMGwxvonw9AfTsIZa0REy1LqK7J0nVvOl9TZCM887+8EL
GheUqCV7hCKSBcPyTzspO9SY+65b49jzfHFX/NG9jkxKyGyyUAwSQi1ei0H24s5e
ukBjZYNViIBKQzGpTcEv8OKSPDiesllCpJRlbxFtn9Gr94ugGow8zDIeVH/DzUko
RMc5XjFZp1mUilhT5NrKM5c1TNn56Er3vHOhx2gZQSfOLvfMuDvbIYmphU1W81Z6
0UfefIHTkqyTFioLa0kZrQmYXFSiB4TsczEEUuvGSxOyi3JihHvoSqwVJGPooAB0
1LoBVcKQ4rH+9t464i+aWx82emMg2cywe8XXzYoxjkG76Apx0feUrFk6Uii25LMa
dBHbyUChEy1mQvvkyyhkxavWxXxmoWCAr+6mJBwHcse/K/FV0LLHp2ZyL2dJZnJA
xIbC69g+piDNyIH7uTum+mx0w0PVDEJvl0dhdo5vaJaDZHkO9j19YDMx+8aR+hzk
BLaAF/cMnHKLcN4BcRtfIZrjSOGUlBWChFy5BLhsUT5g4mZoD0nvKCX0V+IqdheB
32eI73XRHF2J26Plidrb0FE+dUtrlUfVjoXSI928lJfEoyzWdHqiuKr+HfwhP1qf
9ejchE3rvMvU8mFQ6TI8NodWb2uD1B+p9/KCpashaWlwAvt9CkxU1DvtkJWl3GHy
tNgETOs8UvWUOBqR0+KUtYMXww7rgWcJoNTpWV9o2+WMlzlGWQsrlYxmyr6Idp+I
++TZNgYM2N75S85eadA7+v4OTUlWSia/nBEOpH0ZVT0gQA56xKmQH2kcTY5bVVbp
NwGLGP9KHRkKGLEAfd4x0A/YYc+l3o05w6shN9OlCryk2wUWNDTDZHb6M0p2+PJp
Q6Jek4GXyivLYHUsAf0NY10FtMKxMk3KkIKrcA803VEZMUeSQRP2oc7JPDQxBUOh
Z8FjWOaj6RaKiLPe70dzHcTNMnFNkIr0LKANbWEfsHK4hnjsjBUHZ7cGVUyMBGWJ
6bV23CH/3LWLLGcmmNs8obLCcMbEFz4HD2RDz+7kdnpRf3kykoobf4xnASDp0bPr
9CDZHOkcYPN+8f82Ik4rgOxx3CyDV70bV9WqcYUrLd9I3EofeM3mLg1XBX+LkgMp
p3jSp3ETP89Hjn/Ss6AdC2cfOnAwO5IX+ULHhPh8luaBNS7zpZGxM9mIPt+tJ5xq
PgNsVMgWqwuw7ZxqQZAndKcaAqmdkWHPpcstDKWhMELOR8wa+v6iPegGChFxyyOp
WBm34L5jqIj6Q35QsCk3gpdicyNjM1/Iw+aOxGfVDZjaj8QBUxw1Pj7aiuLrozlo
UYqUoL5L/prtO6W48ayk7cDCQai75Nh6oDpRfXjiygjXY9ZXQlIO81HsGDoUr8cB
5838K9XwKBiohIBLq9rh18FmyPpMrf8+LEVmjNXjUAkqqNzUowAoi58/XCkJcHDP
Zbd5CbMwWe5pYSLrGeIa1xx7yrd+Mz0s7P60M/7YFPwnmaF/6ggurfosMYY0fMA6
PhmmVgfK979iINKJKJnJ6GEW3kJ0Gke5UGszt2lZ1y7+eZ09zlaDMHs1kP5XDSQ6
l36inG03lo59TtZgnpnJ0lW6XAVOYbz9wftjYTYjl65s1Y+lo6e+cvqQOHi1XLiR
jg8kkl9ow8oPbTgy2F8BN3UMVF+Iz2j3nmSURRkf9MORr4XL2xYVq36LEVM8h0jh
jN04XCL28i6bOFYLUlSOlVdv/L2mcLCkxZ6EUzGJPEkSJdA2Bi5Ag7KFiw46cRZB
ifetbCB5rsuC2/YVR/W/vRiwMY1urC3grzMoGMPTp1zgY7HguqEuc7GonR6NqLuU
x3tcYUZ8diA93T7hfxdse/zwW+sYIAud3OW2J6cc5E7os6+VF6M7VJB9aoDs2707
2kOZOYQgHARzOsTWCmhvrrUst8C3WgdhvY4kGGKvozhOZI3C6RpvqPZgX4viwmZY
PYkk251LijwoLyzlxEXOZYEMIeqD0BEWFSo9sgMRUB2n8Wh9p5x9jepQFZftqE9i
l52xcxMQV949B0mv/5ZdQW6+dd1Y2VK83M492bWSan4xpUvhQOL8EF6mPGXChGGB
lhcq48fwxkfUAwqKwBGOmCMrKQUnipNeQkigCVP14Xn69axxRPImro4tiSBxhmyo
jyh/Jii656SWW62s14BwHgM1PfQd67UjnONwQWzBILaXOA5mPV1mLEYmkiAJ8b/R
yh8/oBScXq8A1qiaWQJMdq2gUo0HLS0RSyygd7WOQkIICzE0LuWIUUhqzoN9t5l+
D89zRFG2qh7MDGRV3EScm+jnL4T874Jnihs/AxhisgTpvY2yCxrEy8Hu7813usy3
ieKbTnHvS/qHgv+AqU00Hg+7nVbw2c0KPBkSahvRV2W3VcBZReqLA2GTHqdZUUz6
CZd9ttY1eEZsLtQ3RAzOw3RIm20cKhETk+ZgJMHaRs30A1KQjlQ9GQT5A9Z+0qT9
NEjWWh7LADnHnPyscquCjDYC2NQK3NY8cFKOuIMUMgSp9xDHGD/q7jLDyeuXsmAj
MYQcIAisxvtf8cfC5lkQSNEpQx4T3TjsI5NROp4xJbAJ98WWUYmTDpPmB2RglCpe
f/AamNETKa2ThKDIFBY4RwPqMEwnFc7plzURkd7JopYtx4gJD2umJ07RHNRwglK6
x1xf5m+45D1hmd3VXEIgYLO5FDSLkWVnkI51UPuf7cc3w9CuJ/KXShT+000IwQJ7
TsDkP7rgjZV6aUDKzAPqQJDMaymKMQyr9aL5qsR1+k4/MQUhir4d08B9bt2CIFgc
WRACjunMR7MYinFPuDL/uEl2AjTD0J1U9qJjr7jUP32ESTvoQqxd2vSPQaxJHPFf
unIJT0rXzzVRnhhYJITr4V3eDnRQH571J0HrIzhG+uw9vhAIHZxtZYrb01IR3zqc
C7FGHBBIUo/RaxeopcA1L6gJ4ewGGC77FRhtx0VEH2+YtIP75bbiH/NZmT2252y5
1MfDHdgeiAtkzgIDNxAdHatvpPHGp+034Qs2Mzqx/1f72Znn8nYxQsA+LWxhthwT
HZh9zYUm6qp4Lpj5uqG1oxcsX952UPqf5zGICW2yt3NJ1uYt3YCuQy/C4QKs99RZ
Ht3/i57t9amkSKUeOrVsFo0GlaEkMFShC7PO7YBOorqK8hBPiUY8+vGKNxzX8dB7
+DpQfJKPpDMRAxS1A0GSBNXCSPWpYNRzzXh+QY+LKw/AUNWp2RyStpUOmLk1Jn/Z
pRyAhKaZhXLGJCHpVFyaWI5pb5o4IuecpihDoP/PgXcz1Kkermyj4h9gQsSnbUHK
ELXNKcRAbnDktAftuZbW46lTMMoVlwnAASwFXqkL3aIAChfy+HVAKfZ40wTeWbHe
iD9Q1K+DPNqKcxjEMjLGcLbvyi0e84j7lvi3zvalJLM3OwCmn51Nv4dRsVU60Twh
DM11D8zbhEJ4pDHZw3BupzzH8FRpwOHBkZGRqQK6mQ77EQlQkzOXibtZFPfykk3/
hORbaGaFJUC+5OKb+ak6GU/tOoYyZpU3GpWZN8UNTEjNP/u3afApcJp1XKSClble
otyFE1qgb2OzhyTpCCzLiwq0XUBYiL6g8CvDv6MMvcxPIon5Bza2WjjLFz2a9izi
Br3CnS9MsV5ji2X2e/jenuRMqmvCyPHjtvhx2PahC+zKmvCloG4Q9OX64LUmaKA/
HzLrq5ztwFIiIX9J2Rhaglk/mc0xMg/VxQYEUzin51ljKsfuaPesbUdwyE/6jSUe
J8Qrlje261qLxHLWklBtrqRaGbnK2S/SgY6DTTis7j8kmxyoNouPh/0lKM50ZEhS
MWGdqW51G5rHhZNukvn/rKESilfbv7Avi/et7zlGSHDPfQcQqRWH9Dd+5KvUD5hk
mIu6IPe5y8VMWUMa5GyVTYZotUSh2HaVUuN7sjF0/hXQgFyQE0f3DQGxnV9EF9ot
gn0OpqQM10S9ur+M9q5N1a/uTdFbr0j8qQqvwjCZ5Y/Ajfjw8LbK6qnC57KSnGnm
KicHvpAXsCLYSZzC8IfrljSx8YBl0vShH60azXMHi1HgsMj+Yzi5lxjAzQv0Ndqa
PZHBWHpzhzjIU89Y4Nt6qfDHm+7hKDLU/oP1Eyhk5/75btymZwj+22KNV/29Q0u8
dThYdQq8TxF/DeSgQrzZkQEvdap6b98smQt/PY/bcx/nECWoA5FWKfFhqkjBnaM4
yClFZeoJmRey5PiXiWXzfM27yY9dV8vHx9mGwJqHPWUOT4aKUIW66/Gr7CZf0Ikj
67HaXROnExlQuwuSp/oEQ681ualTSswBpfkDbr6l7IdMfRERntqQpJVAa4vSCP5t
qlcM7Fu7dQgmD8vTjVkzaMfyV9heHPIbV8G/B+p/XuBV4LOJGBJG4oMHyK9NpiDD
QP9smBlAM2/oXHsF22kBmZ9dlaWxSbPKLyDHZ7ruF16JFuMbhaPL2h4WQEQtx6XS
mIzPH9EDt4fBJkI7WPbQJ1bkMsjgIbLzLxEIofXmFrksXXrKt999/0yNG7qDHooo
GYk9WTOAjIEqBxaOq4NQQujKnqeZnQ7WKWsXC5mnkOmGHokRO8TefwsTRoAaG5g5
iO8fpH3PP38jbBHEqRCF6GG/jBz3IctUCCUFjmQ8fTTulHKs58QzptLg9PQTeltF
Xp/BVXBYlYCFAfAM2FMv9CQdNRV351wbrORGcMAl8e7EUBJjenih7FqcZ2hrt/B5
5zRdospkj+mSRsgHcUMdbCrjYRoATl5z+zEZmWrtG5JzLeVLuqeQmlmJgJmXG2I3
NtZ45+SObtZY6Lyc/LB+9VVXSymCjD5UqYyQOLDkqMnbPQZT6RcjxCPnBaTfgtx1
YSxxtPZX4qCx+0feERKR4rmAyyt8W+WiqaQalmkwnbvO+8xelnMrLgbx7LQtqlaS
FWgEeGWqYBw0aW10h/B5XoreDsKinwqXY2UUSY2wRXQorUqqTdMf2jkrgJcQzOyy
AC6XFR0e171rretk/jD5qpKB22kfoptSoCqUFoVvlhyh/o39ezqLLLmSpVsxgnsi
x1G+6UmRS1f6Qh1SVeoEpjyNmlpqvfvHfnUGiZ9jHo0slOisYBEoolDpM0pvWXY9
JRJNaIKZzMrbPDfiBUQJR4bWAOEd/s4ZmFKOoeaIffmhvSMQTwECqJZc23Ylx9qj
Bo9ic+1spmjrkXtXPMo76uTnMAlN7V6hmVtk4iz0cJbr4NbAXKRdyswAXhCH60Dv
K5JFDJXoPUkem9tJwPqYXZpwfIGnL6dRaHHWbsjdfYy71hRo0sPVyC0IvmfvsZg2
p8xQ5nvj9cs6eBtDGij23vqkD/zTn4qaaiDA2iBgkaeqb8r//ThEs7MZbNktQmOm
8ewvqfodzoi2uoyxSWdTifQxlS5ZZOCRNwDEvniYMW95IhdeTBlm3hBShVdmZ8dP
pJ2BpppM52yZu6C5Hs0OisIEMey1luzV1Tm5QgidRveACghGsXgJ4C/ipoOMDcNw
kjRordK2slUOyKX6kfXaqS2M0zZC8M/EEIfip8IPPkN/faSPX015Z79N6XhzVwct
h9F1Rv4G2HRDfwbMs/m1Hpb6weO1uTNQcNMG6QfgI+r+9jn2jR8BpHV1hulSKhBb
8xNzJJfDkbVVZZhBnkpWYR02PxtMDGpNMAsbi0wL0K23/57ciBH01JRcXew88o1e
I0GupJHsReqyNbENdbOOvjooU+UKJRPWl+KHAb/YmtM28pwAGJJDP+/XqzJqNudP
l1mkuV4jpJea66tnnf6zPvRpfiuP71/xmN8szlFKCF1H5MMHemP+1GE99b4XO1QZ
Bw3DjwcLlZQrAy9VaYmWQUi/+WGdLqx5qDRIPnndHvgD8RbZTPEMQ/g9hWxWjc96
pNjZumdEXbojyhbPalBEaU/Wa9t5l837G1igrUenaTgXXjeGvb2yEq3Y3JNJPoz7
l//XpmjrTjsxuECtKTj8xWz/EL9SsPAmdEGoi+vLMuHX+O+1sOmaxkPDRxYXepOd
ZNi7ZnMC2vrrMK+q1lQzY93IdxD2vxgV73B6V3hUiWqcwYTB1ZADn60n9yf3QyRD
PKKaqb3YAtrA3Ysoc++aPfPWuxq3CMhrXTrTDovfDUb4eKqHxRSi342QkWB1ZQfi
0cweaHp9FmBScryfzMOsNURpAMO/A/GP9030rWoudiH2o6VVjm64wjFNEZcpf95n
5f+wsvcPKwv7m1pmCYv7Wfg3CGcCV+ZpQW1PcfjfXuodODiECDX6o35Tp+K1yOSK
3ofMURO60qb0JifPnfF0tnV2Q+SVvxFsmaRwd3Jq+f48oyoFyVPgduJpKGzVqKgF
lKK0Nm2G75eGUBt6zaun69uGKqb8d09NJr4j/A3/ZYE35Ks0asbOjfa9x96cCYPt
heoRiswmcvYeSPPwdV3LahyiuEUXm1ox3PwlvY81QFGlN68TcThP+i2Q5oNIAong
GKYoJquJ5OMFWbAo39C+TzNIIG4TUt634cvZdWgq5IBrqhA1UNOWO0X2OOUPqbzR
0JOroYCp+ma2QlpA0X9GM/UvOX6Ngqi5+RN034Sc2C/WfGbkqyQM0XGtobsUA0lw
7t3tlch2+wJaR9br+MjGUuYwDGCaKF1/BZXRQ0Fy3CO1iVGPBxFtt0jIhqzmpKa5
/TXbNr+CDROXWQayltvFLzqR7QYQFiZ0yZGZeN4LBIYYtXQZvO23ShWMXP7ncgdM
ytOzDBWVhWTsbZjFuQGpDs6WHOdPMb76KiblbvyApxnZ1ZqGYp4YcLBQnXJFLGnh
5xOa3vXtC1y71xZTkx9DxNp1IrtG2qmd7P99whDDoW4Y7cIwQg/25Z56hLtGqli7
65cf47rxR3zLazhx3XszRVUVlUhThqiUxFWqBvPMtUJWZzMpbbfMtAL9vBCuRLYR
YqlJ00N7OUsTMlF6XNqxitPHOX/hCJGKkOcKfJxdEZKggqt9DcV5jTcsT8I+UARi
GkjakoemiswyBKTPqnP4jE/6O2s1wUhJYBTKOqJ31aEB16Dngunalwq6BQ2t4LPs
c5fZT850dLBZm+OLs1ak3o/lEuLx8d1rcBYlTC8f9w8vaY9dh0+H/SCNinDqTLLW
/0P5ZUR30kx0dRrU5FCuFN4q2LVrWekBfWM7iq0aYjyJ1Dxxc/uzFrxk5EPCuZa7
GO26d8TTyipU4Rb0CRb2CbXEOBJ76COHZh3A5R9CduUmtbZXsUV/KMC9o12pV0Il
Rhr8nSib7BpGBTjOMvMsiMbOvZnTbnzLsheZlymwjaLLUxUYmOdfHwX/1Eo5qQAs
7GAyrBRLEeIato+yPHB88eXVBhaHoeAY6nxt2HFqS+xgYIIadtDKkh5FwnX6hXNn
YMSj0sRv5z2yV0dsvfvEQPoRVBMbjrprk+d6ECHydSxaPzYiFtitJunVKzqvX2BJ
DlWZP3pPiBa+sSoCh2u3Z9qYLN3x0amlGUp74glSTVLf2SD1i3/sMHBH8uPQCxIy
R3kpbNdfLzKu+92wrGH5cBbQHoBSuCdtxOABTTtS0wXg8vbw73VC3KgtCt2sSGc+
1XmXgtCoBYyx6RA0yVMbMXAiAxkjjZi5s73aBLFlfgCR9BPDY1lzoTduRJiO9B/y
pEyRxPXQ94M1DUs3WWx9THYNtB5RmlEpjm3zq53KkWYXUuoqRDwCOq8+6N/rDy8k
U9L/nCtHYlULTBlE/t62d/tUnMQPVjpu09+WQCG8qhGa7an1ko2MPlKJYmdVICeu
EmQFSN5eDXWAcl2myZIov0c+z3Pl074uwW1SwVSsdOCIYIm+HFSqtCYupGCIHqJM
Kh4diGpwX7zY78mPRSDt/EP4ImSXYNbGzwlSHcYwmPeMqIUFLfsUoJ669TJMBsYJ
+GwdI62QpSCtBUHIl8ujeskkzXeGSEGlKgTM9KKkoBwmP/OWucqiOMLMSjt12ZRG
1p+1mW576VhBgiBu415TBZG1+XOkHN6IIGqGP2gicGnm3+7csdVmGEVQfDAHbGAF
BYiiTOmeSDsQ/BQTQ7PHc35txv2PKJ7wFMCNHSliaQEd2hdUTcAyuMTQzupqGB9b
R7Ia0CLh3M91R3pBxlw6S4rSSYJmDUAAInKFb+ufEovY4U3bLVkVsbqvOGwelLKF
Rcwps295dSMB+tXnJSVlUvjg1+7Jd6P2BO4MgG2pv7KwkGPO4C+2WuT/suHkeMlY
HL+3Mgf2vkuy6PsjFHJOMZfxzq6XMWPOU/LmfU1dl/urYAQNzj6UGuIRV35ajnKA
blJoFxBpbyJLWQxj3GHGZsdSOjqQYW2Is/Y5u7U4A6xPnbkFHSTSKvBBWVJxX2VC
wviIjH+nuwGrk9pfoR4elqQoUpgHMsi1D358X5RdQiZSMDxJWy8ZecRa3hqen+J8
ZcY46YTh1OANvEDrB/5Y3htvlxKOJkeoVe4DDEw0K1yMJiXt+cthhcVTGdNHnPTf
69P+Q52gpayZxhJktzMDCZ27npQovWOu/2hbsOS/nUv70HuVediz7IWaWHy7lqeU
AmAgbtTG27rD1qKGUEicNP25wwInGue/C5WfVHGE4VPe/YtV/oze0RBoPzrVWMIc
e1HNlpEWbv8KF4jlt/13a8nu00UbKA1RE8gwZrak92wkVth3I4bq+prNZ+T2AVIR
sGs/dev5Ur6d2ayngn3gJOfS6dGriKCGtl1Q/Kv7k8vPyYWFYhZ5gfN+1VBWQRSV
alKvyEtumYVtDBNUsmkj8qY8CfVY6JO0pCruZK2p8CdippKoEhD4jR1PfEoVkMi2
SV9/AZnjHvA1Il5B7+Qfi5qnhQwG+jPVKKM8LjafPRWvgIWCi5sK1THqIZT+S04H
lzUeWlewX0eZrxwfE/USerluYr774fqtorFNlBlycX8zg2rAyDgdtzf7Q5xyT4Se
BZgloUCuCf8KZklbGTHsmgAz1hPoIFlQmlpZBrNpUj3tl5sDKM/JiIcyll+rhnkh
HNNxz35qqmJomuK99/U94Hlj10YUxHv+q9EpX56ogcPI2A4faA0E5/wWmhFkYo3D
pAMYGrIQLM5VZhLqUCRM2C4RpNzwPjowngXZ2J3YvR0Iri1xNzYKZdQLxwslEy3H
ZyJhzv+DTmFMmn41y32K9+Z1gMKY1eFO+98a0bGoG+r14SdNg7rGmkNjNVBB4JVT
6VCu8DpR2bpBJZrOjzn4tujWc+CySidUlnNlYiFEnoZmtHPA16/dQn4dwwkxO9ce
fF8pOS2UiBd/pX8j7DJ29XqSsQ1hLSUaa6xrkpNww+quC2UYYEuZiBBCSW66CVwX
O/Rut8DEDAtmdojpWzVy89stu/mR3puXXxqlK2ZtcOPzwqu7gxBBYOWkQYV9iUpb
sp5WaTMmCrbAM28ewMQ9NiLFt3sPukBx7HdWajP2vmhGH724lwswfn+B7XSI71qH
qaCUx237+58244m4JY7gsJ84TU5rYB7PSDE4ZJRYxHoJSMsSIalVLa0y3mBVQANu
AJWsZ+2QKVb7VV7/tdd6v7xtlwodmYCASUljSz3o/nXlw6vjIXPHeJqGsyI9Zw/C
9YoEZf519aQDmtdrbP4+CXJ6JFo/SqsD8e4resC3JxWpaF6Bf8mrs6D9+EqTA8mB
Gh5E2nq8zPXKsOhNKjTQ6WQCqJSVv3YbT8D265gfu/t/TqFRLpPiws5a07xho5M3
gYxNippxshUIfudkvV+Kg/XHPz7FulhFbLWxPCecfMbCXglVu/+6+7QuHZjxtE1S
aZyfiNGxQcapXQfCPH5VBCywSvYfBHfaIwuzhIpWCJz394MBMzzRtqwY7EnX/vT6
OgBy/o+24uop09EkHTr6rJ85eLe25rTIiYSnOBgPAT05sN275jIVG/+PVgu1exh3
4EfGtyycHqat7ysntM3zjOs5mRfu9iV22QYw93iBO6PAk7MgmZplzgXUtBBsgeWZ
DA/7rgnOzSdMzLa4J0RuYLp7lgRdxBXeMNaQ2WorDl3pBzeDlJpBFq3FLpYDsYH7
47LrKTB/IyCyiz4yoUcuOykKHckIBjqgn5QwXSUobz6UWJ056HwuwEsBeFNQZa2Z
6UD5ZLK1HAwieNs9OcKr/SZASTRrKm1kSDDwF853lSrmeoFwUEQ6rTmsdouSJOqc
oQpN8vgqdIpYdWGllDSg5250YNigrt4VC7inNHiK2LFo/YyTqxNhLkvuFD1dv3MB
K+QgWtvJtuMsAdLLi3gcqlKP1PhkIYurx1lF3XZrohGXyku+s7UEh0i0bCV5F2XQ
sWWyNQVq3hbMTLeTeRbBgkuRRhAT7vN+KltVqXcYzlr7H0ybuuG2rG2Bo3aIT0a7
V9ozvkPDk9rOIWuiminpMob4AKbQacc4XOXCTuimgSxOSwQLN4D/R/5XAoKfOtIo
d2/EjmVkPh1j4tQhMRJ+lYkRe99Wet3RWWS2ag55HOUON/BcCXVXXG18Cdibqrrg
O4QRrUrStlj/nYoBg/rS7yjhLiEbk43804jcPt7ideyWXIPqQ5B7l+gSZoMeteK9
yKdMRZCV4oe0OHqJI0CoXdNoLGPTcEJzKANzjia1ORJfQHnNGb2Fdn7+sBXsn4hM
9w903dc+9wqw/JOyM5JfaIaclKvVSIoDtUibI8uQdt2Q8TjlU6sQ+BcPQUyt5O/t
YnldeopqbG+mdNN3vgFNMUOexDpN3MPzpNRpjNBbDNGpclW8pXwShKOWLO9lviU1
ydlvGWrR1lLH44qjJ8YK9MjwhmaiDPW2ENjBP479//+LmY7RWvH4BxRTHWjYLsJS
+F6AAZpROsUgzXanDKLwC3sblGoCo6ubYPFVR1GFJqP+eC+xlNWMuhdHvFJn9ySi
RGMlf74p0eqsKLyxz7C3XYrRHGy4IuZ9wOX+Q6OGSd7jiimRMdz32ddHypvgLqav
UFbmmgXK/HX3gDKiUjLCQzMiQi9kMt/MG2Rd/BoeFF/clpagID9kpMj2NJM156Kd
IaV2LfDZbLjnE/RFVGz0F99luG5kUMXtGpovMlhqoAaGcQEgoxuidsaMZ3aiwqUL
ST+NIs67JuSLa2h63pj/CF1AdgB3kRVwEEheZwdMoK/pVfjVshK6EHfsqvc0yhsd
L031NNo1W45FtyCu2U7wm8z5wlzDqHA/YxixA3fqt2VhD0ydnah87TCAGVKGWJA1
9syCPzmZrJTBgz2GzGo5d4PkcsQkKN+viK9RMhn6Lnt1JUVd+i/gKx57vxSA7nP8
UAGlCTxD9mZXVc3joq+x5RngGcF7UQFWBogfWHSXIa0g59hyCkxSqeiwRb/Whd+d
EuzDNWqwNn+qrnxCdpZzoq+/S2KjdyYcGWrj0jRVRimd8Vjp1m5JweqWsnJsa2iV
wJYT/8aPDV9SDosMfGTzfx3zWsPNfrmfXpFFKXV6bolvVJqHM4oli223yEAtNwOb
xmrwHalHOUAAz9t28ci6Y1l3kKriYzvRMxCzSVLX1pCx9tAy8QKIdPG4108pYdUS
7y5xd34zwAU4T12G/AwQLV1TwXp89+5opfgow4l/XEbAvUM3Bamolo7TAqUHIPNn
DZyLhNOniXLWFpsGrCNMnPQH4632VRqCKbVqTMCXZn8MBaxtxFHcPyerpBofwIbR
7YY5G5R0DglZ3tHeawF+LQF6rWmZlvD2jPdlLpOjw67RwUBM7iFNagAEi6OxO7mk
q93+LdAo15jKBhMEBsrnvDbBsN/w4Rjv85Ct32Qfic52OGo3JkFszuVT/Vt1ZuF/
FFCg5HQs0u0ilgK8J+BiWxbxdXGa4U0QhUeiq7EGk9ZYKl4OOLyXSb8e1O67/TYu
AVJWfH0+MP4TwbNC5bst3epmG7UBBX51SRDIuaZQ36E0vWTyrQzIViwXbMUcg64V
OwN4WTVK7UCE+A1TansXHxTwPHTeTOJodTXfG+Q04vs8pbNz35uDWKcL2a8mVR/9
J7k2Mz1vQEcvtLrveLf1kWyonU8uQhCOb0aSTxNuVVUEig2lPAixU600d9xNUQgD
6WB4CaeLTUv4P5Dy8NRq8OxM1f3yDhMTXzzYz/Hrq2Pa5uqqzty8Z8q8y1TsFe25
1i0eOz/blkNQyQpxJlcLLrWEi+RVGAo/DysY4jegXuzAEvq/XoaTK9wYILokduBv
O8OQn/Q+Xyn/IjlvBERINoXTjM+su8hvZIqzyNQExeC46J0knOgkWwk7OZDvuP7d
PCh838bbgfA2aLwSrYZbMaPQnlaLLHyl9fGd8w3/cuVn/VJlnyJLMHmRtX0n/xsE
VC4PC8+c/VUNPhqmu+SYsuShYLRg6IC7GFf2yBT1rPx+IfbUPoXw/lo2tRXme9S/
TqQakOjxh5fYZ9R4hrBPvghTlF2BQWJQFOzLXrqrmkB1ibfUXRpvRxqp9A7/1K7W
whI/prh3ufR60AO9FWeHqzneKZ7Ko1VOSUhL1VBSNrhgKfZyKrb/xlWUC8NCpS/x
1L3RQij4fHIYSPRypdW4kjgDl2/IZhAsa01EI3ygI+EhwE2OjpeS9xXXzl5SXqz8
+jYrJPb66xIE/ZWtLppsAYTJgdz0YJBI98wMsPrLOsZwjeEd0hS5LclhE6rS07iW
d9pApyhe5YxgEISAbEz2CWHEjvjcdOi+61mzGhKSMfkozz19FmoTEZIxwmvNXTwJ
gz+7hwdJztn7fdUdQNwTyquE9vcE4dUHlmDlIbadiarQnO90r+ZeYQYKU27UU3pA
iVd4/WzaYVJnXHa8DTi9lEpmmcufwSwzrDx89HxZArCW2z/cT43l3y7vymncUmR1
Qj7H+oNyhLBP1ZCsNKwt9nSw4aRAh2dtK5tS/0agr9uRkTVffCSDaHR3pchopQ1+
Q9BxJCroME7K49TE5hO5WUby+81oRO5cRiHHNcOX4sOtG1VcrdKnDK2LlpbzScjw
KXOsZY9wtbKhdPuITrGpsQUfhZzmKQVG6J1HXdnokkylnatNnkW9xPf+LqpzOzs5
7GV0+nxUJDs8JgQ74aImxXcxPA9lWi7pwPp0ERR1brrfs7X0qhGBDYh5JvnNNfIj
ArylGWdroS6EoO4FifYdGKgTupTZLsqbvLir2LSwbAVaNrWRODwHW0sGS4iYErEF
13DXFWqF7O8H+WTYfu2IAuwtsFesCEakkb8vBynMHyuxkxP07UEAboe21VXmdUXH
COJKjjwwvpakbfu+TLO3AX/yQvj59iD5lf4Nj1WI9u69H6ywLpwwmZPWBfuluzRX
sXBn2lGG6ra6x6+Oj1GIjt5scIfqyHYlZnT+tNmDwsMerD61CxMhF0uw/aV8jtXh
pbdDB+hgXBwrxlAsGO4QMpPqinBBmYHzbcqWfkVYbfiWQ8u78wIMzxfpb73SREGC
yxApN04YU2LIrFV9hMZ6Xg67cXwplu/rL1agJBE6iaNz9KW+ePdwdl/7IFhLbWia
y7LWxoKd0tAgLreDjjDJzgQZFyMKub42wBh7i3oeKwKwvAkunCah00RqFe+b6dlu
Pk8qsvO9XnjJ1NQuw4JGvkjArvGhl8GsMaTg4isjbLQjU80fK5l3XtKgVJnrTD/W
I35FgMV8krDbFxJYkd3bWSCngreBcJ+VA2ev4Z/URdwMmZL1GgzY7stq/Cq1qvuE
dNCuwkYPHZBgQdEKWDbB9QNElu/ebkI954p+lpS2EZdB6NJTf8GnQMzvMskLZHLC
fJgmqoSjDnTBrWKaqAkX/1tVdR1uYXi9FLJT43fmJyu8sxFhWogWx2Vd9zD8h99D
cf2RtnFxzDPYUpfqfSH31oe7vSMgai+eXeSuCdDkW1OKMZn2K8Q08aOoGvtnmv5I
Rnx3fYYXhp5wtPt6+yDh2TYA6JwGryDXjdoU8Q+MvzdEXvDpQIc/QEy6OjuOo6Wt
dBO5cH7dw8136+aZkEUszFGKoWCoZXsi6u99c4kuRj86EoT8hzpJk3Up3wKJAtBV
o6JGWpE0YKfy04vYNRZsv3u2JiMrwcIMHM0ArWR9hXmE+cQxTm1BAJaxbUesRpVp
1uZYsDovTBBdFNAkdfVTQ4W/3M+fqbL+7hvFkhtKAdepoRxSweDhM12zr0EG8VOG
/JQ15TVJf1HmIIGbDooBFsSTBXqwtToB1xCYiGYZ3C3S1iwjDu47M9QzyBe9Fa+V
1vKI9rdCFrSbgPGueOoNRnqm53ACjwhCXTFr+zidiCbxH0Yep9EeEQG+4JyWwxS1
Xn6iTq3MijfOmVV0rNztY3l70iCjxIDg/ce8t6Wq/oEzqtmgV5LDHAE5t68s2wkm
r6sWW48CYO6xAPM31fqLyQ70/tLqrrvL8VMvrYSqmGCuwKon6Vv592uAVcvPJ6rF
//fSYMzkAJLFpWxgWmmx5EV/2Vdgc1Xu1dJPTG3Wbs+m5/Xgrj11oepqXM3PwJEC
cjW2ykZ2ZsbpQkhyW0w7IQPt5HG04WpPqK5anIXFAjl+8hyLNAREd5jjL8+D3rvi
D9DCW/6/X9i4IR+lcsVDyR3byXklS9zrPuiP3GTqTkQ2jZ2oc7AO01wyLWdvWmnr
N12ZuTVbd3ALN8n8kuWTPsa9Lw+C6v4K9+blkGOALwa7VWUvmKDS83Z6DfMl56Hf
fqlhkAod3oTETlXb78Q1cbYEijfZelRLBqfjtv6HVJdT3MEx42cjoxb5VERSz8Wg
UZ/N2F86n/o4f/1MhhWhVs+3FKuILjcAVHL6JwvFbciDDxyFOlsQG/XzrUSTi7uw
viOfvIFdUKZRESP+nPFYHgKrCCRudlgrFBB7K6+IUSa7Nz7lRJH278JC0qV+QPIo
ahgA9juDlug7xotkosAB5jZN6Tgfw6D2FmOC09Jwv0GLNDQqlyrrAW8P2AZEdx/T
QbVkZRCF7A74oU6m8f3W39NW7ShMk1uQgHEntP+CiP4Pdhsx9aG504iC4ypeWn8s
DOik85m50yKeXYq0ER7jD8X2vLFZ/IMNu0QNsTgRCNfQsFtmex2F6yzQas08RQGL
Zz4Gaq/PHYjkZGu2sQsGkiwur4ekxJxdxYML1qUFbBTnVgTGhZxNwTbDbpsllHcU
OdoA1kBAnXcR0bFjcXzHS3Tk7XOFea60bIRi7veH6VmoYaNEwKbcp1kqP4H4ahz9
98IS7rXiXkCPjCxEEb5FVgFwGVROO/xX/YZtSbtOJmzkrAk6sIQ/WwHqec4qm9Z1
TaJuFOgYfCHWhJx9AEJyeU7V7XglDdaBg7DxVYCoa26cwHEjgGDk1YAjzVMeI+eV
1/xE8Q6jlKM13jYCNYs+pN8ftFnztSnTRaZQpd3uMLkZAdKFo+xRkkp6rJepSonG
BbdCJNmEFIi6nOykhpx/cJBz+lNotA4y65j05dUv6I0nGIMuZPanExGt+szknXNr
s21P4sqho0kyO8Wej6tnoc5BuJPOLYU0lKx4y+h496xEvldduRV9TGrls43smCb1
ywIxjq//dwTHiwEP5xRITtgPB2ayD03J7iDNYtn2LlePu1NclNw16FzgeJ1erMGz
t4xMWmQqC2bQ9z0h+yiDlGwxvp4hBk+PiHbj9JyMwMN0cfMCxF9uonhu33qHyTC9
43dUjarHwKetXqb3P3zBEiH0/7ckIuEUP8M1SBtNypVIGooMN1qC0C3p0odeZgGd
bx93Go6ILVa5jw9MhTGq+E0pVwybE3XYH18TpGEkoagAA9MLHvFYozHeZLHRyM6t
dK9hUCTOteaL69z9WrC7fkf0VIDahZzJeavM67KkiI4HH0JIBEmAMMuvkMcsQ8Af
dUVuQlP+evzu6/HRmWbataDxb525LT61wG5LAGyy2PJXU2jkw+BGcs98dSWsrJS0
WaxP0Prrsri20LIGCAV+K9V4BXdD2ldiFJZT8n8ZHzPl0twq97VHz36lqXbAOilX
lpe4P0cdbhOvVVIdhDVtz939wEFsAkxIaUibMM3XS3f+IP0H6zaYBXp9h8N3/ADY
nRdbotyVjvTXGvfbwtqQSbNbGD1O+itunnl9xBSjxefHQYUXlVNHjeRfI/XjEhan
cA4grOM+kUxckNz2RPk468vwlC6BMQ+UQaoqwuRte7iCOYVOn0t8osTPROobNpeh
NNq2uQeBmKd2Yu6VgHgPr5/XntcSXA8e6Zo7pev6+wCNrx871DPJkruEUrugZ1h0
hvYLMEmKm6AXta5OVLY8TawyN+W4FdBSFb+HS8N5nL0YUCajpsf0tRM6R3RCthtE
C6KyLT3FUzzYGMift/Ru/j5m68zJJHfYiJc7qaPQ5BnuKyfORb6MzbvJ0pKC3jSF
Q0j0RpTNhtsaXj0UkhgaJWHP6uz5eNvgdeRrNNAnvS/nba1e2EW2xDr5Qy3biKR9
cNh7S/0tSdD3zpogC/ZBSs7GvGntZaJeL+BlkvxuwzNct6IL2Z5bA0Wb2VpBfEGf
xYWiu7LQ+GM2X3kn7D2KjDl9WHugt9mgAMHr5K2zYgh+P8BQzvLbQXbulwRo7pgT
HoxEh2/+RaaU/kBZiuXIbAIqgQJExG2gnsaUg1Rxc5s0JGxGdhZBrtLFNStIVvGo
tJ3ySukgASxDm68XVdekTAXGr3pZnd9a6XIUPYdQCsvzS6x1Z62G2AIBJ4uuj7MN
9zSymdwfCEUjtupNZsOYyupWZFNb7f92ZT3Y82rlAovQhti3shoA5EB1ahAiheH1
pGd21GmnaD5R+9EL5ebCj7FAVcQbXNKy5g9EHVpJLJnL2veR8Ob/2+ToqX+iuaag
TnZfeZStZLS1qiwP3VDpkrV1Z9Hu1NxJzhY/I7MVS0QvxlLT5x5YzP+rECEZJkUP
IPYtp5d42KbjI0L65DwjbVPmKARWpvf+bJ0QLTkaR60bXe8qtzCqf8lGPDN2XxM/
scoVpEbKKrunHz7+5LAxgjRdopP/SmY7dpwJK1x0aoOrhflwe3JS5i+RwepO0zSn
yyo98qEKWXkRGk2Q7gaenEYU/YA+RIeWNXkIJr7/8S/fi5iCQz0xXGoAOIte/lOg
zCN7r32mIiSw0uRRBoBvF9ED2YFc8B55vBEefqH33VdANaAGfiOFk9KKN9JzFdPR
pN1vwE76FrLLn/+UvmKup1fmQJ3skDvUb0yYTdXc+ncCrrs2AXM8JWn8GPZ3BMHZ
DksiIvXjeqVVWY3+stYTGdqtW8fLaSJJXTvol/QVHcJWSoHAHQM/GCmWawxh5tkZ
R0Ibf+8MlZ2rUyht0LTBanrx78bPiwWDQ4rOt5pHznFzjzD5h+yEmo8aPaNfbcaK
qe5BmbbZw0ZfsBosPUEFCIcwi8Gi63OkIqvE8aNsR1zp4k+X695iCEc9AWLRemeL
fLFzwB1mavlbfCyfpw6Fg28huV/nBRPpSMV6vwgy0xEcgwmSan+tOMX7w76VoIxH
IsvMc45iiq42ApvbwgM/ayo5hle4P1j36M5YKCUDusXMQzI6RMXVVac9YzlzMAaS
oYeF8WzALNsC1ZAdgMuEELBFDDufFf5puojWo2VAFiSr0gEl6z9iHFz3nTxn50IZ
+OJEz6Sj4jYb/Cj561DxHZHKLjb+7kZZ3qoaACClX53FuLxHbftXbiRz8A/APbED
QZUSzogI+LnCVDda/HZiixVis4mbzVPes9da61VpCsia3+z36zbnJ1ey8D10XjTf
CUJs2MpUhweprrw6tTXBHZb19tHiDMJYANhrjI1wm93lBM+vXjcmhEINo2RLlmsG
OLrQlJPC+cncJVEZnAhBiI67OvRItppd/9Xwbt5YL2mwtBdlaxPClxz8FDtHRjWr
UKWYrbECsfJ3bg0C6ti37saaBE42VJrnVD4FBEWcLKN2++8G84nM+6gLS8S3NAD6
4hTLc0PnH2QP3botNC9CuAGzmEnBmUjNM8uHXqbmUTp8kjQEUtfMwe6PGAEmL8h7
H0IX6sQYNIEezxrtd/y+OvuPCVi95JdQCWZ9+I99yCPlkxg/W8tLDzwRS02vujOc
OPd+XyUtwoagWmS3Hof439KJFgXDU9qhKF8OwJ82Lxqjt5tPIPSTeBCeoab8SQMf
R2EoBRzbHsvHAxFb9Th4epDwyPzgPGqV/Wrokq6wKxKRWLCpiiItrvoUb4MYh2vD
W01Nv0+0PNXZQOz1tTc8dWaMw1Q96sOIo9uYNtOpGaE0tx++D5vlHb0mQqRuLbr/
wc50pZ72wEedLG9j1cCWKY0LTnY3uQyE00/XiMG8SFo+uFU8fSFOZ9QoCuxCMr48
/nMgSccctnXzlCcetSXahG22bHcBQW7XdEisr/guFE8Iy0RahbyFHCsw5k2jHjnb
xJBgYBjfJeZ9x0b9qXKKk0VsgFuw2mAObP9pWkfpUPj7VUnJe3WkB4JkNaSI+pSF
R6XByJAIw3XMZt3DIQyVUw+/HCzAOcS8Mv2RBPQFdvVP6jvFdz1yM6WiThE9jEom
eS3xU9eg44oKE9T0vJY8Y+UHQkpTqsGGYiyHSLgAkfM2lVsaSyltdZm6e9uKz1hA
mM8N//JbdZOWaBtLOZLoK/fp/guDpH28Y5PzWHvafifb1fZJHTNpEJa2Bxd/rAIu
hyDFr0pgRXHVn2mBd7m40GiuceYmfNIx+/GH4mmZqHrISg5gw431Cs42v8MN+R+Y
kTfB+g7UBOM8RIJ1JzgcpLzjVigsO8IH8MnCYmFkrlQ86yXLCbLWVzqVILczjaGt
HQpvtIrU4/3MBeLcjaxqXnglnFiMtO5JNe05q3XCcB0dgM8ztsQcCi2FmQ1lYt5W
x0+hgYJwsSWn7Wqb0mjiHB2EaQSKbm1Pbo2meeBYy3o+PyP1KtwXnFCuubPJEbae
a3LVP1ooIc2PCFbLwE6DIuIAh+mpUDWXOGOmItPWBhwENAZWZ4qAKtnmRuQBrqkE
BhyfOZCfl0Mq2pBao7LStyh+k9P1x8ruuSKHK0lcZFayJROEEoX7g3JKLFRemcdp
WaByYYkAn02cq+m45hzZgzkvHF7a65ue+Q8PHl6BaWl+TObcvHs2wXDhd9zkBRd/
Opbvp/LZheDn/k+cojWlgMm1WN1vWxovTtbE+bq20Y+uc7bsTWj5rTdgz2rQ++zp
w4TTEEns3CGe+dT6XYDINB7ivApLvEkqQWjwaT1dyRpXrYTwYx3Pj83ErnIdpjqp
j97pstQveaJWAofrvqEGO3V+G2BFu9rA44rHzoVakqb6hTxx+v8NBcfW2bd3lrm3
4zqtTwB+7irEh9GNE0dz95qZX36Gm+eqths7/W2o+UVkXLXuBk/eXJ7fSYAL/xxc
Q7GHRQaiuA6OB3J8ISkjhDNbKlLifv3YH3NRNdacJ6zbjXCSGg0oxU0rfB3BTcwM
FBihBo19Y8sJQVYIEoJkidGUYBIXY2QWRPALn4OZsoFOtNsbDsOE2mXCGzsLyy6g
TYdXLGMCylVw5gL61A/iDiTDDQRY5jsUeG6gv9tpOrBgurCiYktdjmR4dWGlUKgq
tbXb2fSb30NbLs8k1+OIalMIXsBavS3cVmff3KiyS+H6v+mtiGkTJdfUErVyFiVL
ulfQM0R+RGcA779Jt3KD5wVW+axHp26RGebpFbWE05WbQHwSGeluNyYdnmtCM881
F9J0Xd+kDZzFTGHxogWnObiGdaAxCanX/FzkMrJ8RmuS8FctIsYlm8jPciimmtmc
AJqb4gSxT6iy74WwpqJ6lnhTnE/a3eP32Z05EE2hgQW42ePqfcMZvF6JMNutACgc
14Jkqb3O3a7tQwC48q+SeStM9K4gRX7iy9k9fF3O9dTYnwu18RkJA8c0Xs2lPQT8
jTD8rTdxPS8vS95+q2TZ02/ItfOsswmvaOQLpsEMay6YFwxVt/LnDvoAsM3Gnm5g
XXyTDg9PlnvT5PpfK2ujhH++NrA7oGwhIIJTzVMicO3QJsPDn9shpOsjLKNvQa75
bXGS5jyykPTmkvxJyEScKJq+Jo5BSEYOaCXFq/TSW6R2E1r+qeqzIJ29d+0X6AbM
akNmcLzV9+JveYkgU4MJRSe7iEY1Uf2t3YPz0Wh0jOAr2I0C+RWg7VZgULULaSDb
pgZMixQp2krWMMOa0X3TOR1FybZA/+KiHW5/5Cs3iZhVCWBSZ46TrnBYboPJ6E36
M95fORbGX5dzuTndmgG6i5th4TtPZ1W+wfLFLZ/Y4tu5XNNCSPk4utPYjdnhUmGl
WWreXi/pckRepbq2xSTiGdOolAGmBUxmbe3D0IRDHycHd2Pf2eTFYx6N7ByGRCad
nUpIwILdJX7oM3wj/g2/y00MKK7RkMf/Bs7eBge3VtXO7/CvYVrq0fgZN3oNlC+L
lR0Fcv4/SSv53VeoZXAxhx47vxaKPNGIr7QP10QYLjsSzBUGgAQvKFo9G/yjEgwp
lscRcqymEYf4Q5ZSfoC5vtKyFR2qH3dODgcEmCdhr+Z3+iWO5Wb1Sbb9JfrUZ3CO
25ldhlojlnVQBlqEcSH/7rJyQvN64N1iERgnmPlXkcPoxTH45eSwZjyh7wC400AQ
kXQGaWrMrneCtKGJQaRH93qISqbeBGn6kd21BOKXqbvR4wXhUE97UgUPL2M8ddko
WDimGCEDoPPSfpKpLtc0JeelhIFuoDmXSIQA5JCNgg3Eo3vQul2Hah17vKgjA6K4
xywvWZ7nNbTT+haqW60A28vWa97hKPSKNBlbsIcr5Z9b6A/kFyBNusYZ2uA8H865
E7Ut58Qjk6pR9dhau8MC/0K15LDP1/dicQocg7qTZd3iLqvfJJCYM6Ri0UqpOvKS
BUZwD7xO5VXgy3A0K+t0m1kOCk6jHe6sPPY+FvJUkTiuoKt807YTpQzzZ8x6WTjU
Uh32zEVHlBr8XfbmWn/St6sWwk2jywYMu5v+IIfgc1JwyU72sFb5bmuQll3c8yew
LM5hG0g+sqMo3CgGbFe1+hNR0A6pwd6v7tTUDxxfq7K9W29Ruxuk98YvZSEVjFIf
fPIr8nyN24xggH7VOzhW99c0kuKU3D9Fe1Sn88Zrw8LJID3KUAl2aMRkI9AvuRL2
3sb7hxOMeEgXOnqdx2ATI/6oFNypbYM/n/YwXRsNhqZEkp78p2Q3GgNLf+e5zJ04
u/H5Vi3jinlJIXGYeSOQ1jT78Otspy1U2DsFQ0ekWtZVA/N/TcSzfCZ7TvW+wFbI
nmqmMNoerSIIIR00O3z1PpF5mkZJw3QVFTOdD1LJkMQ8ILEqx3dqDwR3VKMrDMTr
TI3+y0Po8ZD0Fx8fISypVKMksJCS3GfMy3IpF3HHB9Gk14fa6M9TpJVwJkKztAcC
wbgwj2D10pCUrTJZ3tyafCS5X/lOy36GGmVbBGXEKsisYjQucmlD1ZpWjS/wa9ag
+LLGWczDDPmDOxAEf6g+Wr4U1rl4FH9clL3ms6PRflLgtRZPbLCExXxv5b2ms8/J
olksSeHNpZu/c3T4hMRly5kL5g9W8AKNCS3OWiRSkaZEQQ0IaAo3OC5gJd32WlOX
oMYJuK0BivwAr/wrnRf9ZL6SXNR89IQmN+dkoqxyULAZ7Ac5B2wriJq5Rd1VJJGS
2by50V7WRzvVMhLp2fHizhXsXb16ft+3/E4lEQE2U2SCb9+0rYu0ZnRyaBYVVHQV
AzR6CfXvpzQlxsaYmsWiAm76VyZoKFRkBnh7TOc9+yCuidtgF2tbTKyBuyoQ8Jec
KCbXMxs6sTbbOJ92Fs+ipiwHgQ654sD4fHeoI++c2XZGcKex2Q+RP44xnVmPyryj
bSGm1Rhon9ybVpnfxDAFsoJ40wUT7VPYPAZxEHe9mlmmLjMxrpbqQO7/Eq0xIrH5
eCcsgeDO8xO3UnOVcbz6JLhcEkBBLyN0TWGTkDqcPBIQtcy8YGSkebHuG15psXGG
e5ldjxe/YR0xmMucPMBdUcxnKMzGUz+CB9CkC8XQwRCr4GC2LPZWk3i5D8wZqnsJ
nEkSPZnHw5/12fKU+1gTkgpNpnZRaaucyEiMvG6dF24lwg+v82jFN/180HoDOGRu
jAW13rtaJsjJTZXJnkr8Bb7A1LOZZLxa3gWZsssxfH0kF0IInLWPgOzQes++NuwX
RIyvq+Y8uy+1mU1zxL/kpGmyAaCXYNgtQYCLx3vHIghhifQ+/teU4Y6QyeflIpbA
wPLJFEvAAykSDwIx8N5SFbZnEtFfUPleSL9gyQrovHG5L42Yo1nchK1u2yVwv6g3
ODDD6FRyaIuZE3mYXzzKhIjZGw90kHVBxT38Iv9uoJpqOfOu+GllqMJD5lD44qhV
CiJcrvV8I9jBWttD6xunIMKuMs7B93lMXaJJRsXtUYjoMqCsrlBT4VOBuBAjVNd8
FC1tOvE+SN0GwO4vDvd3o86ITVf11WaCoybi6caMONvh3JN5LY1xGGKttqeGcbr9
w7se04HXnCT1zhwiK+rF52Ad4TD5kxE6HhmGuAxMpEBtu9dqpNCroBINUE+BenQL
rS2bswOoo8x9mBr7HGdvmhIXE6JS7H8M+s4/jiG4j9CmO3oiNg1Act92uzJgel7c
ETFLIjzA/ECMl5mhiSPsI6CFsPZWt4u9PxjPD7S4x4xCEx6Dvg38I/J/VpnpyLCK
d6bS5mMjZDSMroPkEeUkW3c2b9vPJ16Evr18q1SwG3lMe7BYLjHMBJZwcWRgynLg
oGrSztrf+XXFQ73QJ6n9YDIlM68iwsTKK2z5m1on/60m2sLJuZVG6YyNUC8t7vNv
SdC/WEtH9Zl5T0TEtB16YI36/ptkEYePIl1DUifA0Fr68c9V0H4pQO2e7ISivo3s
NzdO3jIMga2vYLY5vV5icrhz2cg3OSSgnOcFpj3gl3GBwuRwdYTjGupEL1qmTPwr
F9fYLmYfpW1EZZBq/FOK961X2KSuS8s8Vls5Gl6QKKdB5+YNAdF2O/D3mT1AaMRq
vpwl+V3I3t48p7vW6P+79EvU9vFPGKST2kuM8Zs8UtENlq34xlaI+DRgL99uNGto
YXhHx8HjR8ZEEdfyfstvqyy5v16DmECYTM0g2msTHW/mrok9Dd1wvMvo5TkF5JC0
z+OD66gwWQb/ZnsWQezQAMbPHwkP50CrX7DTgJ7P8TSLBd0xqlzXVCtpRk65o38a
8Y6gjUFfBOjhgWOJuvp23W4IoouyRUDW3kgbeGkTvJeu8t+TKvrc/Hh0nXVUq+tC
fTHYDS8U9Z8Wn6cpkXZNOkv+/S+QOUXDAfTNRts0LApgvvyWpS9CxT2Em2hSFMJW
sNCDwC8hci55Obk80dEc8ciiOvNsri8ku4VN/e4EvtCTmOt2Fqo0wtzdKmmxdkm0
Mn7+UaLGbbqF0TFmtmOFZwpjQQQAG86XSbkBZP0anIRg3PzCpxGkJwXCgceDsCuS
FVPq+6y/mNywPtTtnBNyOOr5WkdwAUtljQE+zyVrFKq9Pe78THRMbqgwExCT49OW
dv8L1Wy5Utv7WZv+tWDTgp/gGgfjsAOYp0ZM/Lgxii+pJ28TOaqClqu1K/Iifm1i
g+yEARlGJYZ6T7kaNVIx3Wz4owHEifTBBDoLzPCgXVq6gBalJJlw6zUnRqdp+BRG
2g3fr2s3Ig+xHvh/eZHMYXcHQMu4p7IMbnGNoKN5HZq5zSXY2SRszsNctWKKN24m
KlE402I7gjeLZhUG6EWLd4k9qqXafhdIVAHlttngiox6G6pPPwYVVKm0lFz/4Ogl
XIHY+bExWu3swUDhQpba23GcJh3CoU0DbvBJhwf3CNTaeJ4y6g5cstIHDesqWqGO
hu8JzO7DmeFYRQ+obHxwBlJoIhMK1sgwGUkoxAjAXeLIQ6gMYnrPkryXKaQuNR1N
sQsq5iu8HbsvWYEsHC3X8zGGIvDnkBKDSU4+qNUqNqEEx1NEge5DdIxICubVEdwa
VTR1iXBQxn+umDzhfAcetrpwmFGuGueo3cgQg96p0J4mYX2/+dG7ss4HHLV8xO+x
vo1tjEhGhzj0965cSfyBFBcKYfThoAS+GaCoId0ObSwZnduPr89OJpkwBexGfoIS
/oxS8PMkJGAKeeVurXXMVeTN1LeIpEQeaIF75h4QKS6YphIaaQOmH5CTu1+qybna
8FZ3EweJvPhTCp4eafBGZ1AOhNQdSD9g304QMKWbBQ9IDPx0QfcrMjzxbx4cUlil
BVi1wrDhBx6rtu/epfLW9VRcXIJLblO9yF+/wje20nOx5aHZxdG/k7rCH8fW3SzB
7C5GsmE9XwmVUI1T7sRscYfvWUszIQp/XSfMAkvQZURTShZ9rkzXjpCNxcnhTMzL
kOcHnGyA8hj0s1BAbvm00vmtAU0lYCU9vCrcjK8RVyl4vaeJfkpOUC5/3wjjmwOA
dF42rvbDJaEzF4xRjTCA9l/GroJGMQoI5t5eSQeh3Kz6/myXzN/LNWJP8vFmPYTl
/CeCsmfjy+Ike/4kB6Ks6voL3E+GlLbVE0r/5IZXWIQ5LUZ3M7TQTmmwOUOU9SI2
exrhZbjo3eaa7m08ThQgMHnDAEVvrbpYBiWWox1LloifeSohoMF03oDiI+M7uZIC
RAofE3E432M1kp1FAoqS9sj0EBLTNnRTDOodq6slezcPkmC7uIn/0LmG+Xh6LW1j
waG3xBMZhQn5FqKAlcQowTKLj6X3oa4fM/tvGXe8xosiwpKigoCzCSfDlm/QWahp
o4snUW1uvmljDhnAszlEQjpUJnqCmXTVp8fvMFOsSvhpyRzlKHAOzWJpXWaISONs
XHuP9aUF8YebfMo8OBPhFvw3Wx7luenb3PkNmOvoPu7cO2x8du6Cjoysm/p7V3cP
rNOZatCloD6jTwdVBmvHeMszMj0AH6k87kHsM+b6uPTgYaThZuFCnP+4EHmvqGut
P1gYa8LBDt/gjlSa2uTJh6remDYu/XMHV+88V5bGAdGXhIPZqaRPlmbMEhvUBc2i
0PVMK+TOLhGb94LZUqiCyC61J39jA7vO7C2tU2Q+pswWFQWVFswIGOQXA3NtbS85
kJ49v7xCyP0EkLOTyf0ZKAshaYVrb8/2tjwpnqeXQvKygGx1wiQWIGKR4cOmLpyp
ZQFl53NOVFnGL86xeuDMfmws4EaU5/oO7e+elka309ZxL1FonT2LQCh0NOQ6oTw/
j7ejku4Vj2qChqaftp4mlk2HQpVkQnn19OSpTy6gOwA5Oy+O6Ds38xx2N9y5ThnZ
ehfPmk466l6x/Ytpevo36e8IV1TeVU9/kJKULC0CTro/sVNoijXWg2XHE06CK95+
loEFtLu/y6Sz8XIBw+2Irf1RRF7Y7kWX43VgP9fTIadbm94F+bsrEV6Z+UBWBUwu
I+UamUFyUySpkgptWhE6CQxsTTu9onABTFCIZioIsR8xjuELDWv095vKHGcf6JT4
t86cCafunh7r2vZxmsEW9K8RYfvzliHOybsHqFCw43A++NYE1tIdB0TLegG3x8vV
IRhQ6iWwCif7/b1l3c7m9TM3+5vIsecsLpgw5bWqcaKMOldIK+a+/zWJIwIke8Pp
LsycA7XMlzCK1EQVtnxtjFheLdgPyf659VqtNSqhbFXvwE5NFnNz0arrJ/LWfe1n
T6KFijmRobX4SArZAPde7W040XZq+fX88iNn/YUrw0kA97eOgxt9htc/hc1qInB1
4R25cP7a0B0Ew8kfhiOrntTjw51xDXU63dt5ihJ+gdwBCBaBFYYtjYVSvXdwIlkn
eNDs+UcYO7IfXYokTHskp3Cib1OntVWnLPCz0Vr50cOaEmnuDaHyUGPVz4e9/hZS
CetW2zP6hzwMiJI3HPIGHa72fuTizmOQqzJVaH8a53kK3XuraemFUi1iuibyQ9md
B25nZFQczfG8HFywcujOzfttp1RCIzQPYvFvLNiJtq0Ykpx1A4pd/kUSGip5kywn
rogbUVHAGJZYUBMQBo7P+NneleszVSfIQFUgQnt6rBmUI8CKSiy5c3QMuEQTc0UO
paqCv81neCTfdyD5D7PVHosB0JSN6JZujGcu/bxk3qSb/7aIvUeoi5f65hfSA60z
cKESgKhNe8sYHi1JqWafOZBV+HIayTFhttGzvs8/ERZ/oWgK1IEIUgyeBysyA5F9
TfK8NeiHzA5p9ZCstrVg1AsinXk+Dx3l9gzkcicydHVF4r6KciHPGZk8ypkYCcQe
G6VqJ5TmLS0gSZcHgbdXEJcNxU/YY1w5P9ZDKjo9O1Ym+QZaf0Ld3Dey7A62VItg
fGfI/TAx6cyiIsVzAxNfza6XGB2ggv43600blV4fY/anb7rAxTpaq+cyCmHGuhhT
tJ2+5obs9xVhnBl+AUSu1253oHP1dR4T4H4yfAy7n11VGREikB5LNql5qRxPQ6MJ
e+hitgttI7eGhwjMJcmTpNEkFuyuTRB8lYncBkwtvc0gTByQAfwDv+xWEl9Lyqaz
61f3v+XrlNee88slfBqtoOLAXAKP3tkFWqjWnpgRKYaCcX2QY623MddZTAOeyU3c
ozuC+1f88NMZokL21lQ7W8GFhG5N9IwZ1Jmh0U296PlRgVPjJiF8DVjn+4MJg9ET
C8hNyKXkW+e4y4ycAf7gXctMa/8BYTCf/yeZCX16jrDLd313KOXEEP5oEZBdB3JE
xF0oTd/pcRvTz1VQDeUtIRMT5q7GDq1NuGUS8cchPdAo6uw61tXT69Dw+TzTgg+X
C+hlt5hpVTIw6871jw8/LxI2+qVuxdA3OpG99D3aEEAL6GtC6BPI90YMmcG666Tz
YsObVODbTpCwcwN5BinCQk2nMoz1pcC/5txSYcsN+igOpJkz2h9t2pbRjG5A96p0
NPMpydz5xdxN5ifl31iobwqBhWZx18VLg2VOEjqx+YhFrCBeMMe8D5YvPYzJ/Il6
3eHWrs8/wxfzKVH26+GbYK9DhFcvBVGeIR89llElxiPEFV43CqPhij911cLZCCgw
d4WVuTTKsA0GtgjKlsNG/qctSLCKdkj+2xiJTGFGS/k6DfFcFm4+G0QvleOgHp5x
rXmyVr7yL7GFqktlEQZP6YMu82n0eoEhWHEIp5f+ZPmcsnuRAoSZRuQFD5SKLetI
nuTDQQaPPJJIyv2STSHPe8r0z7Stzs56PJhVrAyLPaJhNAfPbho5/zEgBo/XPu42
o2MxGnV76ayb6kUgZBwjMQ6M9pDX5tMQn6Z2dQbl6+UtGQf6QVJdHE+RkeZU5EQx
Ax8+yYBbWWTr6PPpBIn44oimr1y2WzzXRx5UJcalh+FDFJ6JHWRiiqDXLEoCvyRx
/0gNWvWv14IK1v8UH+EwNtWXJk6JRrypO9MxfeDhLhQ4zB5RoWfuC43emtAIU15m
Y+78x/tQghm1MxVHSUFl0fANbLFJhtaY806BgW/6JDp+VwtCG8ZiurD7fUHxiDhT
aZVwLDIxiop5cuklKcQ9cmHPEPBkvGu6sRoQyPy4T/KvJnn3C0ilJEdKV3/fyZWS
KuJGsdBdNP1aFEcR+ssb5baVCKhaz4V0p6htldrzHgEEJanADwV1+IcAsTQOY7Yt
/jlyY5/k5OxR5pbvFP5pOEWtnUXEWeLP5wqietRdeW5GKfJW0OfNyU50p4BEsvfP
SmipHhQezFBmnCj7KNdbRZrTakiBYJ7CBnqJB+PVGSudxiXJxTjXdZjgGDAaAIhz
uX6dzEfW+BnS77yYE6v6Pqnei/FT/tUwS2jhHkcNDT0k9m1gJDBZR2xui65AkoM5
2CAQ6oA6vatLeUUNRI+PO3zROci17w7FqeVFHE/8GYJwV+UCQBuPu2jIfMB1NcIu
qxdXOA4TXf6MptjjF+qtFPVg1eQTq316HgSi4puGoLTzOscF80NCh/8n5eL40FlZ
vQbbxX+NEBp6HuoVncFgLD5qTB40/U69uvYo4VahGy7clyUju+RyyyadbdVS7iRv
NQ3V7BNfO7wDQ9jU7tmqGLDhyKRc+dkuvpkA6wIdraK6cE9+dmfGbbOuzTSxdczj
r0HnHlgwuecaDI0dcTSAveo4YfZx2J+RmKMq4Rj3Jw4IhVYLFJb1RjHxVWIZ0PsZ
5/ciAXcKi+mPnD/UeXRhI8N1rdtx2dKI84mCnSESdpzRecrCWr5+NgjvaXOctGpe
GFuoMq6HWJM1DNXuDN6C3qGFV6QVp5Mbp4jd17U2JzlXoGtXUplpNdCqsUNyQG/X
AwEifrEO0GvaLXRDflKpqBGe3edQ7OH6B5k4VMMmPLbSi03J9EjleHTBRwK0GRXg
365y2x/sEfDq7qRcPriKlXKVdGElfU+CEfL2ZBTw6cvqBkTyDU/VyLfTMS2cUIPl
NOg7Nhd+9/V4izxssWb9iX7Ev+XTtEi4CluHU62b+LSSxzZ/Yr3mf/27TmfpuuKd
tbJ5WquWjM8qswAM+t2BUwVVhvWN8AlHQYA5TagwSPqx1Y2Ttb6HuvX+e6kmtWKj
8Qe+pX6cs7ZSQJCvQwDYjmDlkwQnjFrxxcFjeExn5j+64w2+2SszItdCSrLQyupl
zjBC8q5NgzmA9CvTc6lXm/Z3IpRmwurg9kKseMoMvzQO5nlbhCa0ZShx7Q4CRfmu
o54kiwTgUeJwplOWUMaSbCTiCiBu2wSTjUWRLn9knhvUyM0IkIxPMrwXW3AXYEdm
1drmF2BJnUacQfpyVtDYNtjzn5GQPnAeDAbU6dTVCSb1F+FxuUYYI7HVNwLND2V8
46HD6bzM7CQNrtP+1QQ3NHo/5eUqwfSh4Vs04jPHRoSXyjAv2EoxVmoeNPHGNIxm
lmOiIh2TfIHWzpu7QPPcpl+yI7A+4IS0XuGL3YaQDzbyZAVrhMQ95WOQ8dsr79zQ
hgDlLuzpi9ON0VT+S7QxYfKzr1DBhDdM/lnFo5DfR6LUixYUNtklHMQwGAqrllzw
Zrd4T1oM+AHhOezMBNhg4pxgPj0Lwvx/DUscP6ZQ5oHlBmuCpkffR7U84MeUXQfZ
4jZZIN35gS1aRcNcPW/JSMOJJByYT4qcvV3RJ6BNneVhgq9hrK74mj3IbLg189Bb
ji86Ks33I5WPEWQrhaEJJ0tECc93NsvWK1Sc+wg8RHW5yg6NVzjeNIJK3DOME3QQ
oJJVnr8TKylGvFYd4egRzYgFEIB9n/mlkq8gBGWwu7IJ5905B5rTPYqHkBlIfnqP
9aSYUx7Fw7df2AOI+aQTtCPHfh9NfyxaZZpAkATKRji+u6zRnZxTd7/1tABL25GD
F8hln+XQU//GM5n18yToJdspCgqEBI9QZKbiicTfKXVOgjPjcowXoA+d5TY8lLm2
j/yhY4ikbi5Phn6WApF59Xctbcocl+0iQ+ZLAlASfWfry014oWBCsHEVZpae6jDy
aWeF6DSlTJeEOqMj7uI51kihytl/+s1hFwn6dEFvHw+hl+AT3ReRJw6YNuEuch3k
HouqaO8PGRRfPNboYBk0hRlliNtwIOolXA9rMiHqVxAyx1aES3/7LWfSKIDteD+5
JMU60lwVsyT90hEBBlNDgoEz223gYCqSTgWAxQ99IDpCSIiycoEFGfwrBfiFn4Mo
XJtAWw4snyz5HwO5Uveawmmc6keI76aY1TDfb0NlcToHQE7mbQxvxY3cwudCQ1u2
MxrFzAQFxVPoUjBUVZkx71KwQYNfuWXYmWd7lT4DEuhFu6eYNgZyohQ2/BLgPKVy
egSCoD4IEM4vZ5a04pGk9PN3DyMuAw7HgxPdi8xonfO6/DJhH9AtEk+aYOp6R1No
4oRswtsOnrMYXMlaXguCEwHX5HY4KUW0A/6Y6DQAmmEOnnwxmEd+n8YiB2l+iPyY
9Q0cNNLLrqihc71UQHf/EfpGgh4qXH/LyDU0e7peTd9prpQdckhRIophtJOldOnj
qepKjp5O8d2X5CcW3iewGsvrEX++95yL4ZBxivwy2ua5y9faTJ0sNmx8FWObt65W
CLIDeEVSabivVV+5MG/y/gixv3hYML//bDb1dpgQGaZ9LpKwfe0/MuzZvhTNsURf
9bKWmgau8VZDzdlggHM+8ZXmiJuasdlGM6gZyTuvNDTxtegEqnGcDfmsNl0gib4p
LQiIO1F5CUBbNoYkt+00OiQTwUpXejyEHk3wsdWf6aQZtnSa5Arij4YGkPUi/+PJ
amE8qjtbxGWLAqyHLQMEpP4Z8a0PvZLuxHyMxPUeQaAhVte1fuwgbxIOc84NipVF
gs8WIumT1po72Iy8Hj36yUuRdQpKb5uElbNk9fN9gPpd9MwYYmx2xwmUSaD3f3Yk
IXyi2v0wcEb6m/vc9wcxQS8NhBVmiq3MY8GcQatwcKgm+p6ts0Hqi0Iau045RA2I
58nwupcHXpOr5y6XtJR4KZ+bHCz3jU/SAVeY6vuy9znIlt1ZmiTkKABWMB3quQ6/
uyfpu/M3K6qLpfnERWThRIwQKmjQ4Jtz/YK/b4OOMKIjaPS2KOfjpbFoe2BZPh3L
l57oWfHWCNJiS50SLDd2yXJxIuule3atUWpu8l9mKPt7KkBDUN8meYmJDUbk3z9E
3hMrt6LK53lio0Xh00h+IZKmmnAdvUUNdxNWATUnjsLYrreuUFHK5I0HnoDUMHof
u26s1RJoCGiYcJhZIcqlNLvB8Pod8fPVH7wvuvJjjEENKN2uOZVHQ/7Z+estEGPf
hwfl9zb8ZenwNwvvRoKt5nNlXjT86cp+Pp47ZTGOUusIKio9LftCmYqmBO7qnaRM
1+CRzv3IdzDSO/V2CQFUypJBFDiWR2aX/VvJaR/mb2T0f3VaSTFyRTJIMAAB15bW
J68Dzv/OcoLRZ+YcZTlyi6zA+ZWJ9BWpDI1HvMYC3TxGmiYGnBErY6Bfl6TMXuwJ
64skcncbyK8bMK7AG20q5L5NAjn4BrqQwmnrGiolPmKXpKj0zDnvujnsSqiGuofp
hVVaIM9ZPcZWeI/wXXv3Ni78wV7xLtNib+SVdUQIfenfzbVUPnHVdtFhS2DcJ1YA
I+Hq9ZEt7oIBPELyIRi157nvYbAx+o5CUCFyx/WGZ0rIFB4vxRlwit3IVUtugeL8
XaO5aL2vDs5/EfpEazSaWjUQd26Z2CSbjO9l2BEThATJjNsthbUCMXoIEplMkHWd
0dOUknSvH+uZm/iWCLMR1w2BApWY4Ey2fdrXuR4ZRMLAhiJcTUONW289a/FBYVkR
rXatVjDZ32Aa3prcYb9DrvEmUJMSuCxILm07bI9otFyIIn1NqBeQhed3qvYN+jDV
YE4hyKWhgA7Nf2S3S04NdoiCs8rx2ne360UTsB3+kGWAh5LBbOxlz5sVWBs94i9P
HqsUIJ2DGvZfKR2gIAbwkUscXpcOSZZaHLQn8/v5lnipJrts+7SY6SaRBN/xsEE2
ETy8mFbgYlzRu8doinHsIGp2LlAHG08NjqHegG3qLWCJgysWI2JND3fQQhFYRd6c
Dj1whdcogr5iHTGf6LdGZqZvAjISMQwWVzvCv/wGzWe8baBDNksGVX4I5SYxisYu
XGXQSVVyfr6Ah7EkUnMmleblqdOtxsU924ivOHNGAS5Jx+YdoHdbSABIyxUL2qav
R75xKWzFH5dKFrdoROdhUusdX95RrS5H1xk2rqjHGwP43e1exDfSg0qkhc36Cb1m
xT6w6LhHH2DKgasE/Q5EpQEMSEo/8OrdgULGqFOd6M1lxnc8aXEmom08VEqZqCE3
PgBlJu3qkNE2MWX0ljhtuQqOkKykfJNn5I6knM15VwN7/5erl0j3C8Lrvzd05fyP
l75CguapMBhoyWV5oadQjIs82lcd586muqLa8V3Sk5Ig4WwroKoWgQhRvGax4gLq
7ZD/2YDxLhiXgv3yQv60+HmLtXjP25JCiRKfLRDIrljQPqBQK/WQGFh0vk4xt2DV
7kiDrr/3826A0leaUBphbzvdWttrfUH+/FuAN3FPcLbKGtNWJRvkYhrCVkoSUtda
8cGlyB5lANBCSARtF09LV2ojBtcOW8HjFDaJsHYCyB8JUcZw6Jtz6CeXauyYK47c
B2+xEw7VHneSLfkrelwcrrEqsEGLGs85m4wLeQTx4QB4Ar1uRyinE7zNp+eHnAat
kcS7HN65UTlf0XpXRRCSBwI+FH3jSGXxUlZYPTpAiUjxIRzohhlclnoqclRJXesR
SCb+u+T3y4USDKN4vTr6yeErGpKUfevqN8+pKTZ4+6yFXyuMv85J48gP3kfqBFgd
zpKRdGmQpOCNR5wlX8WZAeh/9YVWZykDuosUb7lntk1YyclXEqpxMp+ljKlQ7+6Q
mAbZQaXNgdK8YrIY2PvFdDyFpufNZTpg380yRo6kGfvGfrTnWO66JqUWzVRBJtt0
lsPSh4/wKfQugNnCVwuE05Rprx9FvyjZ4fOmz7wS2bFIW7ZhSn96MXy0YfRQ+u51
a+lH8NdEXU7vti2Qwo1ESS58zLNyvzV+l8oSFGFTrGzov/5ULR+g8xdYz9kWDftT
tgVfhZnz3Ngdx2YIAF0p/vuDSC22hq/KX/88cWK+2L0k4qPCnbQLPyvTCDoxy251
uBMdNTmlPng+7acHhp067jartnLtsJCrIt/5QjHDLV7Gdz7TPNEUP7si8hN2tNZG
fzTPTP8KdkonlM9hlNURNIohURZLrwbMD+HefrAKkRD7oudQ41+BAJ3DfB9+XXWm
0WSiH8INlplH1m5Y+eYg5Yi87otu0h3p0HDc+8xC3zekEW+uriI2uoPbdrQqi/5w
e2XWphS+mX4ElJTEOvkThg6KeNiLNKjnTZxasqAjCerZiJa0Bg9HrImiBmPzx1km
4RSdgmRg6PEZlgMV7XsHEH+R4qXia9Si3f4zAgP0YKS0kdVUDvwXcpGeW4t3jzXS
nu/cPRD2gY9wYIivFqPg2KyR/jeDscDTQG0dYtQFzhTB/EDi79tiqG3iHayrYds/
50B39ek2rUp0NDoYChzsqD4V9VPA/ONpzJ9+UGX1Q+doNFyPwy/+pxbMA6ea+Sgt
RBHNAvQ8I/nyfRayzutp4rWKP8Z0P/+fiHOM9KmMsJUG6oohcsdVZi8GJmC97G2d
hhrDn6+MxFbshaQaS9Mu1Rjs2IOD+Og8Tmc30zdVTcyuXHI70MdLzxIs3sxi1j6x
YTMPIo6DTedyYLx50R+mUTyk6qSAQW6nC46jpID2JuKBIYN2b39i14AxVtMsdNtQ
4s21BSGOr1n3SOfdHjGq4VFDH4Xt/xrZ5qTzaWbAAJXaEFS0xH8or8+4dv5CjseT
fPpmwQpPPuwg6BNqLxwRq3lxY4ywGa4uZp0l8+rpMBSrwGsEyElpeZIB4bcX5WcE
AWCIzbRhhjJlHlVfQzV7QRdTi5zHqfX+Y0xRT2+gmtlbMzpvCAFdg/H1bd2qXv+u
9jfCtViev8WqLepk/P56ZtBayoOLhJM4OpcR4GmvAXIX3dF9C2z77OWgpNdaPvDO
EBeOyoq9CNJqnclzsLFs+TVBjlETOCrtgRWSCIB5XzL8iAlxAGuZCp3VKFSbTcYq
N/pQ9zV82j7MlrjwhPDSqHYNGn8bNRV/GUBLphtm6Bqa4lotqDwgA58owTEG/A8z
X+HvV/74haor/1bwtf6ojVb5uCgeavRNNr+RGvNcXPelBuxn9W9DhljCSTUXAx6R
yCxh8/oGZP23/755b9G7mC+oYE0BaclAbRsN1+G9SmjjPWBSQpf2yyLWKFAduFGG
ZReg3WW3bSV4Zwt0tXDe4hFtMwgzbu1kFkKN+Ob4xnFy8kK0m9mHg42uUEXGOjFE
P5LpC0N7n6FNyOPTN2isnQcNllTIVj7sg3dnys21RbaX6nOjOJfu4GBT37aeNnbT
ewwdjfOXZbiT/9jRFEAMdTcU664CyuNgfYTjX/hk/21oKSC8mSaQTSZ2PWR6tB+q
4OSSDWWX7ajlIGYUQjfLd8cAKYIUEeZvj/GupBLylMd+cu8vw+zeW4/AptM3EDN1
qMoHgjTJ85iP3oBqOrzMWQD3Jr4l9lVM4XQBAXFpt7rjb+JcPC+esrFcqOSgVQyq
DbWpDamBDqtVQAVOKSvwHOi0wHAgj3CntgLstd+zrybiM3Jmntll+h+M50TnN5aF
DgQbKO5kCOqhR1foqNntOzvyNRdud4HOz+7mb/ptmZeRiUsPab3XqZAvp7XIlnFS
ajXB4v7yoac56C++CPq9r2st0C2rlrMbmMnb9pnYVBERetrZpjaeqRbcWYN/nG94
0quZj+TBTZ3PhPMtz0bjAiq3V/VHCbvJaJPK9G8qInRyHLcIMtYW3T9GMAXHoQ2V
+Le/mGwsgjzTVCauptOp1MOqnTpmVEX9VOyWwjd96KM5isADoI85dduzqPhPNfK6
LtEg6p5vPgoY+YkK+7v54okV8zwYY4dzPFWoOefTsmlI4DT0vJnOcG1Ol+uTLCAH
KVWm5SxfgskHBjAq3Qo0EpYMEGDzsmtZQH8QMCfBPnG12DocDuCUuiD+dogGYtmi
AoPHJHV019YRVDnYMXBSHmxGAzK516/uKJgcRR+1JcZF3Vqfh9aKi6Do759V2lNA
oQVbYLtutbRXan/wlLDWpmVBCC6ir7YeOUr+nWh2x0a7MbYnmfcpI/a2HBgkeo7S
7sxDIAhOltlNDHPLwySEFIJZIQe6/EjGTbArKP84P7wz97wqbSi9EmC41kKCbJN2
ENiADqEDLShjoybSEqOYmNwyhqvlOQJxLf/0uSCQXbDdvgFYtDfqdq4f7YTtc8zC
8HD5aOGaTGcS2k8CQ6iL7z0In6jzH+pdiNlqLh5ut0J7dCFt8z9/D8YJbVDfgpFW
mLl+DoD2jmE6bU0+W87NRNSYptsAD7LGKJgU5nVLWGg+atIVKgpHjIOFBvNz0sUF
kudDVTPokgZL74mUdieuvk7qsvF9G+XC6GBrhYyY5cY7BjSXQ9XCHWTucIYxHBbL
1a7S112KOAUoBrm+DDZzEqrhfC0vFCjU7mW5RiYpv1+Ge/n5ES8+WYXXla587G1K
B3SkNSp7eXh6GddHuh5+8pOgDp4B7wA69IlLYWwkI4pVwzuuK+50T5MxN9eVTyQ6
0PaE5ve7H/tbUTD1uBvnNHVW4W/7IBp9Tt2YucJJz+SuvfrTokMKDouqNP9pJ7wj
seEkj1wq6ewZSSqCPKWtzboe6MJ0q2pspR1UqRde0FwQv4OfXO7XY4UI40G8rJkC
pTq7ziJTEmIo5SqWXnhjfo79i2X/aQkd+CFWemVrGYcF+KtnmzdY8jjiToYH3KG5
Hnns8IooSzjkyT+RwR6rSToVA8Jp0FLnfgPQPJNYcCB25XFuoli8Q9RqO+ShYYE1
/27s2dh4I67tEdTO7F2c5H42mgnsgmFNlJAJl0Psh2IMUtp69uDuBj9kWqtPDusn
qay2sgN+PbXysBbDshZ3b0q9A3ke4BK0JdCm+ta7h76Do1jz3Ls4CTmuMR9d/ChS
0F4QbU98+ufKfxcaLTrRWfdH+5NoI8M8NMwlGzgi4e+5hDThKkBgSzcTy++UhLa6
ngJJsj0Ziy/n3F+dWhzmWEaI9ZgceiWuChgTj5ilb885ENnqH3zpSUt/fkKYj+7V
10NLB2ts0Je0Cg2FlKU2njYQnWW5NimFDV3PTT4/uXSxxbB6RUUVqRq//S88Ss1B
n1Ldju/cB4ycrKdJBXtf+rLTUmlwiL5m+F3xJ+7vsOXiOaV7mXSHeQ6NHYymWGEr
2X+UeleRnyaK5x+9CAXBwJi9Mzgqr2olrOt6vkhoyWQf+DHgl2oMCzUOAg2pQi0/
gwA7Xr6YHZkmpmfIo0VnahEAcMK9i6GZnKkSwj/aBSzTMxLKr8lzmSyFCwSd8u5s
ZjsX/Ng2ARGQRluJQZHXqLh1xHSW0sW/Bt3Tgp0c52wkN8JK++yKnZXKYP0TEiLl
TU1dHFyzt9j2+Wu7GSmFK9qatSqHSaiKa9m0ldPpT3vlKlXFQfdgxjUSmhu8TycE
CgUGzpXg1mv/fH4jBcRf2pxe8ak29xIpVKCss4RE6EQvtrg0WHpABzHLlTtyptyP
RPKv3hDUtK9smBZdloKnqyT6YIb9jDbT9O1J8+cALmkZYPUx0INzmdnyb9a89aIi
L1Ow35FbwGqglaSPHzSViyzzeihbBPBaKHuccbUV7xr+6J/gotisd72mYEEQIE0o
gFbjebSUOMGnGF88Z1GS+XxLsPhssy+woXuDcYfabld5CULbowoNclFxzU/EKfLC
oCDfXG2CYc3u88Q2fHW5K7ZFbzWGfvdx1fRpiIgkT4IV6pb16qMSAedwI7s5sT3K
Ma+RxolAlC1P7jE1Zl3eH4trIBCNPTFfJX5FSXR5QjO7M1L0Drcf6U/TR5n97GnH
XsQqzpzBdPCclu40PytQHxY7RtxD+HhJCmgwjOOJEZAdmuaSCB1pIVauDPz4rMNp
wUzQ1R1FXMAELX5tTBPefz1oi31XzkL1fbKVtUuQGOdyubKdoQYQ03Jlg2XyM06N
w0AiqTg6R84E2qYTkBpDjMD5zI7m2cULHtH8VXHDkdSQOpJZ2OOKZvPHbkA2/cop
/9ZP3Zq6sKKItIrplkCbtFbvQhxDUNZOq8vTb+bmuxGxoVT5gSwKxtAnCjgSmcys
AQkne9tL5vc3JLV0wdyW22gpUpqpwjnAQRiKcmdUhDWjmSKPH04J7AiZZODaY0PT
YCVOvsUxe0Bc2leECMCP6DuPYJfoKC+/YIqdiTtsgemewwQR4oX3ahnbXJ6ZU77n
fp+8lJHdu1U1LMWwIX9fmNhzo2jEsKuOaN3f6Yck6VziPexCDj685YmdtLamtVi6
z8TDgTWzg6/0fZWEJ76+Zjrr+eRrMeQ8MILrj+j7O6vK5T84lrsE4Cx4dbjyFDnd
U1VucK7/lauMWcHEO0LGgmIQTdCdPYNX+LL5BYCAX8bqAH9/aLvK2gNAs2NTmpwU
NGn1x38FiC6FvphNTrkgJM5n2FqzRlf2dsK5WUrv5dhJxNIHV6CnIweazZOJXn8r
JG+jM5Nn1A7U2YOGNZmQlJh6NZrpktBbTq/4Wru2rNxCSX44wQWxmC8AGsVKhyfG
RWLDv60DxHzKm7K4LkJ+7yEaVcPNIAaXxMHJinwpdVI5sBePgO1mHDfwftweOC7X
Lrr36wyq/l1har1TfSue1mX2LJ8zaIKySiyf00WpQ+v6qN/p9AkYqdhZKR7F7/zx
OEgJDRIp/u7H+43sh+f0yZl1JnpzRU2lB1fNRO8IMsFyfUvXWbKqvGnQZ5TwnT4k
e+jLktNrQK0jeEyg4hbmHuF4KM25agTcIFhche7+ArmzW46eu7M2EV/X869ZjjVT
I2A3JjYWVa07QUyk75zrcy1S1hk/yFqvDXZAu+cKDm5cUN6/39xm9KRewCUxDRhY
eNDLXBwfHE9KtCAbL5mv2diiWQIvAAS7gej3FGx3U2QdzZNMZLUriqMWQzXtJ/zN
mvBYcjqsTgNF+eHNdpXOnLYvv6SJurO/C18Sn9tQEHBQdU07sgsx0GUVcUeEtUGU
jlyD6/jSK7pXmIBK+A8RDGQce4kO5v1ob76XsjCXWRqO/p2gX8hLn4GBMdcWC+VF
7B3/+t3QnZIHpO3Wh/0567cqJZ24xUjlZKSRxT6iH2MLhxG3LUWIeWf5CuOk5c+2
GZ4CQhNtI5O+mfTe/VDSwlYRURfmQivwe5riPc7KpZe+XN12Xv32E9sfsj0yuXc9
Q1tl9WpuvdFmaFGr8zdnpsTJg/c33MgvA/TV8/qgCj7kHCFsfDVhN3SY2LEac4Au
wbByOmwF15m4JMNfnUcy+fp2qokvnN3gV5pV/rKsnzbpkrKQLlatigolK9YmC6bk
eCQmwtcEMFGlz8uU0oiBil+kDl74HHtOEvybf0vGk+uFFY3Byc7+QIHFPut9cUFj
X4xFaR6nURNF4Zjot3UOdkShGUtLso0MYLTeAm/cq6wjPqLYDVV+0j2ShV9ICccI
m91K+Sdkisj6yJ6B9jUpLIGUPhAjoqFe0XYp5t2UzwX2qnfOrnKDUhH+AOmMmxW6
CpMAVWsBaOS3D9cANlOE1+l0fpkm80GxGL9jDtT3qL78WWqJSf36vrBvq9P5uvTY
omj4FgIztbVTgDtFvRX2wCZTl762nZkh48o/kI8qodojihn2CNYrx3TStfE0YsCi
V0vaujmLxw0oQvRvnQof1J1JuuHsL6c98pW0H0+FZwBStXiisv1UgbV4OFDQZHDF
dVpjCHqBYP2wepGw5w9R0sqMP7zRTuu4nLdusQeFVsII7CEFXo3g5A3GLw2cbUKD
au1yY/dpu561nqHmjnGFjWuSgsSauXxtm6VQGlNmUbOTEw1bXdadSXHBmfeOnahi
HCWDT2MBU4LAewPJI/+eoUn25lY2R7mat/gTd7MyQ1N5k3r129xQlhgbGG+bX4td
BeQpnh53UWaGVEj/zBwHWJZSOMdpPSfvCUjT1kwBMnJT7HZg81Dkt5c8nMy8TerF
83fY2X0vSFj/ULy3g2DLopyfNwRTY3BYEwaOa6Pm0jt4m1nLnWzPteij+Akf5xdd
hzxxwC9Wrmneh9FLh5N8nlczkFY9qW8G/afZQg7CBfmspeh1Dxb5AYlku2tAiCLc
6Ur/na7QSQwVbAXZtr62dAcuGFaHs9U6zwDpNGwzumPpHzPba0/6UcqXuLJAvlF5
CgPv3CWqpgJ09ZdJTlrowak+xCj+GLvI4bu+mH1ui5f1LUeUdjMxTmri/TjWBNG+
6+VmoYeh99rg5tPY8Jn0oja64pLFKaxUbXj8kNWxjwHe7FvMj7SS9lLgG/zwZBRS
zCBv9QdERJHsqQh5E3JMROUMqWNWMNHA2Tld0Wun/qRBHo2Zu/BY+oo9BC8xsoXH
F7q/gx6q5gdUCqXM/J5Qm/JKU2IMQlyssJhGfXJY+4Rzctq9Mpq4+kKBiWAFCbvz
MeRPyv+HdBLpsYBH0jmDrlqvozgPV4lWZe1ea4CeJeSMMdSaGi7tYNVyTuM1X4za
Pw2c0pWWr4XzPDHzpneNQsZ115trvLD8hvcZnnlAAbqiNSVL+NcX/+9A0t0Uh3UX
70b0LZHfQYBwQnyleWmE0vdSJme59LJPuHZrzAASG7mJJXofisjWnCU0f/apO+OI
KOJ4AoJwDBTtiPU3kRBxl0ZXpFh9/naS6ga0w6nEpYiGAHj4SDxERq9/njfrg/4z
DDaJ1VKr4AmdP/JJSihfYOP6qDVemSErQilPFnhsbDWW+ekxdu5WRwhmFIYdjOAe
fTLoF1VwIunUpOURvv87KnoIks6DxG7U5M1wNVPH8ZxSgeSCoIk1fO8VezKDIBH9
ds8uoRmCIW/zaEK88G921op1Mj60KojO04w0V2CDsWcOOL51g0BUrhXAw66cgmV2
cqlRlaoT/bfDxl89qcOyqjnhJFH7QZwpGz0KSm9E4mXaJW2ueigJ0NSRRJKqopTd
I6Aac4xDSo4q/EMx5Hs7xUf4X9KhwO3dPoRB/ZCi1ZHuZlghgNwmrB8f/GnuqO1h
mk27dfTkSTOtKpVfV/7pl8wESt6K0hK3Qss5HIoc/jruNgnwRXiKWr0nE+cF49Xu
b6Bcszz6kTpFBM26QRGKvCC4O38bhbLBRvHYlTJwnkVmFS949Ko4G103NjdVRxSe
NviM6vXI+rShoShn7l/gjNFF2aN4a+IdYwENRUXueaSLYu/ziXix+lm4SERAQg7N
sQlBe1UvM6C7M8CxHpovbAn1jKO4+FbJ0X0o1m/g387V7/bsGzn2t3wrdUwP8oJn
T1udAiXs2bnwZqRztvVavRpbG1utcEP2XOLTmaLbkCLLwdwQk6fFivC+8YQeaTCy
PuwUQv+Ygclqf3CbROPdqgoHOf5JzRSFzoh7U3wNLYCR46WUZnAJ6CXYJR0JL2CT
AljcZdYepjMzswOCQhqXGVsr2D6r7ld6eBxMOwyfMTuIeaBP37TO9diiOhyQS8ds
6W+4KgF3lP/gco+2hkw4hxSBhD+vXOZWQPp0vvOp4g6S+HLEKVThzZtIxSTD+rc5
evPrFc5DWJTwJJ4RFn8y2El+Z6x4DNvX6+PXwt18amaPN78EGv0OOc5Vrfp7PfQU
7HTI9OZMLv7Zx6wWvXev1WVpKZaCv2UuUSBaeTBsENImRuQYTWu66fia2Bjyfn4j
w9oZNNZgzYQF4Nsldg9WgEcI4g5NK6VNN8uzCX02yURq3TvonxSWjyKiSaipc8HI
CW+Jyt91USbXfCrMb3StyaRtRxBEUreAXQf9ZSApyL3MGnPyKt2esSZCK9TwMwKH
BmFpo+ZKt97lJwpO9qFTt7yOota07zkVmCFLjc+t31Em+xmUTdH/pT7ySLLzpp/t
2cXr9lA+L+CydAJewWtyUW9Aj1bE+bwZGNyT9SZb2cctrl9/BBvRQTWRAz0I4wu6
ku2ALhvIjk9IZQ6ghLh1zvnrKXSDydYWsc6b7Atn+8fF4DzNjw5o4zsiOeHaDd8W
TEYdNdnIhk0ahkv0/k/EXNzw2cdeb5TBEP+HNyzILD7Wf4XBdVKel/n0Tce8rF7J
7HzbZd2TLtNTiCrtps9mUB3iIPeTwL4SCSSyNTNYXxk7zRjMCvY6iAo5CgiCBr1/
jV8vjxIQ2oCEFODRU9MtWFxSnzww5ve0/6rIJ7+G612cqZ/aTxWDBVfsy/DEa3/g
5PAaFtAl/UdYwwzja7gi25vfy9PcVGdV1Q/0P76UijHhX5LZqdCk0MZ67dl/ivLc
ZnU2p8hrGFkK0NBgezP6NPQ2hiiFV5f3uZK541HJ8az4esz1i3C0VbvALRFQGbtO
+qxARTWMDYTwKhk8x+2GUuNRxuZroNx1iFe+SfF1uKtVMCvpiHIcAB6aJN+jMyPF
xEp4Nsy5rYItx3jG0v6Ib16OT2s4k0aUhAQvo//Qh6dfbuE8cCpPMUaszSk7B1mW
oZQzVQRceHBKjXAdlmv8qGXdmcaqiwavaIyjL7ZNY5/8NtJ41mXYooCG5j1ugHVD
X+emHDTgnvBOCrqdZMEmHLVOfJaqElt4oSEhzT3u8OS1PUhMcGMsGv3A5g2r25X+
rsPTYMKL2dOnIoYRye3wQkiOn+8AHCnAPI49IdmfEUAL4+3wjW1HWjiWF/j8cNxm
7j6L1S5G8Mrr9ZhRqt3ned7BIAUFUYx6aSeeNS6hCCTqOcV8cmVrQxPX5kl7kJ5/
Dyo8jlw4UGnt2UgZdYb1f/TZSePV/fjSIkBqQ33rB8cUJw7VukK9dlWoRuKpr34n
M5hBX8YscheyKH231wjvn5nCvE8qv7IRxSeulUyX5MbRxIqn121cvXIMJx0QdqoT
4pBOhGVDnhUmNV7wUu0Ea/X1IGB1R86gSq1e47mZseG3edHSP3HLEN2/u/l//o/n
fdFQwU0Py0YzTXzJpNy8Ojy6lfp2e+uHyNxg9AuIMzX16ctsSJK9BrTXrIVSH9rb
XPcGPNqDsKoA4pIjlZLNX5sizeYhOxPiWB97PO0VBqMsxBAHTV4mw3E69R5FUlDg
oICNWlYdOKJL7WF2qVnCcm1ZpNsOIw5LQZ9BOXB1CohPA4dlpZXvxKkr84AIHI/0
4WbX15BjXs8KdAe6uP5xpPfnkr/ckXzE20CVHh7tnZ+vHaikR14VFpSXvEp7+W0D
9k3VNnt5hiak17gg6O7DbcwFlB7jnuwJpBs1py9ma0QqH/FuNRNxpidmVHyt7Z5I
4JAYxd95NdmTo85S5j6i8KsV/qWWJfe2gOJQD7DnIVZxpSKC9aogAv1j3U2prcrL
OzV87M/85eAkQPFpNBdaL21xbgz9o5ESP6gTNm3bvoWIz7qx1BmCdWXdxHoydkpy
QLMmOkXyXUKsot92v5RvOJDs/HBhmK6lkHT2WUIc9EX+hr26+z9A2nuqMtE8o+Uo
oWyb//k1lg0kvs6fqH82PNhU1aGb9lFVJ9FdNJU5ctUtTOzvpJEe86iMKWG6d7NK
dK2/6JYBfXA8b2KsupJzkmlFaar1fPsvA5ZB22T/h4MnRRm6WNId/8feiwf2Zd2v
Go+lePUS99kETJSuonczEMXvDVOAebm6Dfl1a/ppSfK/yRAsdyyvaZ3bcY3fR9J1
xLYrH7pO+hN6FylhhG4BgkT6ebTin1dhE3S5kYysT48DDXwH6fAA2N5mge7oEUfg
RJANxv3SrM/mYPM7Kmll4bM/3RBcmondDdrPUjx8Go77lgbkoiZROSVcQsM7POCH
UHBZoVEqkm5HCn6RH1tnHXZBKzHA0IMryYVgbVdye3l8uLpyqW7E6qrX/K8uJjN9
cVWXw+wwbCTfDVfToDD/epSkRKbFrMm/6jIXloOJ2heTVOpPZ3EK1t+ACpQwqaqp
jbbY7Y0CF/6k/tP9Y4Fstip9DI3ZwUt57AZNYHKdjYziM47LDbN91aKgSMnHj/w7
V1Yd8Gslg/5xyynR9e16TQu0vCE4VR9FyNvCiAzH6zZQcnh2fPBn8EaF2jq6219E
OWBWojnX+NaJDFYTnbrlBcceZlExD2/ilAVZ0SBxOqgyTLL6FBdY9s82AUHL0vfu
6jrjpFS9MQKVKafmU8obgbQjmak0/yJyfUUOJt4aJJYPZssNjZjlkRTEPKXGQyMz
QIGq56qxxnIPcr+XCQKtS+u/iLvtGnwo92Ffl1x5WYfhGiY/uYOfBw3/QLEtzM0r
ZXOTR37ZsMQb+g7pBpPU77HHO2/tMO72Dtnk55jOJNatWXbTMIOSBVVMAoomtEF7
U/Cw1LSAN9Ay7Gy/LxCsTLMVRpcg0ibxR4A2PeUr/f7EdJkhzpRRggzWvlz9Tt/+
Mu5jL0rhNXmaKozvFRM6lyrgHKOdXmh2mVdayVbHAkMt/diyy8/qDv0gEh0JEMQX
yBjQ+edJoT4Y43il2Jjq/vA1ip8/AFVuaKcY84zNX7+vrCZPlEg7PwzPPx/cEHVU
x03wxTxiWmfYnfxxDnlVY5EZQoKlS3dRbZW00hVkZTU9zwUkIygaHy8BNUp2D9N7
0wJgvjBs9RV16JlXz8Wfov/dEU7EoamkhOtQCtIiDiQgYwt5TTMV+CWH8mBB+gKB
ZvMZk2EcVcz+UJRj2gIKrKdvAjuaVEe3yenUliuEjMz9HonsxN9ScliUi5I5KcK/
WLm975ZXYJelAhYcmswwko8vKHrB32McciGIftSu22JPHe3VDJiow4gWZbqC1XxY
FHR7kxixv0YXXROqoTto8kvXQhgXpl2QSgsCkIfwhS2ULQUEUL4eQ27SHhPQJs4b
uJRcFOf1psnY1epBTHV3Lx1ZqwETV85dkx4ntJGdeJPacPCf4ucXh5ByKXbSpgmC
jQogZeIfF1pVO8N27USzndJgAxN2viDSQDRX0QHnwxkD7TjGDaWFt08M2hJnThA8
s+HcltXHWaII/CQ+pd0FqIzXuN0qUVFvR1JoviTMpHYysb9PIg0WYtEmlR3B8+eB
+GhSqsdeMHW8zZ2URWyMQ5e836AuI7JysIxUE3lFQl+YUWhFakX0eS418U+fTYNF
4M/hQNmTzkmsi/nubFxt4/YNR3fGqw1dVZLnz7FEvM5lfb6hOFwpBTNmeNpNT8me
3bczjbXt3uk0Upvf1EqbeugdqdwWuHw/+KVY5dH0sqqJQ1vTIaJ5keMVPgZTczj2
lDAsAdhHKhOiO68sqTrgBXApjlC4uf7I9YNrDrSEvi2NlbT+wRJQ4IISvWRimvFq
KOFv5+bDrH4qC08MgOxhyNP4lvA5AJArTUOTPd+7tPAW1NiqFrgvuuhELF+KnQBL
jNVvgMt8oI7FyfJWerSmLB81X6Nanl0Gurb/zM3DckA9ZhXyZfXe6z7g8gxMPg8f
/m53sMdMUqQDAPoMGVnLhA54cQS6i7kf/978ayJxPGAvw3NMrJt9yvCayNMVQCsF
YkthR11Whftf4DFtCNrZ4tu+/ZZ3ZoVKkMtJuVWX4IpPoK4/vHOxbEgsiRFYGHrU
PKfd9yg2nLly+gRgcp+E1/0xMcVkBWC28tT2SZmyV6Xcx+MXg8ITQ62frtf04pcG
+S6lhabjZlQfi3kgYiOVC/1EeY9QvfHRI4/Lk8S18PxN6EA8EmRqVZC44SwLA7ZZ
UUzOTpw5WpyVLPTrzds+bVexII+VaVCctquVCAf8oQxWwKrXQTIH+y/gS9plPE1B
ZTV0tfPEHOyu1LMRzADPVPRDotzMz29CarVp5FV/m5i47Qsa58L6t9IhYCyj6Zqd
6ewj9xpGnvmMLX7+81jtjukN7NCiJ1VP6e9aLXNPazjHtHCiYp8naqQhdq7V7gZq
ZtL71MCjlFBxrdE5oLwD4ttJJdrzsM62wPTc5PY/EKtKLKW69aXrOJi19oEXm2II
CQFVVITJTkex0A56dJNcq67J0phK7X4A5MgEa0oClebfaI9mQfttCc+sAeGC3YrZ
vQ2qaHUnODb6BY5rK+pvJ8Qw621r/WMLDA7WJtm3VLh6qLoZCrEtwFiB4umexF93
zKb6J+uZ7EGVdtHTnKzRN1Ilp0dlmmCRrkFiJz1wnetyaL/r+W2tr2m/7s85ei1r
0m654wC3PBtRxkPOLDVV2DWt0MnsdFF2IBdkHSZa7ki4uFnaD/2ea0Ym1bj0Esk7
hUR+7U/IFgmNtIAvS/zv4U2U4qnPsrdC7gHA7qcwv2gOHYrpRBG00KbIafM/ZLQR
RdXVWGJsvOanfU+RLUHDLxuYA1/i/eFnhSEvXnboIT1LJoSgq9FFBKlW6eGv8W8F
mFYYy+QMz7AFS6DbxyPO16Ia04rGzD9bE+o5RhWSPpylETS3Y0gOvnRP84UG8WjF
1IsGEwFA3uIStfMTHpsOEaJoq0XOrW5WKN0FMGdYPn1Nu0XyoWidGa6IAwGk07so
5xSVC4DX7x4IRGljnEMDKchDoYojdWlUgeeJwqKiDoUH/F+4xZvz68TKMeVktmbO
3d1OuNg1Bkf28GHx2K0VaZvRSg2unlp5Ti/IGL84TIMEbKCbvB5MWw2JoNGfctjz
7Dig5sGLK2W0fYgMwDkPCgxE4BNRTsjKg4RzPEOJWF1jeBS+fC4eqR0ZMeONOyri
hdJwThm+i2c6YAXp7gkhTqlpnm7qmg4w4nV0Drzz0d7exrJwMKEmZ+YYAKqMEYZO
q0ZXPb7gFWnl8Cawf+UHeH7To0keksyMcukrf0/4qZtTLRVovRVygh0KonD/y7+E
Joo4oXrpezq5va2auAut6Pgbt7rdz3miRjXQW1IOb6jIGjv9+1LIAnbH5+iuziE2
aI3iYu084bVieIIDj7xpFPZD7NcHIEz41WQqPyqsik1TVyoAqyYzkXaejoGOPIc5
pYEkRt1r8eQ+tQX81iBTC5twmjGmR+dYAlXaQ/ey+BZnw3udcqHqrK5e/aaPxmDO
wBmUbI78ttaSlPhn+vb53noGa3xfU1N3BgKHfHbczZBb1U6n11m3ZlkqfJY0vL+s
hete1TUiWW3nLKKQbtobTsfKqCFQWG+0sW999szRMM3tWHtO58l1ZrcuvPIKWC5p
Ebw/6H8cG8XGgfpl2JetylBexGoNH2PI9WoNCvvnSL3m3hxWMpNdUTKljB+n8Jif
MWHq/R6PwcHBc64Oa+5l4zRhiJxJ4VSFUX6EsQa4z9Y5JZ33ZGIMcxb2vrGG1W0i
CjRSgYoz6XAszQw+Ms1ugLEn3sL+u3RMNrgNGbVitQ5nps18BgcSRliX7KD3gfJK
3Z6iHJlQNK0k1TQmyF1Gt/lSWqKR+5HV1dK6HI1vZbJilx9MlQmGrvMW6C1D/6ZI
yM796v68tegdtys++xpa6OpdsOtnzf0Ov8AQHMh2qkiv7rnnpgPjLCSJZjd+LaAi
4JZCRm8DoUf6C8KmF6fKxiKHkf+RysJzPZxwbaRhQnZTK1LWQlreKQry21+XVOaP
dQ90+YKw1k1sBjCM135DzfN5WlpO1C34Oxd2oD3YuukjOVDYSEA21bGjhU+bSIAu
zWxgonjVUL8ezpZKLmOmJ7Cs9MDW9weGVztOdlB1/CnmTJXBBEZ+bX2fLC6IKs0q
2Srd/QiskKr2vd22ovosaGZZtRAI7dJFic7i61mo536rwI7O4xKSKRxEjruy5cGw
+MeXXIpeEg1ULQF9aVwJSYq9p18nKL13TAKJdR/Upx7enrDVh/FmI2XdRo+7dtPN
7seF4XN4ljcWhYvbUs6fQ1FPNU6qBBzkMTzrPRdgJPzrwiQW1t0EaTvBVlpVAIiX
oy6XojIua+6sIoy9zVF33kGon3GnUPY6t9HApKNZ3L82K1ulMjaFP2pcEwe1XHBJ
hFqu+gXbzyPBPK5pOOIi8wIgcC48JKtb6MfCWFgr6zp77HDijlQkgoyatf3LMPfd
lxnWFcYz0Eq9z4IKRLA07b6oT6AtwBHRbGoQBVyhV0inqN/f+2Jc4vJg8rKtfzrw
y1yPgM9IBVQ8uEJjcFInUTdlUTJkDPaRbHkekMUm1HAps4v/Vtv9BAq7/wzAVblz
ZVQtuvZKtFi3kLPJJJDYhP7X6TvKRD7jY6zMUQ1gozn47tDoz/uEqG9fM/he7dj7
TVhFKnzphEQuGNcoJfYzyZbyxoeiB7+zBkmXmmdtGj4R2wFt8hMeV45EWHFF3jTr
vqfUPcgWM2hSHXiRJdiYJeQhcG6dsGCucPRenWpsWFPdP0Yv+i5MxrbIYXJzf7s4
3c7no5k4NBiQ0TQ92CpIT7X2Ojp+1ydtvL+A24wbNWmxhVFVUvS2lb54Nj/u0ot4
mVliz6ZWC433C0Uweke80xvDajjyy8mwflB7wyuQMMdSRK8o3YSY0bqSNFPd/gEH
OJCGohXMiEexJ9w/K1HON1Yg8MHQXr5+isT1ya6WkHbYpzyGNS09QSdfrEQq2tFm
LW0wpTPSQkGUD/JBA8miC/Oez227j/uYCly4ndVf0egx2IDD+73fCgM/b48a1VOL
izvg8n152qXBlzfvAbVHwCLZ9Gg8kE40SFQnh11jVQlSuG13Hwlk2U3IxMQnODCe
7iaBpev7wsqRD23haVR7OibIfxgK1lz5w3tTFFaxNuZ6fqwafIqJ++x/w9/nOxgo
H4G4XfAf3wwt82YfLgPkzYlO9zPocmb+sNSPi+PKsiYxDYUzvxNAhC68ZNyeVeIO
kHQ7k+aZ0Dz7tG1UVYxqVA+GwRBna2XQTPBo67a5MeRVzowjHqWijVKL3Djoq6LJ
EvwnUA7df60YZeUmcHrTaRrKSqCizFmWJjnn0MUpOHtbrITZEUyb2VW9ijdrenWM
oSJTlah4ugLr9RtAyUlzrzHL90GzQYJHBgzLx9z8TRYPUQxOkCWFh/LhcwR+XYS2
Kl9qzKDgjAOwtrjRsPQj6bmPWUO7z89RTNijILdZJbashi3aHEHhlBNi/JiIoaI/
olhqqyjbJkloYUFJglziqapxwH+/MFTYOManbxFnxXf6rhk89w3xER8RbvMEH4DH
rbfJUrV0k2NFNICzWVC7Vr9S3d35HB9PmTVEVL/qRyAl51Ka7U+71yUklPlLzwHw
IHUm+k8uKomKS0B5mOrgkLV02W2GySgB5cr/nQMkMZX5IPw2pb5FoZIklBK1aR7z
sun+h1lLDcb5pXTAQ/3O74GYKPTNV/bDc5GQkGbEAT6j5BJSZOLwwdGo55Ey/dWJ
UgrAaORSP9hfXY/EgRCg2uoGEQ92aB4r8vrxFevbGZaFb5uKemaQBAI7cDOfbHRw
CYeYgm4OoBLXZ4PW32+mz39UeNy8zlIMswbVl+JRPrEAy4LUoPTnNXRAT3HNql0o
hFEs3uyTuFNOLgWxWB5XUoc/w5Ah48UKLZc6iBbmRiDmDOObsYzdSSioVvh6tcTy
BI5z7FWoDRROZELvLU6bci4CyHcx/MaIuxXBwP87Fdjhb/Op2eDx21df0NDEKL+r
bPmCL1xKldTl4ZyFp2rVPUpkskYIfkEda6ZO0SC676lwEuFupRX+opToeBCpgM6b
y1rgS+8sWw90K+TtleYTvi+WM8xC5pMqGXZJCnCL8Hyegeq1Vc+ynDiVlyk3Sdki
XdpNm0lH7EahxRZ4WNBz78sL5LWVPhz10XUyimph43SIMbXu8F9Dd1Wjl+ZcoGzK
TAxmVdork3Gfbh5bReUahybRGX217p1n1pKkX5uxjkADgx0DoBVu/tnVSLLI0a1i
DTNpygCPaDyOQfwZlwGMexqL8tFPggNlYAb+LQv9/SuMRPoZggHeOFe7YKi7ajcg
YFeIzU7QPokwf4DSuRNZpUey2T7RtTJU/D3ZBxhWWtV+xGueuRUy9IVDDKtTIC1S
5zE9f/3Umuz/N3M9ek0M9CEdZHPTDT04ctSY6XEaxM2b48rWG7fARsQRSYmSPlna
lM7KSn/8lNP72ktdv7H4T0FFfXOp80ppRncWZPTXuXWzRO4B+zkKh4ysQ2RpynI3
OZQ14IHYdBXDGika1VgGhxs5C55B+wahOiKIJN83L7xxn5xaNASXDnUyETyVZU1M
YcnAK01VQ2/q5Qe4tfaGvi5yP5EUnPWWnz9IpOp6rK/HgtP9Zp9Ffrscc2C3MnCr
X3TRc8jO5usBCg7LMJJNFUI/6c3xGBesuXhAprcWcUV2WaUSlMFIEZtWMRmLg04x
CMrXjH9MdhOpEeLc2FjmgdmgCzfLu+7nusVV7ZZPo++N+8Hz+8q/HT2zx2fa9EeD
P8KyJHnklR9+7G/31yQed0XhbdIJUmIE8jA1pDh1Cc+FSJpHO9dMghL1AVqI1lZ6
ZobZOL0VwO5EKBJ1RItD/ocSZaiOOAKncR15RDU79ofXMUvB2ashZUl0D2+4Hs7k
EyiA7qoQAnmLJMKbRoy7z1ociiox69UMI8CIA5qg3vMCP0oit/ZEapMIDSNO5a/v
m1RpgI8WP77r/tdHsVpIe+yYVPmPrAwyM/cfuo/x0disvZVfg6mIzCU6wwINRcby
bo/yJH09JqQ9dBUQZUhjpxoI8kQeNVFaSSRXovdw78y8sx15NB50njnr08UpTVtC
ucxf3yCPdMmI2UqqhCdbiCdb7IxN2MjrKxB1qx/bNsucLJRaVUodk+mOyy8iKKL+
66PT4IAV2CrbhcezHRxq5uWAYPCj5HZxZIGr+XZDeLAKtdyD23YAhHk1raM6jouz
nUCiDxtDEFB691o1bY1oKh8U/pfOxT1NoUO1IGt30gZGV3NC5e2vp0pTD/RyMara
ioRzMI2B/oT1Rc4TB6urhI9gKsJ7Gtvc/QXVOO3GaPJRqFU9t/atmDDqxi+YXAVw
LoU1jmkf+7R2KfuQj1wa1im/yLgDIPYKWLUotKVUG3Ig+JWbU1itYqZGhrScYqiJ
2g0VFW4oPzCuZk/4W17KZdWMYNptB+htriSvRroR20/OghbIvAphaO7zOm7lQ2Xf
BSKHYFotPXVlwrmew0pVjqzM4cIK4owfpz9AYForRgFAl2ASXBdTho+7IgL7BPKb
5kW25uFldFFVGTlL+fEZGLqMwrzMrcmBnRay+VOw0x6oQdc75CNcrBM41H9uUWa4
hpszAcmdTdHjy4knWJEBFBFJgkHW3IyCRMUJExreLQ7YsD2rFgEjVpvnKnaJJvY3
gs8uSCNcDDC+7NQ4xljo0nZNxuLOAJR1aPuVCT+c/I3umy+UnY0wRpmM/Frhbbxn
0Av2PovyvSiJFG3t+taoylGehsFqG5mw2t3SRlTUGWZDleCjQiZyK80BuI4jvvD1
B7YHR6T6L8koR1K3wPztet5l+Bk25b5IzSbCnILWdDXAlPG9r7K65Ld/0CiuD2yi
9uWY/Zx9Ye62PopZG0ENHa4fhURwUx5DWzGjSAh4FwNX4iQ3GKNNTtWcnaiQ6vkC
fJK8BummIpnA2hNxGp2m21AX932BvsVvTGcEzzaKRjsP2ZBWlPTXG6uCAZEFv2js
5bHZiaIfoxVmizg7Ienbtgw81knTzIo3lbFhnGzc3ukkyTREpnv6gGQfkrfM1Sim
ZlB0V7KpFbi9DBf5xdNqQrWJ8UaFNMsdf8lsEMz28NNFXqXTr3MnGF+PnOcIXp5H
VRNF08nmuDRsaNxAA8S83SyfESi+VQsfmmluTpG0K/JY7BBlX9wNId7oAiTSmu8g
MkmerxNPvHo1Li4aR33HNp6/RmtBnki4t9k6zW8dAU0X7eM9N8QYpj7uTrXYqTdZ
J2xwyd2E9W7VVrGp+Six6pd4KKrN6XbA1eHtZiwKrcNu1RJmJFMIwwHFNyDXMFiv
iI4Q+ZZjvtSIbwf4Wim6GKUU6Yq+H52mmYiLs2HMIhE9pB6j5pVphrNxVZiQA/S1
vC8BESazpOu96Wj+5bweUgR4/YhOAjMMMwnooHNIRQ/6SDTZGjKpvzg0ssre0Bt0
n/7ODf7yizHKfE7tLJ30pGagblXXGgWyOUqpwXFVRFOi8qVbPmujVx45mkCmuzKD
JUH0Yo8MRUVe448WuYkSgDkgIIvMlyzlXrqjOWu1+8ifcV2dYRxaf/pfXsMtvd4t
hGjmXnWUh9pRRt+ohpLNfkESLqTlSV3Hy9/vP8i3KrkHwCUb/eDewjT3i1isI3GI
RhcoiK6u0U6yMKQcVTeDFyrKOFgfIWuIfAss+k3TPkHereBg4p0hI28Pj20bBjlO
kAwo0yFFZJIR7hqIa8Tlmp5H1Zq3SfNghhQAVokQeFYQBUV7Tfe5wWI/L64MWg70
+uz/738IXB7kWgBMnPAx+hksoMkpg4thzkFWSW7ItwC8maItBYgFoDI9dXTgaWx3
Pexu+Xer5FUQEu+gFr5r7+TevHLeJdsKewgc9kn+m+z4CTnWupWsEd4Nc9z0or4+
FxIiR+PGtk1vzwFFfM5tejmQ64cU7RDlsbrlgLMcPqCOYaTobt3B5+UJHpZ0J5ty
YVhRxKa5yGhQ3T4h7XFxKjiddb2Fbh1F5DKb+a/5UBsEFszlJk4MZxE3K6hZ3psa
wzcXtSxYs1D3W30FcVQIwYn50POsXmRS7Sl+AZCzE51n8CRCqNAMy2JMSqkpnMP5
dlsARRFtpoE+YIJlNtKcJxsxCgbnJOnFXaydISERfad1kNdSbJiAAmfSW2suMBuZ
xykvJeUb5osxUBiULTyJ3lEqRbzhByBWujqv7a4Sx5pKle1R/wcmTLJC5wbkON02
KdQasfM/FVAsctqrJdXgYP9zxeC7QNUSD7CzZEemSaJs000LWVmKXeNqJ4II3/Xk
ag/A22o2iJtBxBPiTzuVuDscSQXoaMJopK1oft/VIDsjjLorYFLUt7XsqrFZ8e9g
Rx3ZV7DSzFtaMDuOWAjSvicnLPmDUvbFyxtLAcLtfuiS+ruezsbUhxAPtXq5bqOp
2QRC2t93WGlZi83LYqI/cHKOYg6lwWMpW/wdqI4eqauugUt0KN0xn96LsQbaWQhr
EPGEL/iAi06fFsz2eUQUErvNxm87a24ni+kTcApeTtB++kS48MoDxifu/5fB0U1T
GQkOFxb1EEI+naapFiJAPtQDm6zsuqQQxJLlIo0QzU+k2anwP8jipd+BQj7FwXmu
rXPyh7ApcK1GBmhxXsE4+KVxWQvftAi5qbFja5TNSX0Wj1zRj0Wi4bclHA3mgW1r
fD+DB8uNyOVXM+hTMoRZsEcYK+zLoL0YBgOdqwU+Pp2rJyU+TpAcojBdRJjMrEaO
trjWdUlpseCRwaSQsr202UBm6A1FSsgSv9mlDXtbMSmPQkFN/vRXZyxCCV0nPp6W
FJ3z6b1qKqkx6QQ73/F9ZnNkCWgJKIU8QVo1cz9b8vXb0xSr464uVY9zQzAxQIPs
A0nnrHM9vOq7692i3v3ssDQwEKLuDBGCftVCtrtJhSwsC6HnaXKyqtyVMfJO5aOx
8j79z/6T+cYAVkYv/jkIefey329S8OvwMJjVobiLby69v/FDO6qieIEbQHGUrqdd
VWwk8GHowTyP2gVYe2748YJkd7B0eRNE6YMQA3RyK/2hgmo+WAAra0cPMUpiDZbk
BYvBr9V0UYwBUuOtW0lgVusEdqsOlCwDN6WTK7vQib89zoM5uz815bg6tj5i9xbW
b6BD+IOaZu35GhWBUVodVMTnwfeE4wmakn6IyphUM7rh9tHPrvPPyY6xvruDs0zj
EV9CrxxCa1dDujCvFzLFyetlHTavUYcuZDbwC4539AYjvzwKXhJ3qwSExK1FbT5R
PCCYs6m/KAgG+xDPP+jBHKm9WCXFdZfwl6Yn3Tu97ZyLS/HGB/jrGvCVghsM3qyY
7u9aMILCcvrcLclZTovgrMUg+hFSb8V2VO4fYLs2LhbfpDjYWdk6CNI6QHKD/WZE
De3o69DfUo4pcYgqlslFshYcTiy5z5er2oky9C5aATgG9vQ03+rsYgHxtzWXaP/y
Mb+buyvSQNsPFEIKR4B+MZp/vbqfViHqFikzMfYvSzZF1vTWo1dNcggYwCtbpGAE
xv1hzWa3A38SwHAS0MP5bpJLSO4hcShKSqziUneqhjUPhPvLJz3dIeWQURcdA6WF
cPOmg0OOlCgBNkmIP41wbu6hUrSEiBxMMP2dixAeX+6z+FblcaGhmZy1+5QEfY8m
doa2W/H1PZoWh35z2d4DBKOMb1WOLFp97WAB5S1N8JEpKNdIWE4x7MxNQDE4Btlq
dnc/AGDKwAZEUUYv1BJSZX11unbDqouPLhCxKTIHPLtBUMOYdMZyRP5NsrEtB6t1
RNVyGY0jJdy2h5zUhYF4RtOtROOVYbrdbUG1f/JUC5othBbLZhbSv8SbZ4Vn5pwZ
U4wYeCVKCFhryBQckrvi7WKWV8QDvUipDjByVYFhuh+7ItP1mHEKQ7LFwEU5ODWf
fK3I+Sao6+THkcU1WNXksNOHTb734t7jHoLajx41jpWCME9lEJWjQbLtyJa+C2dn
N7Dep4hsqkY6P2WUKruH7x5zksy9A3QDaYY9TM/a0BNe1Qu+Ybi3uUDbgjHy7cfL
zrpmvm4WTBycvpTAGj4fnwB9DsGIe11vjcxvgsfKeNqzV9b0Wl0QkIPV7peqwM/c
Bt/SZbUPzc4KMDSzzvelKooMrw+vKERtK+WsDIH1V6kXD1inIPALwBVPwmJ7WolD
XnwxoAwJsn6ES2R4uDV0JYYzO6YJoJnVO/WD/8X6pEsOUQ1I9rBHiYL7nUgwfmEC
BVNP/eh7IaYMet2HjqG43VIweqaZGbPBrDDVuRNZMClD1e/mDMQmobroWzz+6/2p
mRAKVtgGoH5U1AFZGBpQng6t1lXQ0ZH4TAhwaA376exUV8XSqYrBoF9x22AWlya5
SdmcxtILpm9glMYJylLMiA3SPAIbuvYaP+Y3Ixc+lq4Zzx5NL93s5BICakJLtO0M
EQeEhvVnMEQUyHBfmhLFA7lc12nMbhh1ljOHzoGO5uTVOH/AyqFK5VnqpeGytI5s
1dII56BRzCb1LxEbyKUp14o9ZcdpAyCTZ1/lUr2a335eF7cV1mkeFxb4tdrYScDr
PaaMjZLqj5i0Uw81VxzWtEiZIRPQtqv4szk0+j9P3dHmmlXUGBeKF2r3MU8t/ZWk
XBwbEoSwGAr5ATGKcOiFyPiJbOr92AFHrtsffNgwkzhXAp2x2rKobJ/121jl967g
U7un/DOO79n4pTJWnELqe4A7kgM7C4zelACjCu88xL76pa9gpEkWq61PNcli3nfG
2VoaJb/Z0+VIvF3dCGQM6C3lfOjnrSfc0JEJsouPK03qWiEWd1zzRUpK19ee5uwo
4QfBzn/yeM3xR2fklwzS34KMmcg70fwcmhMihttrJfyG4LAZw0kKGbO/OCJnOJJd
FFihkaiW2gvvtgcZy/iYBHEnBJFwBunMDpHxeR/EHRI0evICeo3rb11EsRarqI5z
M3lFLSQq3dLbB9Vrs1/MHCAmdGEYeSQKGjrXL+EizGvhEkiF2DklQUnFwgfW/vKk
pjYuWxQWd3vm9sLlGR2TO2/WxkqOjEDOptpaUoLX8rhdmnga6QU/9QL1ZL7JJuJr
zHG7NytQ22PvTLRecP7Tv4cz84/9uUvlrG2bQ/q2fEiozdz+/Y6OMYvZ6uaJJG+T
jP0eFEG7v8DeNY7tBMIafSgk6dXECprhvT8FI6dF91Lq43ZQeP0dMwa1cmf/cQBD
7E1TgBQWWLfcx1ETOumirpa2fL7IdFW+iqg9yJJHnVlc3BDVGkJ4VGYE0I9XTbRm
EhNRubjJOO10b4uYVJY1Yr4ci9gf0C1cTa5lsCvwFs4LdJChQdiyy0PAgjGHaD0T
+bIfylvbgoobuyB1n4GDbM7ohMYKeVEU6bD7ZArKKMjf0/wUrUE4uaRfYPxBCSGh
8tOXGR6cNAKpKgeY+MeqxZl/7X+731q/rcoHtYeHjC4H9R7eVODXqXfDMr6CL9ym
l4BzLxWa1wSTx1E0bXGLBzt0PaO/ZC/6Mp4JhIEajc7rmUHl6ldX9rF9H58BJhdD
CCbA4KmMh+IsQU12jcSvjhbTJIf2hzq0ygP9EYOm68UNlHVhBf23Vd0Ddf7OBc6B
vJJBLcv2K5pP4U/+u3f1FmM7UuvbeoX/rx/Wbw7pzqp2grF163U+6cRT/lbMq1Sh
3OeRkitPANa8K1770k3JzCaAj0YpQIiDJKgfa3Pf789rznM0h4dJMlzMeaGLUTeh
LzKw+7CDJLewUkvVDPNFslYFLoxO+6ZQOVHAL25UYxGOgQLYmiEt7M6qvJnvCP7T
zzGdVDxLuYVmRL1So8sFeopgjs7F6doa8N9Nvojk7yR5h5Fjbxn6EWszVB9a88T7
smD/8566sQ1vLG4IDIXdYy+eggkrpda2HVaxdn1NDsyVgY1zrJjfCpRpTwWsUKXN
tN2LRZz5Qp32aX+KcEUVb8Yr7Z3YZSiHzMP6dQP1IdWaFmulH9bXxSq4YQhWuZVy
r0g+0eWlDETns9R9plSQ9O9IgwYpHNAN/+ephLNHKapBiqmz2qbnstRaOZed//WP
3J6ZuMB2lMD7vvVwacV1AWk/fRPjiENE+5k73Qi/W6CMhg5oscEUmWLRhPZEli/A
oQa0SinZUyL7DzzPWTGHQyyENtgH6F3MbosaWmneynILvBnmJoMvJIZWsaeObPTa
OGLNnrhInOJxf2PuuM8f0Hsy88CI4YrcNCt886JBMVOkswFXkfxuBR07123LCYzT
cB8PqRbCo8tYJ0BdkmqzmTIKDdTzLHNSS+v68p5nphzGXSAiFUhWrSEe79/YVhrN
h4auEW34B/apnFebmjI7wEqQ8Pha1gKE1mpJbktkvGUk56Hlj8ZYQeuLn08iVUua
K5n2gZ0ALz/MfdvjAgoAFsPiKylE65pqTKtsuBRU2p6cWqOgtgfZmotyJK95tbMc
gihlVKNSR7+dFX7kdTxHjNb80rtdDPyGgPPjyOb4pdWYHZlPKUOYMGBgv2UM2EAu
EmrF3vo7z9zquLplQcnR2u6j+PGM268G8NL6J4cJcox5rNe9gRNXXHX9CXmslzIs
d5ua8dt2gjvHy4NFiiaywRnSBVV19x5JQzlh24b5i2ZFYoTAO8SiMPFii8Poiazj
f3wY0YApTrEh79vD63q2J+c4XccH3EjLfkfoHyVgh4n15PYAIbuaahYC0Vuwp/Rq
cec6Oh/M1GQNoGHgDKHCQCwXRZvXr+pT4rxeQuTFMN0wZ9w/LUOVrX9P1xlkqoFp
VMnSE8E+yp32eP/oSAjEqoIgmpuALiPIUWlahobIB/gzKTypzSThXVXanvhxPq10
s1b/y3gkKcSq+EcdqxU4WZA+n82aEVf0MkMBHLljjsRsVv2X/4kmhqCT5XYqZtI2
pJ14tSqmzMNRV2S4tvFsN+B3Wee5wQ+JN9rEYeSSXyYuJ4EyUzljv5tmsRMBCX5o
rXlWgI1JEHwukwRD7BRvtofSbHwU23B+Q+GShyDpdKwGkYcuqZNoRcWpr3EC92Md
Rj3gaaviNGMLw15M5lyb/uSbvKL8mPR95ZAVwGjz4hVQLQv0km8WzFTa33TCg4Cz
tN4h4MYJLNR+giPC9i5jZ+Si6vrhAB1BRq39SjmGCXpvdg+W6hjmH977wyVkZoNF
E11CeznfUU0d1VRsE1V9nADbwWFDUVzACcE7WxtalpZIEWPUtrl4ZC2kYZ/CI9co
dAmMqZSnVNwubCvU5xOqOLDWw9wgmbmUvOdCAzzlrwvs5o/EDk0OYSBQDnEdQe8z
mwCCxa9eV6vTs4u937LX/TY62x1QvjPd2CFfE3Upv2LuqItU8FYuDIr/z5OYmqU9
OmaglU/AZLWeqPFrfmU9IejPD4Mdvm1KX5DoO/18ZJ8gIbjSMbcsFxvSD9nxsLJZ
/rygvOVNVP8j/YiKQoEkdIpf2eU5GFb4lxwbcYOYU1jHNg5RiglPfhSHFxyxdj4z
xT2xkxepyt1KU9R3UaUKbkzFBL7IZNWqWIZWLpCcDywsNV8h3ihmQGzTGros4WLU
34ulpi+mnrED3kXnam+6KMKfSjwi095Wv/gL1bXYfgWSQiox26uAVOT9SGVg49Pb
Ovk78ACdaW2dm3sfS7Avxz5nBbo5YdD8nxTIBq8rlXJtOyU+KAkhjOgt6zSfM603
rU0pKRnEod4iqgGrO4hn89vL0LZE+cenR2+ayhA2Tx68JTbmq433gBJNRcMp0hsP
A+bWull5PG173DVBGTqSsPLpCigIGurOwMO3IPZqaCLbByrCFxl9Fd+tJz5lyw/d
/17kp3ZiPVz6IlTFoT4jf+clQh8Xcvzj85MzGIrePc0sWcU8n8WhjyoOMkE+1hc4
d8HXJAAft0AFsCfvz2ASattRNmMS0T1b0zIxrNaaDc21Y567b3LLIAij4G8CHT/o
kNaFT1SVzCii9H7hSScdo/icld4bKnNnokIK3QZFHVQuys6JZpSkMFQ+cp43tq/l
+SMRG+4uFPCdkdrwaJzBuIB24G3muNWE/Xzct5cpKWi1t+McK7JjrdUYjoydC2jr
/wg9JdpoIjcl3GDEos0/SHFMhSNyxLRUXEBrOBDjuALRy1/8SZGDjUg1d0yYYFwu
Kp9w/ZtPVkknpVB1k1+1C9U1swim2StDXyeahb7xY7lMhHtgZl3Rsp7gOffYHDq1
UO5pz+7H5cPyczRPv32r3Zy4oAWNWvIPJyfTB1cdm1NtT8qR5BvGQrcQmzdZz3Dq
3mE5poGD9tlATgyivpCEAbYHdY8js/diYAmZDkifnHTMVvbJrk4YBw1n2tozH9mw
FU9Jft3eLwNbhggZ+Nhqkv65R+wHY//czKf9YYIp4V+Zxm0TanCNnDdwBch09G5Z
H44VRidNeDfncpspOsba77mrFPq+rZXX5JK9G9e9UkxzGSRY6A9rRF+P5g/m4Szd
55D7/fN770hLQXlXF/uh+HtKGFCZH2TIu9hlfcYECuNHFb/nUC3aSXE2NqzH6WFP
QOTVVtMgiQMOKdOIxj0rohAI7vDqvuN+2wxe7fl466sEpvZ87SD4i4sSRgSrBTCV
aOO9H3r2mzu3KZMj60at92Dozh1hvXKCP2e/4KRu/NSPihTeGIqyEVa+3DQ7JoAk
rDHs22a12UC4+dff7LhcyVPJWUjabA9PHJwNP++reBJRI1lCGWKxGSwYndJT23Hs
05G9H1SR77gAISM7p05Lly3O/Wxw4CgFpsxVP1jqhxtepq3yEo1owowaAMxihMw3
VXQ7t8MXK6CyYN0dJgy8afqFV66TLOIa9fNHKsH532KC/7/+W3ip/+AbQKwTV9zV
IEvrbuWHcuXoloiSjfdAX0BLmCTcP2tC4cgW4CJA7E9XC1TJKpT4P7sZ1cq2s14j
98GuTLUwnbNfFEKzQh/aVJZ4fUDFppqSsIvb58mtcFihu1g7vG71/nc5+mE1KZK2
UmcvSH6uQ/t8SkCefPTFBOP3jG89C64Lf2/7Po0Dek+MHyLUVaBPbW2AVdB0TC66
kVKaZFPMdDFUp/4dJEcm1FVZMcAgl8O4pAqPwmZBsn/6SoJdZ0eyOkoph4+Jq5W6
qOQyF5d8x29b9tMIqOMsaZR9ckqJnnnXC96g4vUlZQAzSFw0v2IF5QJnyHc62nHb
f+x1dkz37T98S9ZiSgOnxb7mbLUfjQfofCz7xlwHMESE9h10Zv9wymqfwvi0g2pP
rrRJFY6zwS5p26PEEsxZlk2Nlm9AMMgJ5cPLRaf4eP6lSJ3Zg43edsUGFNfJIAqp
PCt/m2ldCSufO6FnvrYZ0Zxj+hPnhVVpLXvXEmufbogmiW2CWctOfzsfpECEJxMv
TRlqSGfpuXWtUaYbAPyH8/HWMsUd8c6z1B8b98rHTB38h6FuZ/qSPwoRZuSF/v6q
foyQTogCBhU83jzHYm/w2fE843m0JywRdnVXgYJsymeEAI335cRdjCs3pF9Nn1DB
tx1UK0MCVepvW0VRENIMV9V4cLg+328oYltnsvhoTxzf4urluJFGNWUT+mqxXfk2
OAblTCsUs2FxN1VsuycsVqmGylZ2vay/FLabnhcL8Ih5Axafcw7nTIh1zAyEyXEt
1uZq2mSVNQcsLm90l35Wp9VKY9P/NvYD4vjV+uqhBYnImU3kTamDF0ocP4Onj1p/
htWFQgorCd3PIhDSnvdCdM+94nTK8SMtOjBJaAQWYc6OOEOSHJt/KvI/9ypmM8Q8
ObWU8xrrK5oyzKKl2E+/SXLZ9OXjPuVmFMsBz7GsGgqmWXHnam4O68VFjEJzMUsa
DVRUGgEcpG/yGrdxPZhUZ4Sv7euVlRa+c6sJdwkjW3W+k5lP2RcWdnfbHXLJgmJU
DuVQY8S1SQU0/UtT2Odu9/WiiULVAX0E3XooFWCUSycqIF233J1e8P8JaN7pgcXA
ZaBkP0mjU9Og+b/5+BcIk4RQvMjtWrf5pVr3/AjHqCeNC5e8pAsxL7cbIvVx1D2d
Ltr57Yygta02c13JmCXsfXkVL0j9GnvkJW1gaY8nUmMm3BzrxWuaJO7BTqmv/s5r
ItDjwehm/aoYIQLSTIvE/Q1J8xpvxNFeIz9VpvmYpavkDc6GQdk+TCAMqVz0ALPg
bTrqPmTBpHoYBGsOWHhH5e4UtliMliY3RDFPlrwpF/hbLZTv4nsz2xw1WPP1JK1x
dXw1u8mFXa0fIGb17n9PNzOce5uigDOtBIL2GxNlW5kYUTICtQothQAICcIN2qiZ
/yeHqA3dwvoP4gbHulWplWQJkCP5RXB3BDFuNeuDp3F4WIliaLTtFdrGjrIP/5dK
XXdhe7a0uhNAC6TXDKqjs5ksepyRUyx1NW77kvWYQBL6riOMFZ3NEbjKaWcBd9LU
QQf+GXEi+ft7MEiY2sTMPNAEMcnwKxjFwTO7piJbo7xhizbZ2xiSQ+0CUaTkp1bx
dXsFS1+gZKcqE9PtYoEnXxA5oCfEHiUbHA2QAiMzd7FnmuLiK5NWSQBbDs6r5jm4
UzonDLo0rwtZsxe3lY5KHCoXArYWCvLRBnmbNTZRg4ArpTQnkN89vEV2UvEyebBO
uWNVY1V+zPL1LIpV0tu2nlYTb11iEodPhvS4LX0oIphZXVRLnF/XFJVuYgDyQLVl
PF50D0RqbzzsUkV+YAalXgIzfKipABwbdeVxHghTl7pW6HEr3wrDavSeCz3O1qP+
u1LKsEIgyXk0o6ud+24IbOv0mOjAOpDXhT/GuyTCrHANKHkxJuneG2FvZoxTzK7u
ZZ/lNB8p1453TTpeBu/HUwwX0I4eKenmt0n1s/Ox5vf02gmtV1GtTpQVxgU/BSIs
7gB3oWet0IWhR38lgfQUh2CVBq+L4JehD76CqSiC0fL7ttlIm/yZDyT4pmbyr6cd
rk/wks5iwGbMVMuKu9KmTtKcCBlXAC/H0NrVvsTUE4GdWGO9GdyoslbkOL5c5xdm
jE0z23rXHFqFQwMDzhi7biGbqFCwc5bmowQL0eRFhVJj5S40hEaxcMJWBedc4eH4
aSJSkXcuqNG0jGnpH6iyUTnX2sMwq4y9bapnDqTYCcVFFGwSAvHCeqg10VkVLCLA
QNq2tUpW40zJuDUaeaySIepfF7IwlQVhQriL/t88PX+KXKt00RKAFKn4dPhsaOZ1
SL+v9u+mcBkQlz0QMR1pTHaa1iR02zRPD7NeGCJO/RvTnO3gHlgArQLJ5UFqEg4U
6kVeVwCmX+ooBx0l5StzcbVUb0o3jL1Xul7D50zL4icxdtLkaRsw17WD3AddlcZ9
pFfmV62qWG8MHNu3/Z/qf/NkaoO5sRSzrTTfvDtoeRSEbE063uDVS6VDljAQTFxC
A+Yo4u61Cwgc+BIS0SIAbtbsL2Bx7X3uUkeUKrPgHvzVX6lphmYe9YgRs22l3kjC
vwkSAsjo6z8hRyUE/12Ve7pqZRcwQNq9I8e3HNRO2Im5aYZsPFf2OlIuUzFIkER+
eqj3sSk+TzNfLN60mJ7gwUMnmAgBOdquzAwOQTPBOohLHdqXM2gH7ZJ87uzYu2qq
gf9tb+/dK1I4cqZmwyR02mAtKkLI/9lkQU1aTxJnaEgcptlJ4oFtA+d9JkeRmnty
W9u+GE96UB3f/snFF5yxF+c1KYLpK58RqPIi99ieu0sSr3NlDAKhHrTOkv6jSAEP
8BsPfeoW0HQ3/aaJ9+F4bNF+21i1fUA08Ns9VMhdDmiMuRNyhjTnwBscV2mApmAY
qPz5To6/TdU7UAIUjwR1xBUQ1aNTcor/139F6Ta/hHtx7OpHQM3YAsKwvPEm2QvQ
3sCjfdkf0F7DJGFWsp6aHzleWEK3+BtNOzwYKpTu/bR3U0TfAVtAVAirmp82m42h
rk3EmaVdiCua4dOnFx/ZYMT914WSwJl0o8zFemazjAS3UML4jki0serZDAhyJhXB
uIWYhsoMmLitx/839WThS9ZNLlXVYYIeooYeOuv6AH2OmMRc35EFdC67phNc0P2n
2NYSW/K5oTm7NTx/PIJ6f995pUcxKYtylAZdl6ctfuzE09EknHdSOAgB2C1CitfN
vNVoW8nTLkZCN/jgqtIKx0aAUE6XvKvObwjlHxAVVb/tS4Zd47bKzeSQou0m/1IK
b9EW9Ux0wsORb6MkxpNVAWOlLeUWAuKc5gBtYlGN9L2AGpPu3dGJDlEf/vWWb1bR
O+z0gYVLaBiuaFwK2GuyrBYPDpXxvYvem6ms9JTSXRYguvOTycC1zbZxZD6p1yEE
4V71w+V0Dd5VmVDattl1f1yvIqJGwIMHdOraNE842dqnd/XzDqxvhbikCwnCODhi
6OgT5PavMxpxEnhpYpohbbEieC1Ylppc/XR0tsZjXegWK9mfL/Fbqz8ZKrZJH0k6
wNxdGVMC5n5Cx5XpHgGnJNmwyPUN5qIHVTXmsO67AdUawEyHhQFWEJCEQNyJzBGY
kzkQbhHNKTGjNu7HRKu/JDHsmcSOzMXc/C8zlCPnQlLkHCBM/tNQpPw3d4iT2KGI
J1ijmEo9dVAQ34Dzw5RQUMCm6kjKfMgorCXLK7KHjOHcdq3GjkKvJHCUjxie/CZM
UBzr90z/Kz1POziD1MgKVIBV9ukwfSGT6HONm9/NLQo/UyIVXxuIHQMPh3ttJfT/
p28pOIjByZGXcsjln+PqMyKC3M//2LXb/XIKdwn3GYnHBIWmg95T171YJcHpcZDD
FcCm/s93KWKOpxX9m3UnsTL/0HAT0mJEAnPFaR2ZAUVSVP+eDCg+f4QYACOyMDFN
E5qAZSpQcldSuNHOMgYYSgjtOQq2I6++fsZSVsZBQIJa7vIMm1RMgNUiJ18aWrUl
1Pct35seuPplI0ZDbAtdTSPiFczlNhawrmcIG+OEElVY4vygSwGb/X0CGmtnPQK6
fsN8eYKUdrZ/ELLThAozj5GqAazDI9+yTbddAUCMCmZ7RoEWd7lrnuV/zo/YcvLQ
qCid2rlbkkYM/uU3L75HAeuQ1m1Z4E1zGBDLUd2/ciGIqR1jTI4wcgSPNcTnX6ap
Iq1CT9TmOvOGyEA5M9MNSeQYdlD9LpXx/oPZJfMnFkvMA+vx3WpQy0juEC3lFVhX
2/cYDw4Kr6QJGc1sBmS66TmaKXAJ6KZLMwV5Qul526jCMog4OqcDBh7hNqy4VCBi
9bd2iJ9A28EIaEe1nILFGxMlo1SgcuzAoE0BLOrRn8V7AZTG+XWCjmbO7VS8a04Y
sOOW6C3/3G/VGRuW1nc8QWXttke9ZJKkaoEdJHD9oYF7msnsCO6tKIEoihAxiBWt
44bdzqFzcyGmC8hvNaqvpgaLMt1a6dWvy8Y9mKbeAA1FL7iw4i8qj2Gm95Nv6a4b
DEhUNDEC3SE7Gd9honzRyLm9RDVWqTkEJQKy/bxWRSjbuOuN4SPMGdwa0OmMurQ/
S7Xn6ATCiBrrtGVfbd4JxEZtk7s2vLQ6tvldxnNw1D429Kd6fwIpJNwzKvG3x+1e
6g7xV4a+NNDQD3HEFpqwgI5dQqEA4VBH2oMMU8SKr4JHrNlf51G5fZ5uelGjJdAg
kjqdLREdsu2L80hXJh2MD/Ej+ONrPQxfTXd3uteUuYoGT0k0VgmZO519tbBZPUZa
LO2VsDZI9jYkI50KHhsOOlpas0OW24vpwgH5/lesIpylsY8LycgB0FI4XNkMRaww
9VTGP2NWYd6Li5dj/9V14fkCd7Ql1xxcG0ckb3ewYP1Kf8EPwi53bUNvCpbyrdLd
W/KJ4pf8ZctlSM1SyJuTq9HmrQknM1CjzsyIkLURAtwxr0ojjWWbAbxqcfHf+aD5
J4WGFaYizNchC8dRWrQMYGx80TswUOxQEgsXUJxs1i6tiyNpHkt/oO5/5SuMLNhE
pIn3uFGxdHv/3viqNIlUo72J/hv2vyzTE8PJArtN3GIqNJnAOHowW13HjtZORH25
y5s1uPujj2k26hvebeZh2FqwL3eneauyAyXh73k5K50Qi0QkH4TpBBfquRK82yh+
2tn/bHd+XD2ZGht3yfsXutWz/x3Zias5SIHtx2h8QcFDA1S8pGEsywltdw3rmfyZ
Pm6fBi8KRkOptdVk3AXjlAnhREqXMlYFh7ceYSYkxJblwWR3JFMNSUITUY/Avw3M
lH8ZDNS3mbnML5y+v7xmXoNjKiYDtSvlBog5nUNpR2UNqGOvseJioQQdQmzjFhs2
o8fi3lJ3R7conWO/RAxjY1tg8ofkic62wHNOb81tEvS8itvwzHjSda/j5n0ivlDd
6soQoSB4el5Ge4CWceET7oZjWkW9kBcPUEqtBh2bVpS793Sa00ZDzpC5OPQx50Ea
1SdkwtqM023SNse1o1hRG8/WwBeZ3s9fApDj9HTMK40nQCMjTv35Bt5U5IAEjsVl
SoZqCL1sItStHpneuIilK8q1aNY14hetaEd35QqeSWl+XfjjKbdMRM+2JvAjYkXY
uYfClAZTUaAdHGgz0a1q0khIrVFH3584otkMFXw96ucStuDJ7t03S0Zd0NjUz2Xs
OCntex+viCa54CHC1xDljyiL/DXxX1d2SlMS9FIehO+FsV1Q5253whBSkOVYpMva
c3m9vzXVytlkY/lX7FSDH/rsnCW4HcL2l/iN0G8qn40mYt5Mhxj9Qrqw/2zO3ejy
WmwReiPuw0BdJURTN7sVBCY6WIeauQS086JY9HI0yal3RKfyRjVzUzi6UueeJjif
NZKuXni0QRXmeoNH43roLhcdTg6N1dAxw4OQOdBRxqvzZ0XT1xlRQlCyTTdlk/4J
iaN/i2Nyn8LrKSR3ZawWBqtw/TMO+DoHDoiBk/MZaM5h3755Q7WSWnRHcYrzsiAp
16DnkKE2uU3x/zl8HfDdFq1LiQ+tTQ/gVOF+CcsBfYySWdcdSFnXDGRKS82O1XtM
fH3TRNtl9w1dbl6j3p6zztTzXFA84V1bmnSX7toedaQYRb+Gue/tp4mcJ6hsGHTL
onKVNaX8ZgvHWjdKCZ9jxv2iNpB5ov5KuCRfCk+hlnz9GiWxf+qivL6DqfXRMOVd
IHyyHAlgGS/yS1Kepd7Ar+4yIxepDmqxgs8HgrmVp3g26E2Kzzgk67mCXrsKxcHD
Udmgtm8xTruJvpDdFlIssFRIfd6GB24VJ/y2zhLaQWu7dIaVrCBP4C28t3sCd+vQ
+PAgzeMCuePVAe0yvvyY3MXWyX04Vx2XqfQnRI3YNtSxSni1fIZuCoEIFHeI/nsk
xXWRvf8myucIZospi2oOrDDB6Ik6Z8wKlEVvVjJsATFSVCrN4UqaxeiIja1v6ZVc
KRbkMSewPbtqZ2jI7OukB34Tn82MNY1L9noNw6DS8H1+v1051ax0tKBRFoT8dKPQ
IKrRcx0bEWdOV2/CgWvdkLdNc6Ha0qU/PGwbKMZP8vpBfcC7RwqcDxX6QwzRGZEe
ySGvLArZir+W5syN0VFA/zP6vaZxTSSgnsUB1d35WDqhkOqwiZuK47EJEtHC2cbf
0Zcgv2/6VVILW9eX+GbZx8vuXAt8qHynYfV6vMn8mIgpkwFsJrnuTBaT78/XDarf
0nkTmOi4xcndnfg1MyPcwGl2KAlGY1slReYiuEyKjENA9VGwA82noxJN0oPK3w+H
xezN2u56yqXgT2XXYTu7iDWZUt0JrTbnnpIN9KPE5Ycw4g2fcytdvhzMgy3xpTNp
6GeSeZNuoKt1iLFnMmvHk0eejGo+FT5Wsnf5ukEXp8v5pVoWamdKY2EsyPo+8lAs
070ZF8gJ33z0W/X1N3T3ebx65qhEVUfWlETLttr5BpH0yMwuhkioBSjof8YVH4gq
cLwS+m27inqi1+JG6bp+694mcWIjGREswBG+vp7R07CXpwrVSLxJ+FB2g9Es4X3l
mQ1k947yFS1aMNO+BGNRV7iNJCaQvmnAixDVM9wOtSO+rOEYTI0xXUh2HLWF4Fqf
swKYKEsD8DnG1A/oE6ORii2AlVFahTDvEGsg3LxZ/DUbZK6VbamQ/9dD+0E++fcR
4RjmsEjJCjp5v4X+CU7RYjP1a+LYtCDdMb9F09ygoaKl+g7Z6FBHNBkqycfGflkF
GXaOwcUQyLtij7DG8f8784rqkPs5ooxmfxc1iovOnirMHxaXdpbJPNZCthb+3KMU
sHoCqUGJDkoyRWFjF9A1ZCMZRxqfocrlLKNBuiEo6diB+N4Akf3SVmm33XhDcELf
Ac74qu+GIGmVqI1FdVeO6I6zdBFQH6dxD8ElyoRB5+zjuEwA0hslnw6a3ISZnlu3
EJF2asjLzLomkV563mevqw7dYpeO+bBsODAJ/T3z4XcURKcJd8Ur0IOmYU313fp3
BFudp/jn1j4XaOr5dr5jbuFNn4oV+rim5ptC7jkI3monqCpX9sJSvRQvH+i9UR4x
ABO6NDqPljL73fMSqYvZSNFteSTV5bnprQEt2CpE4r2qZqFh5a4NPdVx9d1CreNg
iW3089fpFbG0CwMbl79EJ6TAzintTVDKGfH9BAwEIVl30PJuQd9twbJQpVlxZXwL
hm1u4xkxD6c1NwVcIltjeuOX2FW0ZAObJw+VoiXhaW5pYpY8kZLNKxmCu86v+7si
r93duU0CZ4B/kmlr6hNiVc5YXXqg3lhzrAorJvrb+u/Sqdy48n3xMNBFyC8mbLTC
Gkf1XkKFpAJRWxLta/tC2CsjgaObJfdTGnWcC+xBU2yos+O7bKeIBTflKg/q4M6n
ZV0WTDmL4KiYh3Cmq991NiXJ7qCzF54wP1H7G8iADtql5zuetHjAZjNNTRrw3TfX
ud75p938MSDbb5Q6ccNBd39Sj4Vl97Azd7tyg0zHr1S67CA7rPgxs612ErOPHvcW
g3qbhF0xsU6ACFLKhcNYbLDcF5DGE1NaAoRVXMgIFFkY3Y3U5AnCk9fykuqii2yN
rKzr+aNPRNsxvbwkG/3C+54PD+TU7AVJZpDwLGyeA/ufgGiER26s3X+NdeTLz5OM
dlQwrAIfngIXexRbS9bj8DjFVhjQNhqZPFzrRjSwYHEiF9NIYfAxgqkD2GSbPDAE
NmlUs6dVNYvQf2leJ3ujzdlDQHDg0OQmvUR/DUOR5UqTZt42RcJiaRw4gsn12Hu1
5y8NQAhpll7omJiWn9O2a+mAbpOSZkrEhI42OC2WnuspVWbBxBKHbhBbwMlAL/aN
/kVpDIEyad9g5vsZhHRMkp9dSSZBYmK8Y3KPbjA5RBNgdwC112xQZtUkgoBw4Oi7
l8d3dD7cQWWhuARreU1hqby7d82B7j82RB27+X4sa2+PeLXGpOQUrTEnb/i5MZVu
zOpreL9uJkUE7rPUxRRHxIfjeJ/zcmyFNhaFZkl3P1ej594RrPUMghMP7k/9zrAk
Nw1kRiNlqo8o9m06cJ+ueJlpzM+3f8SRVhqxG9AM1jCO7vUzcH5XXg8HirMQrpzN
ySQdq41A/s6dETQAO6GwZnYnxaDZuxoiSHjxPxLMf5X/hEQDLOTcmD7aA65SuL4R
LC6jQwsKmcSgG2T0hR+oPEdUsKkt/5DI+tgPxmAD0rwQBI0axomx4l8SNkgi5612
CHAFO6eOQLLAyLzOX6xjac2L0blXnXXvOqsxN0BkYKwlBKR7SVIayem7G/35zzFv
04PY7tCEtQlWpIj+89zSiNCyBgAEqDsnoK7ZZaQFurJ1DMOHo4CfCVeDHrnVtw1h
OXtMEr8vJTroRkWdaZq6ufw6LpI3Fk0DMstxB+g3O5105inoHQvJrjvDPqMFbfpz
aqq7ISsh4UL8ksj43qPtzA8xO7/qYMkOXAoZKYF0HlBgbip1vcSjaYKcI/HG84VC
TIWcnVq5IGHTPuY6de22Uiv8njsX5OpH2APgplSrsxn9dVKtxbXfq6QmQDHq7mxF
q2CMF2AkWkz5QJuA1XXVIBzjloyfk/iUSvkz36HJ1Vn4Zfb80iFYbWQUPswghAA2
iRaTZer70hPIkG3M/EWmCkjJPRZBwjS9LUxM50ZrIWRU4209TjmKl609/h0fKxUV
Twx6FjKt09ZHLSWXcevdwmHQWC34LBeaQDOqacSP8UERjuANUaOv15KxpNm2NSmf
ThvB4aqUx8H8G49aXfYzHa69fcVr7XUmNoBFH+ZT2J9oiTuLVX1meQkte4Z1jpTN
eZkj1n7MWfMBi4nc51q3uZrZG7b6/Ef8LmxijV+s2Ni/fLPHAg06msoGgU16nDnI
RkdQHErdqtsw7UkXd8UQUGUeXvJYQk3M7rarZAYaierzzXOX+kKk8lLgpcf9Hl7b
0gg5kl8v2/dEhfXyOtm38S+8woz3akKbponIadil+flmKdAUqrnx3SjhdmhtXjY2
VGex9UrMZywPpn3iBZOjhGYwZUNu9VY2wPO0MaMwu8TvfZwvUe5Pnmf3oz2m8T/x
esPg6c/tEWmJRbPGwKHhuPySOsHWyZYSBlUcydldXkHHAmJ4q2L4c1HtKEj0fOR5
bOgCA/fXqPZX2jCAFmPy4SkVBglfSZHUHQKsaV6X3kkBPrznBEqiuqAbsTqoX7sV
tdxK6XY8lEC1Vh/ALdeqvAlC+7E4fVPRjk+wv1a0nRIVGqxwm0Q88+hq+QA6Jdlv
vcGLR1FELFoVjv1QBhrWcgU6GsCD3ZsPAEbuwJORJtPIgzw+Lti11gjsvZczd8D9
GgdMl2GOIYe1aNcu1E4crGbRn6xNSAU/ARCKffq8wpOX9+IkDE9Xc96JkGHqHqP8
o0skkvK3QqBkkbNEG+zxbNss6uCzYboob297XjVPBGzgRr/E3v0SYeTvb23EYedH
q+USw5RqVseek+Wtc7t4+JAqphdferjIMzOWelx33+SA7CZ05Q/4ispFFRzhBjHB
HpH92/awpY8uQorD65+A4++6vQURxXOHo8oC3/dTj/ze3qnFuBj697MUQX+WQ39C
QqFrSSryHB1OYXcTAabF9AD+gLDH7uBeiM9pY9lREuk4r5D1tmNOjsvwuolpjapy
QjqwGhtuWZFF+jKk5V404lqGvJE1NLSIL5WD20IRkwTkGH1bDpvCrTlyr3jav2Ze
fSZup0ElXAx/90MQ+JZol8vQ2RZG9FOEjvqlSQrNC1tbvpKjEctSPW8o2gNZXZJn
RBjIdHSRITgBnO9FIqJ1deyGcl2jSR6Dea0goOAFmFEwM03EzYpVL8lGbW1EkYSp
cy2CJBMonUFWH1Qt8qra3xAYglzX18f7stpJXQmUV7pig73/KaSS8MyB+K7hh+Fz
VKEp9U+jaeTL9v0EOQ3x5+JEl23seJ20NTjcW1ukYsjBW7vnEJTwAN0/jfecKeR2
39NnQiNTcVM+NlfMrCsFyRMVRJgGOTYBLjPRpZU9CD7DN1NyP9lDRalxHWFhEXfD
5yB8vkihmbkWr2ybZOImYKoVC7bJvCXiQoCG9Lgt6rPX/as8Nf58USjLJoQdxNAg
OqC2VVnnM34TCiinPDMK//TB81ZJMFuRqQZzVk10uZxjh9ya0jbc5D/ERsD/ht5v
c0QGF+mzqIqXa3Je0cSXVm7oo2G5PTpEmpx+n7OiqnjHA8mZ+cB75WG7F3uPCiQM
olTCJv4vdpoqdCURfwl9n9twqWDC8d15/VS3xNNi7hZJyV2+koD7ZfJ8gaqleFIh
6rPjNnPVhcelm68BKXlMEYkdjrTClCbwJ4wd/Vq5xLGy8tVJNgteZVCBOn6byeey
YXqmNZ4eSwwBsGyyvRorjnl+R94ofvEw4yKdrg03PnIpW4s8sF57/PzUY/t1AaNW
lkfuqAY3g68dduS+tgAGJLeiDJyRUJh/Like05ZmqVnUGmak1nfZt74mvTF0Mypz
HerWsdJ4BiHMnlNKkmIrS+ls7igZvbglEOpIZYDj+b8NiVOsElB+Y2xlQTfipLpn
QAdPwxky2TfNIrnJ4f1d8M9FD2tCqXOPFuH8dzb72TvNvrIXoH9Juh7R7ms1cHuR
1tQ44GFsK/dm/Ws3dGOf7Wpzlseti+4DQ4iDOdPG/at/o83cdSXfeYzJyJE+L5je
oCjwSzs630x/ZSTwiBJBZ+iBWrNF5AnqCqvBmExyRaHOaSazHVgLlMvBY0QNipXn
dzkdVyp7DxMzUQxThR82n/jYerWf6ljqEUuFfLes6QACEqVXgOWIcOKMZwoEXpcd
8zUQiuPFSTiPm7JXgc1duNNCKCWd+ci/nM34x0NBc8TFBFKpRLDtkU2t3LcyyI7B
8o4KFaAhiSODmFKDz6lpcx3iug5zU6ZORzkdDtzui2IMCm9XsIgHlsFqv1VzmijY
qJGtszp/d2CN5Osr9oDGAGXo0a+SRuyQHBejhlMlyoNpRFB14ToQ+RN8UaWeeb34
wIjLJlVeubr3QL/unDtCaaW7HQBsjr+m0la0k4u3snE4BYwrley432kqud4g3eds
KGvEwbwMvFEUpM202ARA76/myJnETVewJTTushPPxDMv1jwJtGK4OhMRS4nX8z7k
cn2TgGLsKWnGcZkRxcN/PmQCpPZQOFsrRSI9BICfa1vH68gE+riWWmZG05Qy4U8G
7JAyCtGwvHVBJQD2zwNke5Yuel3wRenQDEqLDDBVxbKLWPlgKSEpxGKggZQiBIN6
wkVBtAe5YWiSmNJ0kMr4Ku2DBsLX610XSlnlDd3RUj9p1y0vV9if4u0tFeO8Eqgt
HoesoM6XyFa2SnaDyYoAK6GZbVkXPEdqhkLmQlnA0TWOqvkmFiYxOnvzJMpMNZJn
4sQXICsVTMO2pjV6pwFLZO5T8b+XV0jQwlSlxeAXjEoNeKdhonmT/yIyLsjFfPxk
nMwe8pWnVS07VQp6G5IdCUSq8bTl0oSn7pLwmvrVDr+jaO8gcz5XzwNKo/8jzPU3
wKRJ4ts4VnMj4LL1SDakbYcE2uCnXGAwBzZurelTrUBHDjCyiCELcSo5Kg1jCm6e
Pp5YZdJLR0fKtkwJMgEdJQVkR5RyNUXwi0wn5/L6mJs+aHMABFig1KXUzmbOZlg7
VrcJZyTWoZ+9UW8xwh+G7I6i8ZdEo7xOktAFT5AMm9di0nx3RVhgu/O5vtqcO9VB
CIRTOLuF9X4gwMhfmFYxnpUF+IERmsei2r4pAMrLblH/6JgQ9D4vka92Bvzvv1ed
KMKc3Jpk7j+MtW0HW6xQm/9sLPycwfAW3RRFh2uHFlqg1l8i2vsOm2FfdscEyU0X
pUE4XffEWWgzkkPDHPxtOMXfZdqIQmMxwplMdZNHTvO1zLih+v9YLjXmHpmm+gv1
nq/nv0Q8abOVBQQC4zbJ4pQ39x7c7/iqIo0MfkWIGVATRADxdrjwT5ZfO8XyPSar
+sxUppQJh7oPLwu3BnfMaBb/4do8x3SnPm/fB07bGP7if+/00Z6TYLPYB9d4ZSir
xEU9FBOrLfioXZG+TLBxtlut5CR4Ns2AE4MhBTVpchpCNf02sYKXHRtPX6rQoMxw
XoWPwadfgPJ12PxX5s+d3FkCS0wJxJvLIx7S5CGsfamXlX1SFb8SGSREBv1/d2Hh
hWpTRYpW3agU5U36gmviM4iSDwAbhvZFO9m+klNqWwvPhIjo7gXepBb/7cJmMIKD
EWUXbnznGI46a5e2fa0Ey+++GY4UGe2NWLdEJ9zgFvk3k/NYpY7OJZUvbyuenTs1
IfST41nY0ruMkW2F6BUlQT/iwccjem6lUc0EDm/XX+AmLxl7aaZHV4B4dH1cHcGS
TB8ne+6CnEDIOa7JN48nPAyiC7+0CzEoryjksrPJtIo5CxFN2oOs1AY+6TDcxXKq
UDjlsA1iSxK6ZjjqED2hQkdqqMo5ZLm/NmoIagIb5MKMHWo/rjThm2qvz0JLxxl8
JM/JF1aIRYFUot+CyWjyaYMDcOWpEzlqoOxcR2QiK4v2mjAlmBFHGLHYm4Uvz4SU
YCDaTB0hkL7VCpNRqZ5uWpHimq2OqBj12S8gpvToskixzEuFy3R9471QhDffoK7F
rebOmZ6YOMV/05/njeC7siJcoQ8ziEFvTSEgvfs9GqnUo37/st0WX3WzbvhtUJB1
vGHqNYZM1R9d664D4flLAQONNBfUw7iSTvk3E2Oc87pI7G/kp96lqEVmXm4NMDQb
r6KfUmyeZRTOf8B2kbRmkn/qEsG934GZnug0jRB+wFMM6sL29YAOquU+iO2Nef0o
n4/ERip+mMO2qzmujcPShcU0swREqINKS2KGh4NGLuVZFs6swooQQS2Ym5FSsVgb
NJvPtpVMNUHIrCop0qctAfzzKYLtFOOEpWVCGv5nOyu27j759K6jMdM++Oo6Wmgx
P8ntvFsrU5H3m3n0JXHG5giPstDd8EUYJpyZodrGk6z+EJdVYTKgm0lzKl8lHTQl
MXatP4QkOhNtAik6F9QcJ/8FeZ2EzJ73Z+AT+9qGdZIy0lZhP3/efSj5YzSbjoy0
n2YxWqz+lj/vcdsfqzj5cSI3oTHP+U4F2joZ/zxQ0Y3hZMYvv5B+GNMUgTXHKXbm
WEY5k0IJouN4asadPhbfqaSy0Fhp9YWEZVIUTL1/H2tb59r2P6pVzX7C/wbgu43r
YHt+qqfV52y6JXpqIr/VK6ifaOh7+8BE0J99r1rk2yb4gxFyzrzDYJ3pJRpR43l8
HBhfr8ISlLU2s1385mQQsoWlZprSDE5u8o6BNHNGOzC2qTHHVXKKunjxZaLIp2Gr
XTnO8NWUUiKGATTQ18avBArKhX2H0rPuzfveTxbL4nV4CAFCv4imHoPlmkMlUrsM
UMYsin45sl5yZ8tXXGuYMP0jSz8z6bPzpfB+QX7eCZ8fLqYvksL7Mmdz1+qyxfRw
oKnGA5AO70fbf3WLcktjzHjiowsJXN1vSw2U6hjKmdpFJ0l1l2nyux5Y9GnYFAZ1
HD2ZdWQIQ/pujHUkdz5RFJ4XARPBysDDBtN5+qamhkNqlobzVuMA4jcwvIca8SwN
EgpxQrg45KiBCXBShECMaA7LDDxGWmNn4CjRWPItT89E+CHTdnZgmCvY1D8O6Mp9
W+/oYJhj+ldW0eA8P5pVkEZfhX9Pxs1npVDlU0R0j4OZhrijdWAghGKEI+SChFkl
TWWbbZ0mk0pAo4p3dPvEWRWHXc7a9t7Y9NZgkmQ93Y53saqIeC3iLdcX93A2WM80
VoVObyhMaD19veQiqXUfdC5aVQzzkveefqzwWsJFMUM4g/7qCd+hTz/PkYbWiXjS
OLI0rS8MVbgHF6BHUEW07/vVIn8caFjWTuO4jgehuCaw6mU2p1tWKI0ilKynr+Cl
6d97IokE70HwK92sFXywo6x2QdtL43vB4t1Wknwid90zMMsY3hyD9kzdMvDqTyl1
ZW3pmnBrmJGUmLua6aym2jwIdG1jJvONMx5lwa1w7rt9+NbsDPoNoP3U9m9f9EUt
PyKzX384DxbEOW6cjSh1CF8tK787xLXDg82tPeVHCkPO3W8yVHSH+/4U0bZGHELj
48dZUhGufKcZoMOylo5PHXvAyIh7fQgMfYNHvnzDGs/rC9A7VKorzq9W8e4x2DdI
FJ+G07/tPX9ACdWrM5ICYCocipGQUVuL8Gs1jQz2ak7Xkvjrg+PT+N5addI2HvfF
GTlP8fV0OD84MTXEBHFc5mAn15SvVd0MiG+ZwqOryyxK3IwIhzZ3SAFBmD4f0Yo9
7BQydWbfdLnPuEbUU43IjJmO49tJRegiKEXSEcHsLUkQImdcC79SPFTYMeOakkGc
T2lHv3ldkR7qbm/p3cFFA3680oI73NSEu7vxwGG0f0v0Dz2uWsSW54A7ZlIBuWb+
PD8CW+RpcMuy2Ks5qM3BzguoW2MKyOrQ3xBj/SQx2ArvBk4zye1bZCfEfvbfy+RP
GpSXbh16WWwTN3QAk9jnUKuyWFaXDQZPI/r2qrtzSmqz/2kwvI2TI30OSoydMO/x
QO3SUMXmGPGGV+q7g74iaviDYeoBvi58wYQ1AWqPA7mbZmjJGWjD7HvqFHciI0QI
rRaqEOUxLEikxKyNLlLvwW9rL0/vslF/x+hV7zJ6e743/GiL330mwuOtZxtoD4qr
mH51pbnN643qdWnZtlvy7ThWAo3X+xAvxC8UtXHuyCtJm2s2Yp5e0AdGeObwJvOb
Qh8C3ExfUpUrH9TnxENBmraYS4xwY4qa27R2KnN0gVYlO8vQyHxtNXpuKZrzPWJb
F84eq0FmKWrgL0CgTbN7Q7rXfWaqqSZks5fG4ue7tB9jTTGSKTsUyzrKwQsd0eM6
b8gQMWFyxRscC4tkXQTHP8reTHkAMl6X3+lRzZ6hLbLDRg8W8Hw1tRetxczMCZmO
wrby8MXcVqgnbi86exCbcludEl9xeIotsUKg15IQ9f6zGrwsjLMo310Ssj+zcy2J
kvivlYMSvKp6c1srIcyHmuqYqcQLKy8G1nk/CMRT1fyQ6oC9qUWLk8pzdmrtdsdX
WOPjmSCZGs1EH9Eyknrl/237WT/p+I+j9clcFkTJ6bEi2Un7SbehGs0ysyFesiGq
zMWhsliHHDKdbq3x+kt45QfoPa4R+9XUCCHYJT3juYISFXswBXJOx3Iy96qHSCwF
4THra3OVAXH5/7tgFNTelYxV2WmIo7dl1SnvFNyZcyAroCSy7M8ky/hcl/hl/thv
Ue5pFqpOrXEaH9D7VNqIblg+aSoB4BW6K2txm0DzSRvpq+i7hAO73d9b/zfEqYj/
zXyLBP8nVF5WX4s2g5rTqDVh64UtvJSzUL1jZDwinkWyYZgk8CIkZht/c5pgWb+b
k4YVA9sMzvVpfCICHlSjX0KptxhOXngL+J8bfVwlKekvf6/KMLpN92BumJNPK9VO
BH9vvxwG/nFIX3QJbjlUxlMUNpoZcna9DgRqaNcLZaTRFkGMjOpfY/ngGUKjGyhG
q50Aidri8EYK4snh4POWGbZ0hWy0LAJPgzUvZRsGKdzxXuyy9ihQh0tln6/jymo0
5I93Sm8g+Ok7t+z24Nx+QWEwVqU3BiZ9gihIuzmeF/76xLEtN5ANfjRh5ZbDxMEW
aJbgOI/+xXf1Bn+aKfj29ZmS0nqiAUAKmEvtYDGBJNBeasNvFlV2/uEAdT/LnHGG
aMt1Nf7iW54bvjkh0juC36wmeCGKx/6XSxfr7PGtjrTNIAVpQkRuW3tdRkEZhEQk
mXJLzdxPNDqCBDGaTIXKzrTAGCTvE5cUD88j39qL9Ojz+DG/LngE3HAq9APHANz/
No8GnnT/yz4hot8Lmx9V/UBQIA7k7Nfmtc4+34FvD6rficpPDMzHLfx+7kcq+z91
XnIPsFXDU8LEqnN5Mbn+bGukHUdRJ2vmgjz3o8tqY73fy6UtJRTWCEEa+6G79hmj
IF8OD5EOYM5i5+22qmluv1avuky1VYwRZ5lamPSoZWpLvr2xjNeSfEy2DjJFkfk2
T/46vxCePE0Npe65A4m1Ea3Mck4eQUDFS3N1T378STkTZnS3TQKH8WtKOcTNEFTa
TIotY13POJuM8CJMhoMEgySg3e0a7c/ZukD/n1gHrCohYcCMnnYu1HGOsnDhq/Hw
9R5/gcYmcAjqL7Kc8/8PeVrdrequ01bVlwXUzWwoITPkov4GhpI4B3aXdLzqr22l
3xWaVFKlYikTn1eXbTZBnkrlvKyiGv4f+R7XdMPLnFs7DqgOK54vdhfhnr2WA69V
x9tIXTMqd6PdEC+W3GpH3RZ1+xq8wGZibtLxish25C8eb2v3HK0xgPM5LW0J67m+
+rbXYmX3E78wK+C22VfPIoMH1KhZWdBHie/vIsEbNH92gq5AtMBfCkV6QuuMv9Z5
jPn49M/CvgC9P8sZe/ywmEZGIduC6KC+nkSnVdcooYw1b4yCzRugbXUezpTyCOgo
t05ZACZNdVW+yOJR/Gz9D1EgfDTkgYYelPCiVh1KJy2xU6QGRRZXARPiqTN1sKDi
xOm8l3rnsvxz65fdWShu8nVqahS+0FyT/0D9o/DBv67mE/BqLfpkGm6iUvTyp9it
7FuxTWxMAOeFvFogJbIZ+c7yTjON+PUiuVY29xEPsPvPXrcjyHNP5Pn/d4KmPkdx
+oMMXw3sY7xLZ/oC1qOPC8JX8TQltp/62Vmwr+k3BE8Rt4qv2xxX0ym1fxKQXKPe
d2jv2LIL2jQaZOTVFsqVHyNwjW6UDn17Lb0b2Rz8ZvS4nLSEIejcGUxI8E3ssFrA
OQVryFOHmjFdq9huiMAKHDJNcHVAUWToA52oyng+80HHFv8NqRtILmzBaC3UR/3r
MufjkMfc05zqOBB5ldXRiJTJUjmWo2eY4xi/R86lLS+QAsRQuc668QnFh3TMI+eY
8//PzezFjXFRVPuc8Xs2v6kBXucpaSlvJXJ2/pR5371/Fi56+O9FcF8B4tynGKrB
iQ3rvDcTXzgvbtLOzXZhcwaYfpMXyqm/lzHsY++lnVLBTH+jGyY9E+0a4uhqVyds
A2QdOQBz4skOYCRbqsazKjol3V/HJdo6bEugSCP9OlQ9q4EscjPHmgJRySfA8g7q
p2LcyEBjLyQ70t4ck3kwwUjrrEmX72eHwak2/LASAwB317/KREKshr9r3EwKdvcJ
eQE72feqx3UaU77mFuLdfkXM0BIAFRQaf8sfHJg6ntWj8moQgzhNhBaZfAYgQDfd
u2uiHvSbaRFR+PAK9cyxYAHNEFw36E3ng7RH39VcaTK/bBxGGPuWPYlFllRPUngA
ndQXk6CzF0T6tuZJjaliA65gudqNP8ziL/PR6L5fzHL08hWmRsFabDFoFI7q72yE
NQYYtY5Z9j9gSBuAnyJKeRw6Kg6+kxf1/nsNilwxGxDVgNQiTIYHKBk5sTH1Lit3
1/TQILST5t8ZffwzwNtYwHztfRPoABL8V7TZAT7fcIogZ0ZfX1uwdemLuIngtUXl
60pG8Yf9dmRPlqa836o5h5TOkDcR2ys3Vi17/Ps7ihYjjeiReGaaWRSNJUY+ahoe
Ao0TDMw6Gxq1oThpxodWuVT7xKEYek1Xknc+pwRJctAThIh95jZ9BA7KkRHii5JN
0Ah0xgp3ahcvx4v6/RppO2Ak5ZZsjy1O/SUdbCduMI3ibj/D/915Mww+zPjJU10n
a5JC+6TOsMmtuCUwZ4q1sOBhgdpZJcWtJ+3CQ5WypBoKM3JqwOGfzQtaYHb4EzqR
MqHyKTmOHXbY2rQqs9nTLeuOSEezmVlAeHhPYfQ/m1HkiULSgcDZy4JjipO0LvXK
mHxmW3M4HaFMgeubmVoCq3g5gnzER8GOQjmR9bdUgPGL5VRYkTMBuCKnIfTMthmL
9GfaN5Vl5Z/KxnAykslRlpf49Mti9tvlGzBG1CzGEovsKi2vzq+Tb5qQaF9s86aT
Eh02KY/RaMexENgVtBxfQfgIghaUNFWWrd22tCOmqJ9t78D4aEhugvZ+DM2FOkEf
dl5f9zUJQkPxhiqEClE66akTbWcNS9bSkHNt5ZJh0wehZN9x1y4332lXtgCEJwxx
APHx9NhD57pgawBYCJlfzvQKMVXHuRUXTq4TpA2cLw2nxiITjES8LswexH8y6CXf
6tWF0JTKy9HYmINVqUMbd2SFE735OdfKeOSYvMW92ofvxUTJhkMgyHemUgXXwX8i
plkqPnfwbpIzpZo1M8ag5LqSga/0kCMi7EJJfM4tB4OuqxqA9kYz+BFhB11vVcrO
xMUKqK1+vIGh5j0x4QSmwUCk649Vfv3xlhlEbECq7CtEtSWvo/zL8DoCYTDTNaTg
MkKqaS1zHBiTwEzAugqVZ6lI52eBdDzDCPSRi013BlLAXU2VII5y6V5GS8XprWcu
bFCaTzm/Fg30ZxQ27SuyIOSZdN0sstdkzZVHRt3Zqe4AaKSiMtiMEsRQf1esYtE4
QZ4Wo1QVumH91tKsps8N1wcxA3XxJ1xHYXe2v6PKB+dsSZpp9KCWOzEwJdsERW0Y
ts6ZcrSN5cCFRw5qCjEfobouBr0CIhGnhd6dq8h0DZ4rEcmazq9X1BNY4JCxoPqk
0zMISQpeyRJ2Z/d/zxzXzMV6iN87L0WBrrVtlZgxYrkoW0O9coxHAuyEGXkh6fqS
ne8u3fOpXvgQ4Fye5SgDMTwJzpOff7OuLdFwmA9sW/GiEjDEE3myOH4sgp9sOejZ
U6MCAT+EvHGeNT0YfpGiYXHIywsrgG9YV+9lOc4yuZbxgDQPHKi/OjmI/aRJirbO
/Tm2roNu2oYzs8ELCjjah3IJkJCEZxQAcKlvTQetNRE7ZhvceMZSd2ITcT94+Mjx
rruys5GeHfAwwH70AMYGyZDEUdYqEo/xV3tUHRKWbxYZA1eYxr5T+d0IKnqpS0Oq
0D8NNhus6SUMcpQs854YDzmhO2hzcfPGQAaCBirjQqw5iZc0tqCbiA9zaSQPszQ2
y0a5/ZGwTduGw4OvapYbz3+VSk1Lak6CUPG5b4cWfi3wBYJDpCYDkthkrsAKZXIv
pm3foyUi0aDvq3sidDaFiw4IA8rZ1++flMdDosnXqfhYG0jtsX8dDBcOmILJnA1R
9eg0GJY90Ck8z95zs9oFlCAWzrUpQnywEB3qIirsK7lAYNyTWbhMg5XdrmY2l4h7
3rnIcZPOn2qV5DS9WApG0cFYa8wpeVC4cAChIrWLa8L+6dz8BYHYVHnHKmaq4ypz
t6W8xwSpjUITM0bzWzn+jSaPpeR07XJBAd7FfBs8tmlWxu15Jmnjso/oM9M+Q7FC
XFQYGOlCglPxk8Tp7uP0ME0rdm52VLrzOPUEd7kVF2QNCk3KivIndndtryK4f9HG
kye/oPjqRqCc1GPrKe9BzAP5pz75L9kXfT5gW3rVUGZtqbcMVqzlSeW8MrxFIPEx
RJxtUApbS+EsodnZU6bamS2usmIfFJ8ahLiR3Ih5ig7dhNHM8PRLL7N6koSxV+pq
JgR4KhzI0uWnNcBaiW7LPAeoxPgFh8UHw70zpIUR6tvC4XyaVrk9ZN+16jgBIA+2
NKzE8xtz1hu3KTZeaUBsuRATKKRj7Dgz4NwfT3m8QC/Dv+7P9+MJbrUQy3sag9EP
ntvaU83VVYVylXPuCmdZmt06unIrSZY9rd9jvGzQ+s4sdeIgcBimx7ayLWqq8PNu
NOJ8ZVGGzUv/jJuiCcLelq9488gjbBz5Ff4AQ3AcIWb9zWmQFrsD75etGEWjxo3C
Q/mV4+Qd/cgpIVtpuWWDiWbBxGhhHT2qQexuUNTqhRUnbJJ3Qlb3ZJNgmfWkMv6q
nfglzKZoBOF5tPAPWkFCJGSUdMQEMn6pxlf6Thdv64HCKDnw0EcnAxjfztFTzjKI
9CVfKXeajfhVjr2Xu7Pu4Hi95NIjHjYVwUCXMyY8lXNFoyXxO1j5Dnid44+dvLgM
57APLSel9wDaIS2cp60cEnVMNxCrwyF5DU84ASI6BFBPaeHWt3o6LIw7XVg536JU
hSjmHITzttPFHoLrWHA9kiBIaQEEgMWq8Uoejs0VszvMMQB/V1LR0i92d2jAwfMa
Aja+5qjFYWIalXstdT9XjYJxpaPdjrTXyc/BZCOtVoJuq6i1ROkUNQ3LKd81BkEG
gMS3F3v+AVgAequ9dbbznYtZ+y7kr4AA5SlIQerCwohDCeNyKxs/ypJDfDPl/biC
DA2yjuxqeO1OrIHiYC2KqD2BOr+CfIhhwKRyppYvAZnSXtQb2uIl7kq7Cb9EF7PA
SqITptBTxndtsnI0emFAejpzt6iNd52nBPxtiIAvSJ0RjfXB7MaV0Dmc5y8kS+rW
qRftTkw5J42Bp6y+Qw4cLZABNH4HcXpWC0K6qemQodMq8uB/MsmvzBYCZTg3NTDx
lhFuf0Z2bOto33o5XVl/Uy5ubMjWMq//5jpktS0ib2klv8LuF8kDNR/WY5m4WM2c
ZfuhMVFlfE4bUvXiS4bLEkuTKO1ydiMfi/Vt/kgexV4qvwKwYMVVj7DfiLy/SYzl
xoPVq1ABHtjmux+L96FM7NuI9RumzBdL19m4lhge938Z2LEZcgdZfqpq1MljeiHH
+BIDDx1gH3R391Aq/npcuVPUcjA6JkIxXMfocvf1CO6dPi+rT9UdHpZtNrPe7+IT
MXygeLxTpIkNm/c0QfRyXrTrypuA2mZ+Ok6b4NW0U51ENkcxUxPhvyj9eShykoHw
ouuyVK3lMoGVG/HojghVToyovRh1Zr981bvhlZnd7Aq3TDJ+c88GW1BOoi3YyGaW
qRYE7+Whz3AhmlPN1BVm2yoVmxzaT9sgXBb/a/yuCLrl2cmS3TX25ohZ1RGxuISG
3Sw5CKoA4Nhff0/PrUl3ySSWPWDSOtKvzCbjEsLvPyRnmLRJ3UGIbAOnbx3LEt0G
tty+SwoSudHPeCaZVtea1YvPE+YN7qh9BqEdYpkpI/wZmFIFABVjUqCGcqWA9b5g
3KDr1WlqNiU/HzvFjeqQyntBylUe3RiFwwmN9QGhzh734tL1svDq2VOO2DADT/gT
dk9qqHpmWwg+ikIaCkRuRB1O4Ji1fXVFDLSbKOlSzyTDcOGjOJ4dicKI57M0l20+
oNGI6m4MqRUoreTfAZ55FbMLFaFL96q5o9zP0LMREwzGWAK6sxzeoGPaonrf8j7R
j2BdzbWJfUi+20JfPxS/9b6D/6UebQblC5PVuv5oCPyVuViNsECDP97uNRoHFTEa
14aNMHAUZbJuJ5HgCMPb7WOxxuQgr2BQXFRdC0awTZtDUSbbrobF7oW8hJAgEF8J
M7E863zxVskkaoDDZ0Sy4iqJ3szRtORmsvYcPXNawztG6UlFXIYwIyUXCSCi8nbV
6rdvvvD9upFv99lzOCJlk9Nuxt9TFWr0IX/ohcxNj5fFgWQItExjByUWEPavtN5f
WwmR80qAwneUUOMxxG0GgXvi9j3KVUHiitZq1KryN1PrxVd7SCWogxojTQa6eRDk
EaTI/FFqvg/Zf7MQkhL0pVChWaW2YK4/f6+A7WxuMaYX4LseUNwhuSu/zn4pXBDH
rH03Vj7tQBRnsoHu5oKSPhoiaAVkKpxQ2fy2KDL3T+tHm6g+nuoc081uUiv6gvMc
2qyJb8U4GFFvZBFELnWZ+hF+rBPbBrragCArMMqteoJG4W4mIcDQ3BTmrRTjGvLN
jKGeiNq7bSH/e4+fEU+JRuiobrA/SqZKlPsVFsDrfpiYvUjL+mdYdf+ekR48swer
HI2F2RzDv4PYIIDcoYTSoRxyhDX1m1kl0bKnPgJd1/+KiLNIkxrlQrIMs/1kRswG
+aQr3Ur1Z0EPsF4CFJecyng1D1VQW62DOgN8nnM8y3z5f5s2wP9vs1qu4Fmj4tZc
geDi1GAPNaPHc98xjefxEpEuJCL/PKiO0hrwxh5x+zYgVj28DXA4POTFsQt6tPXE
0D/dwBPw9fg+BKjGN4B9EeKhgX1L213s7nWeG1nu4Bmy622PO44E3ibd0PNZgfqT
T5PVwUNBO30SgtrOfv7GVVTOnagrskCMo/67e3KhnXguaIEsCUCXeprsgcvNpEJi
LTHSblwUZWqqQjP4Xuy6DPHJTbyboHvU3UbTplXPuJZ76EeLrgJyNAPQRLQMR4ef
+DGnXEr4ZoS8ZlY6z+K1FMeQ7Cf9BqVCoWKky5GymfN86Y+qPePTZLL1QeujvzNZ
4pj9ZaIulCPo/pXPKTFxpoy5dvU4TzDG0vqsqLnXbitkZ9uf6y29JwXJPb5kV8Br
hDaAqInoo5AaOhG3qtnnavM4MT+T1YknXp2FCDsAyDcQ2D7kY0rMku9QKxJJYfKA
TNOO1lK9PTYXtt5mlMxbNViiqJgkpFMdJc2e4Md9i/L/lnbe7znO/E45tHzBj1PZ
1/dO8tGQWdRIXhR9c9zr1IQPsPW8p2qx7tD+WVxYLDCkO/JjzBIMm+3TK1slC1lF
SOFosOEI8ywQ40ax9+Hn+IGXuf+Lqsv0+/Dmr8QgK80rP8l+bSlT9ALdd/ZZ+Vw1
Jp7l9YJorxkz1Ig/j5f52c+57YRCfUAXr3KVVNH5HZ94B0y48YIg3ONWuw2mR3kT
xIGyfRWpgfNPlp9ktiFfMF94FvW1zV35m8Us7VAGRu9m8CIVEDGmB2K641wqGOwo
8g+HJVQPEkhyhyr7nRALiLXLSMYJGu2MyFAhLc4OqeRAfCgl7Un3/MoyETI+Ydjz
Zgbrhi0sOSmkwEmigw7mKDEPnTio0Fp3kjw1mL32Fy/BzsmNuOWfrHz0oVVqHHP8
CYo7MSjHAaoeWErCIcTgDhTS13INoYRirQksTba3ZIvr9HGbF7on3D9Jn6JjUNdB
I35qb1wGcavz7nyD3sD6qChBsJCYKT05npinxFVE6UrQW9RPKxsvjGxO1TPR9SaG
2zXYyqbx0NInZz9ic85Ef0X3TPJiL/Zmt+ceAtFp87xK3kng/349B0KWcN6z1IzV
aVPdq5i5Snaq5eaflrjg61LlT1dR+Fk7fMj2qr7MTnnCpDPXvDrFbCgqOUYmCt9u
4Y7cH7Eco8Kz8QP9MtQvwzWhShY06Dg//kvPlrSSSoBh5LvGQQcgAvlCysGlJzQo
0fI69uL6rZpR3baJyTp/NfztAvzTVkH35pIiZS5aEkaidr3Csu14+GMOnp63aPeI
zdtFw/jchxwFool0FZ2EEm/4DeIb47gBsIH9K1GzweCLLh4QRyLMD1U+emaEQ1Nd
wxtsJmKnM0fP72JjTQIzbnz38Um9+6lDkacMB1n2cEoza3Uq1BgZQO7zvM4NhGmp
9ogqi7SXaY1GYeOw6tzlG6L51KmePzvGpKjCfHSji462+XQeDVDwkiuI1GTmbS6/
dNbAV0GL6XAe7NNtop1qu1kF/6yqLiFxSi7dzCu/2x6NeTvueTEgTbUEf0vhKdHp
ez6nZkXzXnj5y8IAEJU7eGtF/Q/zEEz2a6fXhfhQJeha9Ut1AfoEAxiJ6Ikmqgag
kLQafCLdsV35LR1BI2L9Pn6VT4wjCeGW2uecjkz+2bNNYP5PgI0PT9WYeJbEtciu
LHx8lOiMTfXmDMQVdygHkRclWo4ujx0io3b4TVttIo94Ns5kBUDoVSpPKuhjzgV7
Lr6qMQvZ+CaiUlusYesF/zyCef0TjIfWXzL2Kbw8tuZ14OwIe9WpDG1ynLHf2sll
+SZ3HXg33QtYa4l0Pb9wLeXNGX2cej/fFQIbovBPCeiAoarmr0o+jIMhcF4DLGVC
xFDz42aQcrX72+2m2h5QDHO6ACZQ+rKWuCDu6lwoPaYKIsbBph9VXhiWTCPKlRq0
HIDpGkX7Nf7vxYORkct7TuBZuGlOvOoKSXmnyTlNSy1C9N4owbm4mSyjH4PxICoc
mc78MixGju0g5etKvzs5fAtED9t7IIXuTdppMzG7mwNHgCod7nGYHVTCKer2M6gs
biibB+hci3eVH5am26FfvSOYwmjMGTP7l8Z8089c37jecY0jWAijZBPrceToqBYS
RvNORzoYeXbsrVPRRZ6Tm112NTS2O9UhqH62KPdwUXBwxtgxdl/pkBvv58mdJHRg
lZPrjUMVs8DkYg4Z6OT82dlrBcY/tQ+KdiRKAsInev+r6JkMDBiuyGMxxt97u6lh
wZcE472YMi2snVkd1gK4vT3Svbv7cUWjMznxA/1+b4ArRWWBCrmcFVoq0oP9NAav
tqoyEAPN1pjDc8CP2XD5se17iDmrBjM5oBlltyvtoANXiQnCAWl4WJ2txDYmvy0h
EHiN4mZ/REC1S9V787UHhWhjt85POMHCkxbo+AWMmvzWsIs6jNNlHOZH7vU/BGVO
TsGze42pNDd0XRqAQq1W7CabSXyQWpHle7LzIxN/Ils8TtKamLuYALIXdn1MeOOY
s4imzEG5VI0l1VihIzamotMnNsYu2vBVf9UpB2oqloYTpvg3/uNmfsy36gyyo2aE
FvKKL4jDG8wZt1G1QFJPHbtwWf+/0K1YMqgz3Ma6zbAf2ZcruOgv1i2vraml/Fa9
XIiZJHtNt2LqcC44dsIMBzNq+FIg/CVAb3ENZiFHUjnpyhuDIgX23n1JKtdMeNKP
yrZ+1ii3I+CAJYOmf7114aZJsuEo6zeKtW4hjShQ8pQsOtiSvexWo6fwg+N/RSCa
4090D8639a4ZEG1K2umYjwQPtDQmGzoodo61Cpxwix2SFZi36OrktmPigFBBFAeE
3BMNa1/UoaYCovICxm9UYxSjqiSHFSyjEWxgi7OsTFim2rGWbAbGUHE7UaHc01e0
OD+6oXgYXyWGm3KHoHNuyf3aPXBZYlYzNVEPNrn39oDu23ZgNeBRi+b+TK2u8cGo
9pjAtCvd+k2lBLTvseWXEQNg4cWi38R2X2yTvOt9X1LXdJcgO5n03M3v3AV9lEls
lbpHxwbqOrL71Sizo3V+bl/TqD2vNNEDA9wajNCManUAm9Qca7OE/Ky2n/0IYK+u
lur5md9GXrDBz5ozARMT6e1OR2WN5Src8bKGNYO5W8GdqjUFFDK6G4NaXzl5YQON
japyNzehdcxEtmYZzlstOKrvRXbPPTcrmma3ICviNvO8x+WNsqH2Ap70GMHkhd+g
UHSZsnqfh13uBPyrNAPr61rCRxfshYMFdjHM3BW/Rur/mLFKLAE50Up40ZHjCfih
Zm8qpiB+LAEwzW+psiiyRMOuMUB8MAKAtvF0f0u1LkK8+luDzJr0igaPsTAu6l/D
mO//lNYkrBon2S5aHxFF6TiOSA2aDt6zlu9/xOFU1ZiQeWry+RPkJZV8oepbxKLh
0/IRO8KTe9KYlrYWTXRPswnZI5JN4sgI9+PgpqCwKIYGLA5MAiBlnnZfcl2WVM0Z
8ci2U59UpL5EcNDWNybjQFGYWRGpDZKKh+m9XYjZDHKc4oGWPmuI4xrknMsvkkWJ
hDa7ZuEFBhdghWWT7cU6FOmbpuUDQFgMzI5mW77W9OC0RNk8RPi2nZIK3sBaEX6D
HjJXtVNR0pKX/fSXissh6kgbQfWwePdWNskknS32Gl+29wsFxGxvjtxqMIboEn5w
eqNV7V/bEtiv0rf3dArtqdDqh5gNsNb6hWOgGArxq+wsHcWYZqC2H2Wu7jxKMP5c
0NCc1Wj9TxINDdB65M/C+pdw9vmyrFDMT2r3Z8iWdZRtkDyHuGZNfDMHQePga8P6
NGm5u5wOzH+46PJorMM9T0N7GZzCvtu5Na0DKpR4kUm/NiLxZnUhoVWWK0FMMZ14
q2MhKjYaqQ3rXUgSedKg1J4lW/s/OyyA/VbjsNR/JbziCZjP6DqX9OQWLBHyKsUL
Fd4pw4K9mzsQvM3y3vcZ0i8ul+MCEeqOQL5Zch7sbGscb05V5TC4os2q/CnwOg1j
aC64e7iCN3/KcuTabc6jDVKR2wuDjV3CvimxeoMsDJ/UCWAUSQP74bfgI+SOltR+
ZyZlUBxFJ2T5a0fYZwz9zoQhHqXk8fspl/5NI/KIm4xrAksFrUpd8AV6hxIOKZd8
dtthHKQRIiwKVRHHEhMiVZWl9JHydyz1JZbFQsg8VIjMaV6cD12e7AOPsunYD/xS
xJ6ZPJCtVytSOinc+n4rV22DKwmqIvOVCV7/dDRbd2xgmFVG+N8yqZ+DN1IvMlE6
vRpP/Je7oKq/u2j87vOS+eOALJKpMWhNM9j1qU8Jwbt93tEQCyKDnFKfuSwG8WQG
UzatHto7k32u7670E2v6P4MWAI19wesdxVSssZxkhFlFHL4IpLRze1dvA+4ArEzK
I3lkccCDO7niHoHwidebi78nx8jTcNZKP6VImH7wM/eKo8xnVKpzqwGSVStbIQtr
TiXMnhy2HWZWwh9wMY9g37EpUc+vlGYURmeRUCqMpIOk+QU84cvTiSSKK9WmqnpU
XWnKIwkk7AYn9GiCCjX7lANh/URb/P4fSkASwu2IWzokK2jc5tmVQXiRrfMXaewb
Prqst+Btzkf7IEABzgZrgPkCyil7F1rQJH9NcIwN/iLn66VZmp2xe+dtLHoZUhqo
Gt9TaVBgWKu3FOIXGAyJ3D9Jft5O4/bL1FUDjPquNNLmngSdpqbS80nMlaPSQrSn
/+X625YI5bGq+wu9jb+S7Knbw3RHYcWatPLtRKKE+PZxGfFuBV0m2650t0DrRk8c
+PRcdoVSsQfCELiV5WDiaP4hCasBQIJxkJEd2abCdCFaNQuCDV41w+izOQuLoLpe
Z3jReQupJsgyvEYMELBr4fGiZ1+tzE1b+nNmciIw0YGAoar8V0WHC1fUTcnr3aUg
AjE937dLqTT7KNFiapBDZH4BF+cGo23MUoHv5JmxW94elCl0qgw74sOkhDfoJ4KD
P5yY5MFKGdeH/jq+n6VnNeyBbhjsB4T6julaopDWnWlVe4r3Q3tDm0qM4AC8hreW
aQiJULsWvU9Q4m4D4H9gyYBhAioK3QjRdQfcGfTx3+uo+ZAOgRCi7V/ENTz2ohZs
IGyfKmodhV0NIf1Qh5ytjA8ZmlHAI4JaRW3Uk9BNwF9eFOA8bqo0VWwW8VRWA+1f
fOkKWc8mD6bDm+eoill8ZfgPaVk363EERT3yxwKMAzjc8EpNCXKwIX9YI8ugM5IE
qNGeWRtdiIh/MfmlguEgc335RIk27hhj+eOdBuGl3jMWwaR/BeyHaunfc7gVwe2G
ArGQ8ZHdKI2fxkataOMKVoYtQQNQY9QB4Ig6O8EQV7PQa8WJSJ2mFyQjijCiwL0l
kETTzuhwpBH98jnPhu7H1VBb9rPSsfaHIyVqYMgtQs4tIFtoh6wxmIZfTm7kfNV7
2nBfqHWXNOY9jtll8tN+50dq3PV3ML9bO8R29qpCxfTqIDa0p+oxKunRdaCUBnQf
XJMM9YpcjD3xWVj9x9q8CpePPKhy3ojc8dbn5Okft3AOFvcu7Wk/yzoUxER/aduU
qbSNmHAJuYnMYsCwgnBRr1In3dFwpyu3Qqf3GGvAQSlEMmxBD1uOAxbfM6oDsIVi
yukbr47s1Vsv0hQuEyJE3LgDg31Tn4mt1j1sQcN2KNZwqtNeurAFoMaTh0kmFmrR
mPzTNUQi92hUddd9U0JpLn1HL19yZ4XtMAI7+1jVeyX/5GKmzwELfcPdF0AUfAiA
C/mM387vOiYLV4sDjl2Ugv7GrTz1G1nwNdqLDDSCIwUxZE5SqQ+FvMexn9U++6mu
cF9+I93g6Z2WWLC/ZkBUirI/BxhnhMhXdmEBx6ekjD6HJnFCXiK0x2WV2bTsL4bj
fIMzBQj3XyfovfIqTjbZPBWvO6jltksWCc7D/HxxvNr+ZFp6ob10hz2EJKc8AjKl
sQASNRvDAw2NIHuO64j79eRJ64K6IwZpp1gD5AILHmmFrjEvBumB6wKuTfUX90YO
gEAcAl9dpR2ALcj9NZn9UKiF8Jtc59RhL4yC1wxV8fvbhKG9GNIbpmaNoqkkULJR
FrgRZ8RaSKY/b15YA//vomvmlytN2OWFI3OLmXdjmBQ6H/521HNaCom014myCpjy
JhsZWHIHoW7hUsJ66XeQaRjctmRMYyFGQjIPQ+defazUIZrZL3lvPrIJbqOuU0SH
660REolhvEOlnS7Y/3DdGjAN38d2uHv2FXhCGbXKcRbGcTUjgChRyTf/vVPSJNs0
p1CPISv1zyXu0xVI3gsPgz7CiwBmHGaH+20/z0CG5413EeFd6e3O763qhOsOF8c0
pfBHx0WvpLd4oLJXNpFrzQZSzgLKvZlEE2Oin1V6OiBzdk9Ve3CZL+01hfc1H0RG
nfpdcmu3In0Nf4NEDyNLy4OVi+WAYcbs0+TDfgI7GqhT8b1LD6RDbJyDutdeyhDb
BOcsfAxldWABkiJpfw8gZ2fuXsJnBuzQM08V4bD+bRz4Y/OGWgFiPh+rtftVJuzu
EYwn18YRE94RuV/Oa94WnL0dJn5TUkYyZfO2sBVHsiVED69RYIwBH1e/7M0B6ymn
oQpj42DGc9v7NxGZtLDCXhUDVKJ8KtdqwQMFCcF2/ICKjXeFTBJKUw0m0gY8KKh/
L05jw/LUPJgZQdc+RvyCuwEeixfMBFDSuP9kzGrdLgQ81y57cUJ/1zmOglN8vOcg
owDfDcy68bPkYhP+XOABiDIW4dtEjBj8Vbw84jiOgI0d8l4lh9xo4HLnTETaoaTG
ncfNtHd4ZF9j1EArQeSdsn3GksSQFJAIOzq7YZDW+b8DExaWyDz5Jt0hNXQIGB+N
yJPlpB7LhekShWUr16npSn8osJOc0ZakLUEwS0M51J3qMOl4v/byVETGwBBYwkUw
9+iCE0EEpel6Z/qlwsu6G9Urivht1ytdz9xPgMVihUyeHUwj/ev01WCxSs0533TZ
d7yLF9Q1WuQW79KvNq9+qipY03FSZ8wZVb0+a7bJIsB5i+f+WqqAWd5c47c0z2rN
HXr107F/4b01kRNl/OAoyxE6Bj4Tfd2jne1p5Wn8yqbf/ceIlhg4ncolilP36jcC
qsNqu9TPyya+RXf65e9anHJJ1cu+Yie8uz01rrPAaB3s10BFOaYIqvwoYzsCLvqA
lcbxlDZPfD5htyDMRNRbr6kVT4kDzhYXg5pilJAl9klrt1+FlB3KIKQ5cG/1G5N1
QsV/EUgeY6DOk1rhR8aqtYbzNFdAUvm+6Yu9sHV72pyppT1DJa5BT0RtSKIk/aVF
yUMPWIFAKLONesXc7VOkfbPURUqycVW6YYfiSUG/CBzkD0HMx1njc0OyXVtT1twQ
SVeORb6pFk/uCW7ilCxmA/NfklaRMd2m5xrZiHEOHO2daIwTgmDC/JXXWevK9IyC
VbF0MwsQ3nql5Cw5zYZ921UgEKWO744zg8veoz9W4gxF0YOhBbMYErkNFJDTuo+R
uygASSTw85bka88POSibEcp18MHIJ2uQRLN5Vl50H0orGq0Q1n6yOKzafMnlmmIZ
3LoFZu6DThS+3A6oQABv+LEUrk6pGgCM4j9lgVzl+fIx1d4S5hmULCMblJ81x4iK
nlG3V7R+T9drK3FRftnd4HQrEzctqtGp/ku2Wl2/CV8F0EO+HtFOFqkkiJxm5zTb
BUqS1FU42NWtDo7sUge/YHFs9tRJPP+pUfsVBZkF/y5186jlV+163n+tB3bNnOMr
pdePLKGyvcP3yE5Gr/fLZjq95kSTLUSkwGOUR0F/Zedhv9LKEXf2k1lz1hQNSx3O
8gy1DlY7B5OcoqhYxFcHqOo/veW1t76X7qUkWaqR5DGhAP8yDSZGLXjHKyo6+7HC
VSPNmalmF0Dt5wasdiyJZO9bByC1WKU0glVf7rMpAbIU9O39/Mn4uA1VEL8NQ64s
ivGfvFYyDXHoAw5N+ToVgP9FnUeYQiHuPUndaWTNL9i+++fhy/yUXfBZfLIa4rNf
PU4FdjKd+h2MA2YcldQ54cZoUeA57znOvjUwg/GAWItu9cVH36EO9L1MnxakLR1J
hGJR76jfVD4z6cpOp4AsgXKiL6sdPuXh2NCn1KdhXPpwdJxnHz2Y6Mx8Q51ZOXzJ
g1siBqLBZXoBRW6LpXVpKOwxnyLND9WeP8pHlsvuTW4exB/2TgHcRxcLJ7Rq4LCk
QY3MtQk2iTifSm29AKG7pZyW4SUGXowVvT6JixVG1pWYHhKl1sde7rQBTC3XGFDn
ogkwIalafqjYf1ITa2XzeNdrrSZ9T/LRFgEvAeXSqMPh4xZCxlTjiU9pUpp3N5eC
l7HtTN8yYHdNsU6rla50qZqMpDbjdUImakXVB9NjA7S57XItHmnAFqJhCitAHYwT
DcSvVxlFMWthlESn4R1EB7yv5REGCJSgYo46tisQtClPjhJJjOxlvzUbjWX6dhf5
r2KzjW9XEMpSBDMZTIzdxqsvj6Jgj1hL82akQCzuXdZv8ijfaZ3cDQD34+Ql3Xcl
+RdVkduy/X2kqoXvgpyfPK85Oi5t9Dwy4++80uOvoHJg09DWBf8JdnsaZHFjGu0z
hvH24V+n6wX0Iyq9v9NvHgPOUhx0Vjr2+P4zk2cJNlZCpRQxQotZ2l/MbVLmZlW2
aY/zO9PapVFm3+yMC82UDWjXhYDpEZAQCsYxxdpUEBVDpPJ+7zyjDU3+6eeOINtX
3RkY4HZ2tmPTIbVbYtgNbp3P+AlljwXF7OViIuCbaPfxzWmxXcwhN8sTeOCBBjRc
ngMK5sYmj9J6h8msrlxFzFefhgbGp6mvuW35QHGtBiNL4A07PniaFgIGDUi8pvoT
rX7N4b+sdM5ztZ29+8cPJmOZNiPemZofZuPnNgU+9RrixlsbrlJ/4JtupKwq2xDx
pAtEP52tSK96DVoNwD5NA3avkgVucgfsaP/xTNRa358H5fJ5RLE4nXTqxI0zdZGv
4GMFoCtRc5wdh48a0FWM0SBFeAGYOAuqORXaqeHljbQrVuVdtUGqnDDOiYcrQQ8d
GTEFqbVg4arR3RFQLMIXLIaGAXc99Zrib9V1h+nxqL58uk4z6AYDDhYzypl49VBI
WxwOfR4bPs3s4kJGBTO9BqEi3DCn+bXRSjJ3ShKuBJSchI6FwKYlrcBXvjTQ9e8Y
77wCJ6lwYm/Xrje3drQGqUcMgtQdz1guNSsyDNARF7aq22yDpA7rLORSeeXBySyW
XmtorLwwkShDlo0AURNvP/wLR/kV/NAycsuqtxrfw/StBvYPU6o0Jwhq6hIBUO1u
3gSYoDt29tYjl6rEN50oPGTUbbA8/ll8m5HSHOGo/Gn4Z2wmgqAB3XJJvmtFQjuf
tknh5N3YNz6LHnrNMDbtnfwo8drsQGDwTPS6qFryHELC1i3+vtor84iP4vb710eY
/ZbVrRUg1U0a+nyGMx2lVxVYySHvNs7EVKEO0EEqYYyOyJi/C2iFj+jnUk24YNzz
TwPLn/1ENJ6xAQnigDkXNtZuL8+tDsiwG4JW4sQ+pvpmlrUoMIzWV6MHhrprYz3G
NVjGFr9Cq/lYsP8T1bYP9JkIpf9wwiPCCSDzWZ20I47yeJV1kvdN2b3d0X2udZAQ
+4j9JS5InjO8EvHOSmIftPxXhYlPrI9Lp36WfFWgeLnq0SNxFzcXoxqJMlUD4bIx
xezxf0BQ6h07bd4F72zNVLRVpadn/YNdRwKMUEPAJiiMuYPulC2kvY+gYhw8r5B3
+VFfbi7y+3JOLAfygAhcgg2meP5PF1dbbOYdzIB3oYRn2y1p5jWiH/5Zm5nyTeN0
MFoa6BGBNFtobyG4xwVn+s6DaXFmp3qkDnzcVwYx4eJNicm+ExUEqkfrEgffIQ+J
Q6Pi69CF0AaouVYQ0Erk8g4nEODyqCJ3NlzLWCGPvXsMVRbwrq7QkMjB9oG011bX
NBQPzCDQoO1QTYelYqv7paQ+vx7+BWbD3+I50CqBdJEaywQaNk6PYm+sJP4my9o0
+n4ivTgUGoj7aM55XQIPJ2+pxQWLlCSXkYUOEtyUH7MPAV6NPeWT7bgv1Lw+9dgo
IbzBfZSDVlXU2kdS3NmCa75YHzKbgljdon/B+YtEwwcgPvFDTVCK6EejrMSKwI28
6Sb5GWx5Yl7Vbcg0nhx/qGz8gBSnB/a83GkuElebX1XcSqklWjKLDrCvFCVhoYsj
FRh/Al53hJwRF6JzoqbC7IbtsVu4+ueisFKG0Jah9rZ1xM5qnY9LlL3RdSxVKC5e
2Vnqf981z1ECl/6/REYptgY3ViETP4LOkzVefR8hlTXJoevxWJS5AoG7TxN2rvhY
Aswov9sruyC0Ac7ODoMSarafWlTPNpMgXLiFhgz/jijPmpiHqO0/Fzn4rxLc7lHH
yX3ghK8S57KpV4lVyOb6n2aUDQz+Kxcyc5WF4GT3hC1JM1wBk36QoSrclP1SW9B9
Y5Zp1KgflznFaxroA88c83gED85E6H/TuoqrCYhR8klRwHVyvcxA2pYs+m9H3U95
tP6ar5Lnp/eNFCMw1b7MeDBJuGDJLylZVgfshjILi2ENeyGWEt4LhlsOlndIvYk8
I2Q70FE8vLZd64aEYjAlHEyHqgS+Rx5K0xs2fOzNcVAZZONaq0C80m4sZDiRnNzL
ZxMREB8C93oxNJ7zcg1Erisq1s5Gtb26Yub1DDi+4/5FSpJzg4Y7MMt6q78/kj5H
Rau/+Dgb34OMTpzOpV0ty5OwaMGGjNOrz+FNRDY2dmh1HKB+0bKRDIe0eQ7/NEsk
mmeFFbdN2EO21PKvyL7zue5oRP2hUyfCH9OdjDC87ClEb1LaVBed8lbip0qbGRdk
0twoJVCi5SyVh1UPRVyjS9S0YiEfgLeDM8/z3z1oA6zMpTIDVKqnbcuAh62Lk9nf
Trj/jggvf9S/GcbrymClATRBJL9CL9esBNQNx9Ep4NKiVLMqjAGVbxW7Z5oVPzJ1
G7U0CdA4uo6hcZRegKDDNVgkdWcjnFGgXJd0v6yKLVaXzVViAfALco0HVqF2I+TT
aQBnAiof56uSWNhikypCo3KFknEqazPD4VVSMRieR/5Ocz42qIPLh2OJWyChPi0n
XZT5cUqdq01kbip86PwHV3S0wSq8TaWjyRc4i9wwXQeffVqCf3oDeqRJSVde9d2Y
PTYJRewEAvZbVkuXSsUXQi9oLhIW9YqrceNV9Mq3W9E2Eblzp/DIcDJglEBaRvSR
pJYsETLstDK96BwmLlRq1utpdbHS9qNB14cY76pbTmxxjPDKG07JTEdMjF1TAAy2
qzT47MIayQiLXMmKiDy+H8zi4VR040BZAFlq0m8Z4L87A9Phjr4wn4n0fOXYHv92
4PrXBv4rYAutJTFMK9jHS8yfTKE3Juqbgpf91Td4c2tEfLQF2a3FKap+E/wV8jFT
j3zXIJuRjSd7RPnqxVDS53QNRcIfNkfgXrgZtmjIsX8nnPbiajDb9gcgUmmQs81t
1kJgJ28UCVO5B26lq8EfcBfG0W70qF+9rbH3lIyZ0nJdHcWmncDVxMYWFo3ak2B9
wJNABVsF+ICzCqr6jFtT0E/fs6e8J3diKUy9mn3wyjF3jKIqny3axTgNfe5q5nTb
+O/Jn3uYzvU0ETZiXixy7eyUgXdRqm/j5bCAloIt5qCC7+u2u9jz0cwLJ3mw4wAg
FHwPZmnM/0Zu7kSXBAhTDnWfQsZYdMX6gUripfF9GNfmtekZDHqQDvfZADo7N0xm
POGSGDs5szZbuKrWS31BENoJMmY0bdvMP9YyDwd4l4uDXEJfpR/DP750xawMmn4x
eCRriYfsbdT9AFpXobqzOrmx9jumP0HiaN7I05lSbosiFl5m+YjRyNN73A3PaQPy
FHBX32FAO3/7PWU1p0wMi6Vx2o4xKSgzvYhYdG23sRHAV4Z4A4L2mx6ZfU2WgFR5
1dW/tF/B0SVqNwA5Ax4tDzY+JJ9JZrLh4dWs1HIlvI01gSMgtLVRKyXnIVEwaHg2
p2fcqah14tjGOU2ncGF2JUSvMsHMp9HxM1J5QqZ8rMyrOK4RtTxyEXMZ8ey2Ocnm
RqTmfLh1SfrxaziBUi+/NW3R9rr2YHDmvbAYgK46j/w0Kr8Yo2eMifb+XqN8AuYu
746oJ94ZzMHY3XdYm0Lx2kREhGbMzWH5Vi0Ho/8YFHTUUOfpc+0hiM53gXn8T9JM
AHdudHrD+k/iQNZnamfLgYMiLZKTMLXX5mgJNGWQmRrzud69z2ZND4orCaowC1M7
dszbMtPKI+VNqctAIXy3dyu5Uld/H47EOGtJUotujt92Z14OT/Fe9t6Fho2Nbejo
rDaFi+3w+6WSZ1RFgAKj7WphWvzMBP6RO+xviPO/sgW6hqoQy1Lb5cJQtqwxw40B
NrG92I+IC5yrOxR+bUBWlp4lu1cm012ej6Z8jHvE1L+RezSguJ0ao69JO1LtzFOm
VGsyemwd7fIe4WnY2f7nY2N0OEqwBnwP9mVKltyre7U2rAK/cBMHVvSmGfpzWKc/
CYlaGJQoUjiUAXmuJ1sDw5pIYoHaOrOoK64HoORo8YWcRilJo10imX0lwJPfrSw9
OQ/pVdBKcxN5vURyQeF+Nxsx+p9xPU7y9UQ/RmV+YzlFki2RTyRp0RcGhI3vYrwl
fdDvOj/KZJc1KPU/oJGKS1cZXNenjloOHZxmFTJPbDF4wQC3igd+8x8NAdCiAeQO
oX+frEHZ7qiyHyPxzuYHhXU14CNZ86VCTMmxRGCV6lvOh5W9sbrFTklq2lszmfFU
ilbCoZYhpw6JUXNKHa54SqgKtZydO09pr+mYajsSb2LFqV8eH4IOqgvxwlS2kWkv
UPrLx2FMwS1VHuvufdU2yCjuTQYyjXDcPRVwxU1vMPrZr+xFTapIwE3jajYSJmr9
X8tHeJa+UvWXNLtawyw6HyzfOgz4v6Ks2r1D9ZTet3p1aVz8XGASpxw+Twisjp1+
CXRPEStcuRh8689soCjzOLMi2hUpWFTX72KVy7RT633z2p7D4lAr6kEZzn141O67
8SnsnJ21eQ5O6HzahDbj5WlsEtdjthdZM3NlYmsm89lJ4tsCrnGUION0No+aLXSW
9pBVAqaTGnslQ2jZbUNDFPx0FYIyF1aaHMFt0U4pGKTq7EKX1vM9vv6Tsf0pJacz
UlWVFqL9ZrE0+bmo+7ttKGuA3Okdlh9xXL+EGH9EuHnAACZOLgkVGWGYVcKg3lLa
NoVNVfpyjLc79qUGhCaaUV6LUBHWQEKPJSqKXlZi5XLJxZJlSCOMyFZ8Cf+s5JDs
H4auqhi2CW4lD99ZJ4ngzE1607oTZs4BEsjpSaQc2nB07ZUJskfTMN7TJ3Fey2rX
MsRQHlfBxyjxqoo61C8JjwYeOwBBOsGp4kCn3mKHSH5Dwe6x8WPnH+dKL7yBpxCW
0QWsAVMxODi/h3ITgdwPuquBQsRtd5MyGdCdB5HoEUJ64I9/m8kiJv4ABH77/rOh
KgYQj9b0tehRZjL1ZaOG8hmG12FBG3TZCl0GIs7RUwHHXyzUoCOjTdFtxImWdlw2
c/k6qtYCJ29P4bAKtCY+kQJy4lOL/4aWxBmsl3KDHMYSPwYFLvadY2Ulkbb9Ey1K
qS38kdx+gI29V4gPYdcbvqgssP7d5gjYBl8qpjJS5+RMvCD8w8R4ZDUpNS1A2waY
mzvP16zzNkitp2dP4OujY+q1+YzEpD79rkt+8ZGNlgOTsaMLFasUtZxeZ8mchMvO
11U1vQOih2MHHsry0SolKeF6nqSOfH4rRiUA+NFhzLXjpdUhgzM79NmEwZYLQGAt
W/G3L+F97K5lpjw+qtJq8Yz2EZqV5fagar8mYLF8rBFbvxIYWUGPwBLGBjuNcSWT
cvPzUB64tLTFYCJ/DVGOIhf7XoQ5va4Q2HP34KsmvoH7mRwOp9C9/vkTNEeXYNi8
w/kXyT1aHeKCHBPJBCU/0M8CT9ddcHUkymQ/XF2nYB/+CWryLijgbM/v3a/Z6i3r
7L+lGZjCm6cRJjcXby55HcnFHKwx8YbytUwxkVD8xEuTw54frE6mvvL6Q69EVF2e
/6IF9fxttJDng8Mgeovj/uMlCTA6rQ7aB4qf/kPU7Q8APj3puQ+G5GDKJ1jzEPgp
wr+rQBAKMtGlYJm9umTzAc8RoKJ7GbZburScHuW3xVzjXh7rucxQP2ELmCXj6RkA
GY0y77YntT2pY3y/oneV0qflCSkz4gneLaoJea6qyQMHkEyzhK6oEdUp6vhHmbSu
J/RNWI9XkH69KUXV+ZpHFd+kGdO9/izsDT/k5ujO1NDBrWoB8rdqxqxHg6NBS8zh
mIaZgfRnBe+M+zAYKVssZdnsBYTRXfaJnxfukMf+EsErml2wQjDUlok1xR0uu0GR
mRzl8f8vXELNGckor2qo76O3ac8ucxUBy7CWxuzYXElBTAr7Bt2+GgPFd57hVaak
QdN62dcEo76U5UE3IauVrGwoS1yJxaU4njCCLHWnl0Aq5Dw9tizZv1BjiKjTnnoI
JvTBk2dkcqMXVImfF3e59V+4NhfqwfpoFtLODMb2nhpg/FrmzNVsO4FbkiGxyNQb
Vffdh+KxZ1A8gulghdEIIzPm7s/uKtw8b+FrKabGLoyl8vqNYFqMtzPgZNYUDFS4
wCIQKndLdIzWlKPHkoZarEL/7SW27NTgaI/rUQwOLIJKSevKd/uYQTC4icJDlCfa
hWWaTSm7Ui4loTgI/sWZMl99tjyuou/xcvFsTjJafLT1F4UoQAoB4DKRpKMCoqti
nCQL1VZx+fmV2C+4i5Vlh4sU+1ywa5DYu6e0nzZY81BAmSezLBUDGHpi0m/tqOTc
3a4ytEkpD7Y48Dt3YY/CfweXbXwQFuAhXFPysJuQwUwNML4KvMIXQdsXm16jY6+j
vJ+U1ITh9GdKS+0fFn+T4XnqSuLVLXGXM0fEyOX+Ml8U936pyge/K67tGGlpM+5J
rVbCAQOg/e13AXxJLE1BjhsolIqV92zvAy9UvT2yXe0Q2GzWOFl6Y9yAvb9PrOis
qyQJ5DTlzlqmDG+cn8Rd0FTeZKIuS+QQYmYNb/RsVITLtQ1PBPBPUsOyfbZsnjCw
Hl0oeTjnSqtZhMEvDro93raqFeDGUmFpsOBKb1bv6C8fdCY/cE4VNB/AKpKFjIYy
Gb39USwDX1hIPQd+Id4ztNgK2TcqsY1jiYfXjRNFGuMvyrLge32Mg28upQd6IQbI
W6/YmHoDaSqDhu14I+8KjGtZDLPlueegKD7jFDRYi2uLL9EP8gQiGeDrxKVv4i82
MuUWDvIDrLpb8phiLCir6ufgbCvW5Dp2pcpSt+aJ8Ji6ekRYN7LOvdk0nMCgwaRw
kK7Lmf4rYZBtuFUAfSYzO7y4mjgKfwwvc4qeGjoItf2MyRXNZAh7KzKMf3m8T+nH
Ja53o/PKCmW6pSZxpNA4xQXyKk80/beSwhuol485bKlm59X1726EL0DYpVyphXcd
ksyjgjUFZD+PJsg/nPXCf4zDoixO6n77YI4N9Ewaf0s8Hw+dCwXrWqOjpA+TIELi
dU/8YbydCUFUMpwnU+Im+i11iyPH7N9QXNEtTbzF9f/abS4Uzk3sqRpthSZDah3A
uSWPRr5UuUCWLJmXMwEA00itYpi5QuOyWTveFQcsl4z+/e/50Ozja+zgHYIEfV++
SwRmsRBm6kF2pBS1sCFy6xs+58GzQl56Ibq0ZdaZbCA34e30xTV8k8UlEIo67nRd
kEXq0IxG7oxf2S+Ory3SksRNRLNrhGwrBmud1awOVbGflJRCnF49W0MRZ35uZTP7
woSzkg5d1piSxTfgmZ1aub4VSFVRlu1GNBUkQ/+RVkGJYtqQ7RyzTLZjp2QG7uPM
y4Zl+ab4omTCB5zKl60lHSWgq/+FiqZLSxwa+QbevH9bHywo5TQn48BUxCj3TIEg
gLA++fm9ewc0+WiVKw6NManF5Fg/oP0S3zk9fJVBSD7yOfoKPKV2hube+mrhPtah
6WRRQqgF8qtijYeahRBQ9SFNanw5PlJ2eB+bmldMOw/BmTc8C2SUFYrBMCdlpYIw
8we7UlPBwA+c8DpT9ZZvO1zHspADyFZ09w4Cx1iDbe1eLNj2o3oTgKF+eCxDs6vK
vOLU0wpsc6huOyVHiFScOPBwaEW4azr/oL2a92iovUWcuDi7NWGMwtaUtF18WPFS
fipPXqPU9sTZLwGUehISL+zgQp701hkfHejWcZI3ZbEbrUt9FklXYuMNqEmhi9Ph
/7XpFYi3dawolzwNlX1uZSzgq42cVF9ExwXzTUPsbhiuyIOaIUMB5x9t7Y0T7Z+e
Z+Zu4rePUdV5XTcq9ZshimzkiNWScvLX7ACCQe0R6u8kTq+/ewkrQxJcBB+Xd3cJ
K5pFOGIHWYSzA7tcnKRuRa+MG8Xz9X7iFi9EA5DPyfyLTtPJ+yoDmDfEuo0/AfiF
myNYnU5OnjAJ2B8KNlSypyAGLRUEoV1g/rp4YDm5lVf6fqX8dc4pSOt5BsW4VY4I
lADIiVsPfbrCRaHs1TsxuI2bYt1Hy+IwAvoStUEWw8IurT45/SfhMptDPOL07utm
3Hr7o5vfB5Cpxv9T8Z1gmMbcdNNGX0Zp7p4ASt+KjwYULWKYXQlpazi56/PmdeDE
bF/7OcFJ05kLnr6rB22ANDlhPAxultA5AjVj9ET3Cz3k7e/CdLBEGoNfKfRUkGH3
LqnZ1tMzRCf5hj7vJKxOyMazSkAH6ymW5O0QL451HmXeUKQq6THowK2DN2+nzIOw
BLfHYO63w4UXDriU4Xn1gVOQFAl1/H+14KPyt+36glFhAgcKYkVXBZ0MD0m0vSCl
+VH9WqSGGQEyPJUA91+9fuy6EsDMS8iJHun+sdJtC2q7UoFkUbsP20FvDSAv72+0
xhiliB/Hn72ESCEXf7BWXIQkiFkeIBSRmOufkYgMhqKHXBlEuy/83LeoUUrqENVy
Rh6AKYks2eBQrvh0C0s+JsTcgW1ZxYVQbngKH03/YBKtk/AXiWwrXOlofMG/EjVw
ZevLkoAvzypxW39i0a9sh9zokCQ2C40d3rdJ+NJMhIKHfcB+mZeXLNeDc84wTCPE
U8AMImaHQi60R2t7u7ofzF3adcMZ3enoU2u1Tj6t8rl96oFYmL2zNpIHCI5TuMfU
ijOiU72sj+y3rbS8l5gZC26lMbrnt3XTqSg9wLt9EHa5gY2OTz9YY8mrZgaNAtol
hdx0STGGbEDILOk5wScjkDPqVQ2YSeq8Ivaci9DUw+7o+EXJBJvTlVO/r3CwGwP5
8ovSfllmCC3vMX9UVuHPbbdkwfdpgKqYiPQz8l6K9vXdGq5eMhvtE9AuKOb3Tb4H
cNAxNJHV3JeK+FVVKo4Cy+D7j126CONrmqCyWyrHuBBgfuBARlEYj+2RaGa2/Rbg
ouZFXlxeD65mjJuRJd+D/JDo60t+noba6XYdaJV7Q1YdDw9rz4RIblC5f+SLBAbe
KmJd0AzjBDxrPbPnH+jInYmN659I6OxMHts1WBM5rMwY5G0Wf1sQDtYa/1VDcaLb
lpvBRfTrye5jLzZPyV8hPJMbsKA+kijad5ZWmjfnummlP3jW60x0rTLgKzvX4OOY
ssNvWHdIAwf4oL9AI7hnIyOc4/90xDCWww64/NuXimrMbyFdDIEFAnYTjqtbYT5g
fp6Mp+gq7UoCO7YdR9oZCtFN4lckbgammq+87g6EsMSGhgTPZeWGKdNJ4dglOqe0
Q6voh9WcX9IjVGjIUuzMFmCWyO8o+BeNGvCjDjSHlBOBJk/l5jHdnE8qJamIpX6J
nwbrU4PiG14jmrhySH22aABVTbfZC987w6c8L3Y1hHXYSLOp46cqCUzIyD3rVke/
9pXbomoGaKdPLzdGeWioEVeoR4m7Q7EeIbakbw28UVaiNx1X6qVPhZyxdMqpjgJs
LuiwwLbqtb03dpsNDimtwtiA6kto8zO+6cozCAkYC8BqdLL64hJQG3RHw8cThjjL
QuKqMUecMF3/KTSJulV1f1LpTBmj4c399ysM49LPf+Vc4cW80hlMvwIDefpHwyw9
0fYLQ54A7cTq9Y8oXUMA/8ioX2vENVFlEbhu1BCJrPKD4uEtT5yqID3DLd4KRnmc
eSvRk+f3kAKg4mTsdGwbMRkqJQOj5lCDYGc46mlIi2p6sVaMEkfQb0b/pGHmm+Ij
eN1uQk1tB50pwv0cJ8LNsjtpWin4WkStpwLRYJZj+XE0x13cshDrk0iAEHjI5zDY
2faKwDG4g4i6MRAX2FBRF6hdYHwo72GNebqFuNTtlhZtkvw060TVKFGOrsk34eXA
IirDaUUVmT7F5w/PmcUqzVPA8QU+VFcDlyYJCJDvEvT1KzfziLhEt3iBTwXyJmNg
Pf/EYBeyOYH4li19+tTZMW9XMVKOg+vqRNg1UFsKZtEHYUjxabhkbIURGBBe2Y97
EEm1/RJQO9oinkIZ8t/sX8Dh3p0EXd23gjLlYQR+Pea34AmBCUu6iUSJh56DyIXc
d9oF230GTGxkjiGM8NtPadsWDVt0aaswXg2ceyQvmGDJWhqlGizmmTDEqrKBo70j
x2OaxDhn5WTRvjCc4kYw61qpNCbs40tYZfzUfWzCIecYjKZ1Gt/e0TC1GbKZGZan
7f/tlRnDv4+CmVtluUDx1srmweoIrjpimUjmWcmDi0f+rpE4eSIvmiMxT45+D2EB
MykpfHwtsC+Gtqd/T0JcvUMNLZ3gFL/C9y81ELvADYpm1QIK0orsyoBvxG8+TgzH
xf9FcOqVCrFpZGUw9eBWGeUlzKrZQpjaTirzvUy3WLbGiX8k1ypfyGBvMHBwWzNf
EG+22DQSACGgL+/cNhifEQyfbaa313y9XhMpb2Yhg/c8jb9ZRZXAXFPfCluqnqSE
c65CCq3L1PWXP8eQV5N1TcStIlig1FGB2q78APAZylf32Qdq/GsxV3fs+CD/aIQL
V1FhqiS2Z+//egkTRZSr4P/GEtcMSrtVinJIgxnp86kKYdW62obo92XTwcJ9FHz3
UIc24k0SUbqF4/3RGMKEsNX1ioWA/ccS4r2ozOTlGIyUvUMllxflhGK5PotbNFjQ
7AKLN8WiChkF5vr+nIIYzX53hl/JPdCcVmjVyFPJq9WAOzCwoxjVOoa/YL+VBF0Z
LDj4463CSj3eDfXwEmR8TYrAdLjbZTzn3WV01t4EQV1glIsDV38VwbhluR0td6CX
lUk4CnNMi5iug8JngV3HlT8PwNL2TCbY0+bfQyQ6jtKW6YMo6gMSewaWZaWf7+xz
jnC8GKbgxMzBbCGdFiUpBnss/fpd2Uigoc4zMrYC7vfH9zjE1K4tltm6n6f0LaSL
6y+LK63ASU9Nqk1GuWrIRCwFgW7yurQa6vInmj75MKtGNrQwkG0bNt1oxYvy9MR7
dl4hDLEk+mArpKWFDDHDQeKwSXP9cZOvgp7I4IcEsmkp5pu9rdIosH+PD6n4/yIa
cWjLWgYre7NjboV9KLJvNj99hJmCeaoVaB3AvojwWCdqq0LhNk1FiG9BkBk0KLw6
8XH609ZfXFbVXh+/DObhAVpv2yMRudKD+tQG6NB+xO4WZb0n1cs8U456IOtN+ETR
+Eh68B9RkkMYH2egpefXknkOOpWQtu4jstSi6XAbTQDZnw34ssT8sDS3B0hAeGwn
b+ubmpRbQ0WWQK7VIOuXZBaKT6PJPtZpLNQapMrS7KZFrpUkcf4EHeLfrRMGZUyI
hLWaQ7BabPSc5bBrvXQzcy06YTF6rvmk+1qRgl4B5tdhq6qOC310o+kYeHkeBPeY
nVsFgh68Qhy5eQYN3jlOlOk5QcqyBn8G8kRB/TdKwYAqcjesRaoNg8mSFochrZ40
JPwvhojRrWBtyAeZrgybm8MSr/jL5glNT4ht8wfgm9GlvoVkPPAxU5b5G2xy+dkA
l4yjLG5UB6vxzHynVF0K+lpk+E/A3dmFofj1YR3JPtL+IcyT5zRl+pheMx4s1lJc
CJeB1wwJtyrGZkir7r0g6EKsMJLVcHueM5/X0t9OrgBp4aDNkb2F2oR9qoUvVubb
6gJynwORg51eHNidJQtVNPvQL5CXcLxRmYeRRHIJZkBSQ6hLU9Ajml8GtRWdo4Wv
R+2QVPijYWRi3wAVYiilOAzwGO1RTrLOOtWPD4W83OTNdiIx0ArB6WPa2yiGGdbR
hGI7tiYRsY+EN8HXHriXgvHLQQosc2bcau0IJRm4zO8fMtymWGaQwAm/GRQ1k0km
Pfmyuus0N+DBREonfc6QK4lMxUVHQuS2Tc1u7crtko2I1kPAlevz/saFNT/v5NAe
T8hdGigbGYNY148kNgDB7DfB50hyB8IqDjwhvaNYJuXZvXiGMqhq1KPh+Klmfn42
szac9HRhrqDOUCPW78BlVtO0mRC+qFjMcF764HcOw2wMNaKxwXSCfTK6DU66GjJL
j+ywzuIKoKfueQixfVrDLOh4kCo3hx/q0R2DQrlRaK9bCDqNtqVEM11pc6yZ5G8y
Swe5drFZldoLcBU992MNBiL43oAdROQxhpSiVegukkMk0gWoMQsaQ3Rb73M7FeXP
6WFMcuh2F5oIRlVsR7zsnpavkYzw/jciJOpeFMPw10xvyBiFG9vKsHI47fvBM0Yo
rdqfmUvYOXzcy2Y82fXIveUs//kaqV77/P62ZwojyVvIssxPI7BdadWe+Q93nofT
yn1SAHXBfdvCL4PEAijEtjGlPeasQN4JPsQjGkltpj1n7WGKnE1uQLQgvPY6TdbN
yT8rutINKG2rWhb52f5fC0pN5Uh3DmAWllkh5TJyKy6dRjLWrGkrDQcpRWTUyQMs
25St/+VhksaHPngEu0Qigkix8ogKzwY3JkU70C3hjmy+4KuooRFjq44oD6VuT1f+
ZUnbpmvzhVahySmX2HXSn/FFJB3jM4ue8oM6iS+E8bUTCRqk7U+vETCKd+zBLHmM
OF4SJsgJrId460NnIPzbpDft7vPRM5zH/bDwkoOTuLG2bLWK0alS97L1bjLsXJ5S
+5z1h8+iS4pRBidDb4Q9vyXfPNfe4POKAtfGJZnsCItpMFxUykrnT+M9327CVrqg
cYRs0/6ExHtHVOlvhOxGqQKXi2hEqgyYGzCpxdzppWTPQ+sSA0LJ0x59exOs0dCU
g92eYfG0PXTkBNHiIdydhYKQrg0SO6n6i0j8zJUlqv0sX7ko5pDPAJFbsVOrAgvo
8wNLQpiq9Vz6GhwzaSpDL0BVmBlD3E3Ql3G0cZb9G8dcUfmEoiu23KvH3JBCguci
ydeaxybJucFlHJarLXqcacL7nbaNY6pmfEjSyMMCqRX2BH1MZZY6+IMk+KiunlHh
S76j9Zo+TnYJ6dRD+y5yywT0ljKY0N0cmoYG9aYIYYsRheYegKDj9o8qag3eXXnr
8tnG2GkkmaCYh1C2eDsziw59JcM0insN8BvCgS/Un69yFmgipkdW7psyjNVKVgxO
WwO7Vn8pGY5kQQNPB/OAfcPgU37kw5w1HdNtBmktKHeimjku2Kp6zihLPGwq5br5
SdPMZnCHIYNeEbBdVGYy7yLXV62UdieOKBMhtwMFARSs2kJQ/GTu7nnbmd6rdil7
a5bSH5wt60P2Gr2gcuu1xGQf9K+fKU9b69jY6owya2zeapVyyEB+Q0W2VFersRAp
X/uXotzhObxMdT481YKIXdldPPQ47S1kLmHG2FMTMLo7KjWaXFB6XBGa6n7Zvp04
UjtHcdpoLy7fB8q7w62jn3oLkJ6Lto8cScmBNi7pMJYcuBMaPb8Twr7j9XgQg8JZ
Q+zBBrPl+maTyZTgeXuHAj0ng8N2TrhsXQk33aGD0iYu+cpMhY0qmDaSuXiegfvS
kqoxstBcahFTAi3rVG/xp6nfAaGSvYdkfeCs8eeKlbUm+OXTdD2+oxx3+c9OOehh
GlH7Jz3keENAVRvBuHGJsI5PCOHzwyvypSoyeMtH8UWyEGjR4HH3HUVeUlB5jCUU
ZVGbs+wPVWseCt3Wncdq/Kq7jzmt2UyETkMtm3pZei66Q0lI4rSKuJ308xi718K/
Sm8LmbrqtpIjF6pClwn/e+Qh74Ugjo5XTZz4UxUKVBQBbahsFRMVo7taK2FO89jM
2uEt8ntRoR7nLN7Eczj6Xc6giYBkZ2/DNXpLIbqkMYzQYLKrx1c79uX9GoRkgc3A
Jh9TjClGSTyo1hNJdPYhK5WyN7xI83ULsorHIIIEmk+bePrqGmEuLp5raHZh8avR
sikTGBPO3xwHmCVMlvdN2zG+oRdOe337G0qJJhAP5tCTulJW6VQuDektekcifaUS
nr/cY75O+x6K+MqDQJcsMHwtw7iE0I2QJjrFboYoiyLiwfUtA2ktZdI5BuNvCMQT
uWzySe/QEAy1fXVRoIHDB/ipn1cWmOYGuGcRSy0yT+xTq9gZ3vomglj909Na2/ou
kJ9NdfUI6WmFeRSXNjGRW2wTSWCkCm7v8m21NlLG4iVY3V+4TatE5ZXFWogLp2VX
olL8UYXpm7PV1kv9DXUiy3xUmKQIXDMrfa7728K7zKwucH0kqA/iyzyCiQM1Vg9I
JdjTmqwNzN8fbTtINaybKYTO4/e6vjKnk0cBsAa87XPIOJRVaUPYgeCEz4DNYpYx
B+V5ZLmyEgMNaVkD5N52gOHKdUvOvQsg5hFQuZ3QnIWZI5frRpiDfd2XJIw3HJkH
c21RZWmFe4GgggGve0VJ2Y58rkVDj3zu6LNzncwkbM75oWFHq05pJFLPu1PAhf0q
prleKBq6orzFcldhgACwoxued1RUf52rDf9Up2Xc16JrWhzG1VGdboK9QPKlxclH
giilTvbRMLxuAqo8xHBdqr1PVGoMJyL1u7/FdOq0gUcDts6nyC+nPjGhT09MhMYC
KRTNHAn2LHVddOJtAA33Ke5DaTVTZalGO/cwuAN5HvCzVmqLdLfdiHPcITUT5kt/
BZZYf9FSKTl0yHXl5viaMQ4Z0LBDQPd/Aq51ps3M7qnCK9Mw2cOIJxNVRXxPdgoO
TjMIFparbdrdstRiBP5f2xlP1ttMyyTsHunyidRjibLCSuikPwy5aIPiaTreJkki
PZ3+1xnMJPLZDo5fCvUhlCn+ZZ4zoZb/5Vk0YSPMTNPzHyPZz4g02ZyV0epb9psJ
4XJo4MlQypnbU0nkAvc5FR+al/Fn83Nufx9p+ZWgJy+iN5CqQ4gwGsdzWC4F9Dcm
P1juBEOSv+PKQdVpTDjIBjZ/mmW8piXRDBhHCtUpsnz0YLJbA1m9eogb0ZNYPfHG
Wae9RH22F5dCKM1yDXDjGUwQn/74y6KkY4EJ80dRnZ4yqGjWCo2W36SzSAwwfptz
/zGoPHZNJCVxTG1IH50Iz/0t0P6t9GXYmx+/Ts7D8OZbhUlSSEaE5/48D8GYn63Y
m/8WehbiQos5B14OBi+3ihFfbn0MJPpuA3cdeXvj6DuJ1TYx5MDaG/nW4vS76X0q
7T2kVSE2Km81+H+c9F5bv18XIMl6fQwrAgw42W7DeVvkvYY8CwG0Wb9449a3OsIS
+oZuCbIajU/8iYd8mUzOlsCsWRytHAAYSNVocLbowy02bYz76QuZfWERdI7iwUut
LGeF9D5FCFu4SwWCoGenrssz7aIiNfGHJwipdR4oE5ICkrBrvpUBl+J7wktVAtuS
xyZHdywXznUbpXxVzK0fE9Q2fmVdv2CPAYWaChjLlp8u65q+i/PFJqU9+Zu0hiRZ
IWOhTrJeDPHUnSHIB+tsazxdr69INBwoIWy0acIcuBys4ouMI3/SUTFq/mVkXGjB
1IlTZmEy7MyLJAVrYwRNcfM4/9BlCBq3Y2bG0Etkp3p2Mfr2hgoMY+gk4QXi4Om6
hA6gBYIRa77iOpy0/QWPl5DbFX1UPPIqU47/6Ic6DuVGATacn9X+zq3HWb6dhnm8
XIXkve3tGEGFBf6To7sjWSeuHvASwkVYPlguUySPOEEYKR8UGd7rh7mE3h1b9F9/
URtkYS47Oq6MOIt5lK1cySjGuB/XghilcJjbwrBcGOPNYBlQMiFam4pzdWZnH5mB
Xqc/oEQA10zMiLZq1azsaKYXPsmu01+H7ZgNjFDTOqlOwX19x3GdGcfEeSBlmi62
7fIdn01hX8liiQ5HzrtadRCoGhE/N6uapRBlS9ot57tdg0PMYaEWei/BGbfgOWuR
Fa8mmd5+kLdNp6OlZO5Ol7uDs+cwARyktHpSDSHtBQAkR1OtzuaVIF4f6QI41gDb
cG1/KVmGIkCMrgu7LAUmB/Z0K1OCBTtQ7TZCEcICjYv89im0Q2BzhzC+/Sh7dVOi
5q4GTCQPb7JRRpK7rjId4hvl9GKamaLTWiiU+kPwJa5YbZPgeEg7buECA2THnx5I
fT/ETzYQ5odgoCPpSXcJXlBryGPe/v0UMhWhe7sLtHD+F987HwM45qlmli+bVBUm
5Y9RyBxffxs1oshEkhhx/Oja0+QonigfvGBamT/iYT65o0UsTCmKqbQMPPupOp8F
RIzQzji1tzf3nZXh4AyA2qo30fzBRu7L9fDdTtvg2k0l016J3LolpiPKWgL+JPs6
+W1nZ6ZPs8Rn8F3Yu2nmIA+tnK3cEMinUxw2459ff0mhg0tsC70CWvEzBxS8I9tB
sftznY+MxYiqbGcDWZ3MaLYiDUrIadKdkDC3Uua1xk86LaF8fT/nM56txYONPt+8
XCfRAPzTGPyY0XQZVi2gSFMX7ycUdE7xpYTzg7DhNlc00U+LgIKEbbaLUgyADTrD
0g5wUiAKZYDGR/WIQowJyDPdQMqwLlWv6Jfy38YVnn0iXqnlqo/bw7O80n9F1C5V
9xM+f3eSjk90BuIHlfMIFbOY/NZTb87MR6HiOonayz5k/ZX8jLbv1nJyvGeSlQG2
mQk90H0kv70Gge1JK175SfRuHOI9SOgksc1Z4QgRtpnaVfx5OHYQ03o397i1+gtN
vOIJMVsIbxrX77gjum2CUjkW5jT2ax6eo8cRR0uXhjGnVGd+2f2WniHw2huZtemn
m3T3bFmt1/KPhs5qZvdOS8f6AXaMOykbufe5AludxSzCNHLILuUYimrPleHjOh6V
+X2p34qMmSRKx8ntU1/W2Z55U6NrS0i1/lSnkNCpQ68QT36LBXOUehknlqFNFXhx
EfpAwh9Yr3343+dTigrUpEHetwETkgujlWvjsuwVh03SUvOlSHOs5pI8eT96tcDf
iMseS0sSOdWzcn8fZljlFa7mJuRxPAW6wtqKji5zV/2JvJIYlLhUElFSQ5dk7aPI
NaHPXakZ2HxMrXwfjt1adMnYDiMgEj/eYOsUTbYxOlmTsxyQ7JgHTp8VrupxUkOb
BM5plUCZQrYbYtCwgw5K9g0JE4IxK64dNtmbZVXtExp27E746H6xTDIjQ/3BD6aC
FZPRUAeaYx7wTTl/szN/A/zfBT81kCFKC+874DTyIQVMjhquSfSgc2oaGVkzADbs
QenjmkXGSDxx8ARB2U65IU+XbTM6CwgyLLX2ivyzfS+lxPnZNCJHXTHs5a0qp465
TgDu/+8LrO1VUiiA6SHUr+5rsXFxmucenDGqSJF3T4CobW5JSBzaJMIkC//BCiKz
OSxg7HNbdyPmv9bjokhWdpCDBfqhdn0bCd2wcDr8rMUAySRYww9oxaKwBBy2SSUH
aqE8vKPDsUIxFVOwJkLE3kAxgiiDwEJTq5uTnbgG2rXnutaB4g1doF9efD0vDEG2
g8sbQQa1fRmkPvMXHfS/bSCxm2W8NloSit/d2ZxXRajV4WQc6ba11wEUdR2LHdpy
xRPrjvEue97GLxRYVNVX9BOM0GMQ4Q6IyVF4XZNMw3DJId7Gbsh22oK5SNdO5IYG
bn49N2wLBflU9sqWojRUZgawC1XVKAE9xLbKZ14T8EnLCDNKgnBlDgUdRafjwly6
SucIC0gKqItia62sSDa4m9UIRtPqZN3g9ovPWmSWh6R1QwwdhILKgDdtcvtHB9NZ
1TPY/iy9LCW7kgjRRo+FdiyUopmsswqnXcV9/dZilWE3R0ofru1HSYxQjsl/Mi+z
nbfzsMXFVko7dFMwiOtEpVQZ1FrmuT5XWoyuYDLZeGKLKrVUJjnJAG+vc8mvlwjB
cjWrWnNtuq2cRT5s8M/Co+i6ts/vNohR3EhYRquMx/3e0tvWxpukcrQFsf2Dh1e4
s4L1ZbE2OVIQPF6orEFT3NGil3cBVGTOMf2sBLMdAXrZglFcRnzCtHHRUD9h/Rw1
guPUJrFnMW1MU2saXKSdk0l6V/fJ3eZqEC3SDThWu5ekvElkKQKB5Tkrj7Adkoec
PO0mjW0jyxsWJmkFOaOYmpUxzd35AWcSW89fGW7OvZq0dJlb67t8HY6AigD0rGpb
WsrLqVxx+yrX315p/tuE3q/AY9sjLFiooFdQOIrCvvaw27Qcg0i0mPuntP1/7AQJ
aoPGlrZbZbs5/HhxbmU429fn74IXl0xkU2vrEmD/7jVhgkfRQSFCBclK6RwmDkO0
bDsFP/Xu+E4biQ4Kad/8Dk1vDVuXIF4uS/C+T0122NFm8humaCA7gmBMjjDygeia
LLZXMmZBtZ54tXM4uHoq47YiGIT7588LGMkJqPbn3qsydVqCLnFZXJvwQ+kgWDnU
PyUzb7lnd+sO2YLzuCArWnzQXYqZ3S7S7vpAoXmOOlTgC5CNZuvzHdEoqulSqn7o
CL0zSOLWMFdxzFXzVFXg7wV6WEg09PLjEhRCf29kpgY941x9qOq+Ko7Oo3O8T/K4
DYkW4RpXf0SImT4t9yK54CdsSPS3v/mfZhdxQ4GWP5ncFjdPiU3wBTd0sydW9/KG
n43eJ2GNO/R5eksPeY7sJn0kOanjoB5EW3oU/2DMVVQvNR+Eq5I8Oh1V35Dex2Bb
Ys5fnpsAQ3XXF8fERjLDTypyYCtWBUPXlbz/t1WPMBvsAP5xTSB0SgxLgxhYpp/i
xIglNyNybgTPRlE2Qib3WGurWJSNGHS2HC4hAsNlCZTIAhj4+hvviThgUke8cmZZ
zEEFiwPE4lxzAvc34TlJnGDPTSs2uZRy1a+KqksNkITA9EIAnlFoHKHhmmyp/LyT
yrS/nh+hwb3cAohAGcqfqajYXYQo0mPKJ6tVZIGOpHi0d+6tBXuqVDbfLQG2MysI
pleO3tQXmegb7BxtSxoZjNOY8FD33cpoCpCuR4McqOg3TOVS8zP3+OnM7SGafeRI
vXvZkX1yXQU/FNrGK76c4sjpl8gtB1bcY30cJZJ8OOfdlIAiw0WOmV4/Q75hjj+j
b/F4Yqj2IFwRi6/69jGsa+WN2r7YueZ2gJRDF47ya/zWgntxz95RrHHe9NY5REYc
stIodLyNY9Jjxyey0CwAbvqHFDupcep+o2jHX7PYk4ECFhHyvr+0fGftKTZVBUCJ
+LZfGCHuhu2GyKnhOp4n62MLF5q6fR7isEpVN3266SU0Xsl+pFL1xZuYRN65rNl4
weHbt0uHaQUesh7HSnK6vxt+Vsy9/YPI6iFHnE0R5W6mYftzhSH4U2/EYJSEfUDd
se7lvCE3XeMEKqNybJ7XvxdkbfafzV2E7cXBwrPF6LEDanhpKWMu/XWPeK5Jp1Wm
tSsKcFbvuZL2Xlvus2V/3VgkYneZ6syR7NEWjJAkXdvv1fn9bCPkX2Y6HOcMptps
5cBW1V75uU2IXmu0eW0PHC6m7sFMvzjRb50qaMmjAwJfAPMDWGWBjbXdEXIQi/K2
f6Z7bVZa0Kai6n8woAnIBh7tEFEhbM73u3FUn6qRdGKJGWAoQWb4iBWpYMGSmeYF
J8fnWMlZvix/b3IknW7g0bCmL5r05LqFhMsbE2+gg58ZKzkPKP6dGBe+Cecxfm5O
0pvRTBqr794UOF9FDcUI9CIZa2sxUewHtg0OxUQJWMsU3XncBi6guTajOMfpFNZX
GBdC4c/NPo9dDjEsDSAih2O5leMpG82W3fEoZK3/dV1Y8CuP6boA1Fovh7gxcAVR
7SmoaNU/X+iWzsZurnY3emADYVqdAYrx5e9aZAmtPj2pOkbWZk0S0vc1CICNdCfT
I3WFIQtOFXrB04vMqpVpx4ICrfyiTZxembkd7fQcGlOZzKFC3wXwebRKCj6N1SY/
IH1rJV17stynYefflNEQtvFrjNKmzOZawcgKNhoIBJlkEyVtWHWfr9bv1qPA9JSy
AdYbkO+hIs22i6WCW5WfhZBp6cgo1uIXvIwNsS54d4xrvgwQmYzsy3+E18oHDL7k
ndPE+h7HtMAQrRHDmyojXpxbRq98F/Gad4UvsF6TilQ2mFZ3HXUfBIjA9zh/yzoi
VJtwwtMWtSz/AdHtjgOy/HsAIETmiLY1dml4LCuY0UHTpCte75O5XnVxA1MHK2x1
zJid+okhxuk0sYk+x7fODJtMUgS78v5zecjkZ9gfG3ai1NBgW+5L8DxOwwYu/SJw
VhbIAAijZtIY4wGABSS/DbM2VH++f209sV/XAqKNnTiRGVtw/9DOnLbYdcwaJVv7
jke7sb9WBoM4TwMWbH75XGZTVxz0lQtaEBLo6VVxxIEqDmVm30d1TbbBQ4FtBspL
1nu4Nyp5KJgR3ARvfO5KZBc8SHZQk5SpaSRjVfM1TGzA1nBnK0Yd5AfPtfS4r87I
nc8HR867bp05e9an5H1+EKdIBSbKeS5Ub0Xj1ZIzjRmEK7RDRwpFNlXFJ9SVj13n
JiS5V63s3OFHNxxsPuiccGCJ+Z4utUHAzqYgpqspbEQZXQlangrL7nV9zE0vQwwO
aOnuWLfqjH6bClU7OYGrbL0e79sLUx/yT5y4D4j/55pVDFjAm/pVKaMHgWuRn4BN
IFl8qBK68EPPy8S0uua2As0SoXRVcK/xExNFSkeoHUHWdMQpybQ8yNOo6Txtc0hN
iT9el2ROm80w5qJVX30f+LKx6XSyBnVQZbn1e7AKQsiTnYB3KfbRgECiEixSss11
G55SqLAaV4P+cQuVdmGBa7a5mSMkOj9C8KvlpX85zAFknPSXE4iPjZxaBNka1HuX
1Aya/l/9ud74RUkHnWN94DT7PGAfOzFqDnHSEae67BMbrjMk8YMufevoSsV9Oub/
gATynrV3t3dBOp81XL3OIOGA7MWm8kBAQPN/b5bw3klODMyYlqAdK3GD9KUfA0Z1
v6Itr7yG8XIoJcAeQVzsoMGCHXUANLwKk2rH6hHl5qIEYFYRw7btDlfbnocl/1oo
hjAGjHeTJ9Nt0o7I4XvG++DYEFvzmVxWqMQA6DZFLb+N0qYQjmIh0VGjxoASznOX
cS+firO/cLL9i0nSN//euFyb/rhNATjxfxHhul0dG9bZ0bvIRISfRS38efo+8RJv
vHb3VSqH+cz4FPO/j9DulmIyk04OdOL3Zj/xgyMTVT5tQalKsSuGIO4fNFnZDCaR
ilqcAD7rSHq/x1J+VAE4w1/IFYa/FBa5e0jLfCHl0iMT0m/kL3MrS7cZ727O306S
ihvjfuGfIfHW19P20k+/F/Z2Q8H9uEfvmmJdQ4UxVynzR7Rb3JHyjWBVtUXZWPMB
MIa/FfmpAZqL4AhxtJLam/q8XOIgKTQV9nRzDtIIXwUAWjFeh8vNVnH5lwHtLcfC
8sg4TfB1ghqGDZnEMRBtb9iFihr9eM4X46xdJ8963KNrZXUrtFfnajxPCvGB0UIF
14zskLsuHWGUevJr8p+Y+3KdYFxbk5vfV4UyLH68BMUW0QrNxbobeYXdb9/0tQEJ
RcGnG5syJJXYVqK3VC3W0yvCVa3PJ8DSt3vxQ0/TAwqL2pPJYivY0giTxsa9odwa
ihzdGyoAY7e0SeuAidKip4wHrwWbaKKactq0NwT/nmZtAXWCCu1ReOKUCj5MSjku
3eFKRhG4dbzLd/9XoTOSLSQJZEPgdx3BWbNXpB3oWc5UK69aX8ndrq8mMwusN8P8
wdQ9fpsTInolPdeYolOFSL/FTHCVMn20C4Goi6ejxzTE5D2/PmYblJfdw0WvLyLv
dS+qbs0lXOcR7tAxiPvkOaMFZH8fJV1ZYa6DxE8DrxTJcgwGtLyXOaFXllf+DpZ/
urzLsOk3mlTWUfuwH0gS3t/smG+1zyTLKU4FXbDjCPS2cbwLiq6BBhLpSK+Bx3Sb
yIgE1xTYqZWX6HtYF3l08XqimE6/pVlPFV8mlQd7RIDCdN0G4p//H5pui4uSc3Zg
x0b8xnRCNTRXT1H0+Z5YeWhjOD8buMXJgCAPw5auvA/V4pU2xBVdFD5eeWsS95he
zLnIFzmMIpBftB8HxfP/k2VTvWVft+QwcpqE4+xGYJEXkpD0TS27tYR6BP7N8c+x
nV5i+RNLrumm6KthqdByyRKY4K+gFrllYPEWeTBfRbV5djvLhwF+crqfn1NxrDS+
DvxJP29JPRo6Y7/nBrk2z6isbpgK+649ryFw2P28l4kt+ox8hM2SwQqL1ABhO6ZM
TbbX00eFHXfkiQrp+ryGHcvBi1nOCVWFW44DUbv0lCS9F6ULfRu6EUqFSn2xsTMH
nMVdLK1VZH56WvG2lujmAj2SnoxTABZxT5f8NzNAAkRj04IL3xIQ/sJ2u3vnRbNW
w8nhPe6jveAz/MuSIf8PZItwrkqGgsY2hxyxS9FX+HB6KT9cgvMUmOaPGPlFmhyE
H2NHa3m4lpSu/2MRbSQ9Q1AeakqN3wf7QKM9VFCejGWuc0WT7rBTtJlMskXk6kGC
bIGCOxcORg68djPI0WEqsLm3BMxEJ2SRWUYuD9k0kfHE4L+NNcFeW46LeVi8ZYvm
RUDC7WhM1PDE1nIXqSp2uEsImwvmw+MqOsHKObDa1YQN5Hgvxb6FaTsLbBKHyXX0
vOm86ycIHkDrac2O1VOqz3ruWR7eRMOoHwJhCe8uCadiEuBt3UB/g5baoajNdrAE
8l8Bnd0O6OlO14tYEwqf8sAIPaIC53UQeavMKomMQU7vBW5Ktjrs+XtT8P3Qhsu6
+HKx9PxiBdgEoejdpKDzGlkT+/Y0tMztI9pKfXEg8aXiwLNxPNmz9h5ExpHHaDd4
xN4s/Sgl2sCAIQySJSz5XpPzRekVfqvekLyht0n76cQSrEq6QyeEogDSYdGG65aY
ldKNk1XihjI7W8BQFM7d8Wq4m4ua58XhncErhTNVvaf95VjxXN58QV9sznern11i
Ztc1oIUiMVTs/XH+dyK4IgfG0WACJbwXgujjYz/hCoV6YJK4ih3CVmDAT9xdF8xe
Pl3Dh8I7dEniXCEaAQZ658WXQKPp/tKeICHeOLO8Wj3p44RGlaFwuVHl030bQIjz
RzREvX8L12WZyZnPTu0Gk/eRFgY8ztYLczVaj5b2HKfGgiCKJsxdEgFwTk7y0vGP
8EZB+9Qr6hnoEox7FdwZCXc9QDA1vMsyCHKR6Nzg2+lD9K5gHam6lDjqim1oVtaw
DDuZiuyXieKShoCX9I5fIVy+oyrPS6gpL9MeoRjWnHRiWRWql2H9P4jXM4IrGu29
SxHpAUnAMyiSFc6zRgm3zdKYDpd+bmtBgjqlLpP6okXf9C+rQkE4x2SZpAs3VtQy
sOG+WfI+sqobDTke/kTqOGzcZdb3hM/U4+zrdnsJGs1hMFE1ZCjV9bWaYA6IcpOp
PSoJhLfcoX/mBggj3vb4lKmceQ6NLRC7tI3WO0tiNk/STGaeJosgwTe+eNE9/gEn
o5OgoH0b54j6hwaUaPMTJewWUXb1ZBSdDGhdjjY1934F8tcQM0LEQZqphuSnMB1+
RK0Ie/jr+dcWKJNYha6afQ9t8bmZYGu3GtLcO036uxJD/yjyOQnhiPoV4yIYOlUy
/WfiBxx6vAavoEzL3THB0hsL4sQ6Ue65ZMpRUK3HBtDvotzNhiQjfGFVBLHvMiKQ
hFR1heYrAJfdBb26ZjkopJunyIxdB/xW5R0xCqwZn6URmTpSkkee4OyN5DwXOCbq
9T4GieHPOXZmN4f5MbTYZ546knR1lxL59zWO71ZoQHG9x/PLkjT3+G9zlQy57UkF
qQZQNRYsOyLK+RuKOFnOe7KBXNBG84Ybpo857a7Lug2xpqwK+Z96UxW2r4Q7KDlH
hTezZYOJSXYdNaICXIt27KjPW7cPzDmE4sSJzLUiH9MF1ugmpqmbCyHDWs02OrLn
PQcw/kBnfLcN/0eE6qi4x9LPqCfaATMmgVg5JjT+EZ6av0QynLLBCtkICwbhK7gG
PcX6Obs8G22I2mLpKaZjOiMoOBfepdYannHOfSpr9ucEFJ3uYLPKXHkKqPLfdyqL
UieiwlFKO2hkgOm8vdza2HLVyScTCcCWtZUYFFoZu/caG99yM3qjfpd/HSRKSYgp
UocXXTKFVCpRck4HSmvAQFNpkwSNum2hwOuJzP7JcVF9TCUQBmdI7FyfB/ZlT+iS
ttp2nSSMePzJaTwHVC+fOzogBv2pBX+t0GQhJ0T0oamIVj0bQPgX02vfBlApT9lF
ay9U6+7pSH99P07nWTDMBdmKhtTD+2930K1RPAeNvdSdC8RimEj/0fClO6znNyWZ
Agp2/fLowcbaez0ldZQ2G/vxHXoPIU1pKp6HeFUVQYh7xEe1JUXZCdvuec7GVdSm
do17G42JVZb5NFbnk2iCKobJYwEfnbB3mQbQVaTOJClH1HvVsqel2ATE9INK1EjV
NvOC/xr0zmwMCk0X4/NqcFQbT2sg8KrEJDVQXUj0mA20bhdF8D9YI6pfoiiMfv1j
uME+1moOMeDIXHaZf6sjtOuoRLiayOMtyuqRIwQLXtkdmwV1yu1uBjHFFOP5yWAC
Au85Xua4TvVdUiJBPt56engmV0q7TWuAUaPMkeqPTPfyIkDHlNljfUwgJZNrPo5a
b6+SwSY25MiCKNPj+n/Lt4LTB7Q/H1G/K36y8sdZ4oVezLhBFoHfon+hGRvyT6dV
UUQYDDj6HTSTebWZtKOp/S4TzvsaFCWP20ujB0E4lrgE24MOQI/w4LaQWJLq7rr9
/hSAY01qdwCBWfQU+VdRqfeuGxZQLio0CWsyrZp786TFXmvfDaS/Kt+cSya8XUHk
nEForduAMVjo/8JHE86uDG4jX/rLkUAwH9FzjyrJdHT51DA6ZOvfoPNdiUPFBF1/
ScwWcas8meeXi2Ag0gOwUtL/39Vm+aREosghOgPmZiCy9rGt/s9UR2NXw3Ch0rSW
0E+T4z9v77boXpzoUm76rt7cuRyjkf0+GBclSJivnZ3dlhn68w2C4SecxB0c7E1w
F65mSYagAJqIDPg+AGRE4CR6LYVAVuXsloPq5T8QRSaqpK4L5iI0ZKT7EV/Nplc1
Ucwef8K/EgRGb6q1QqMhxGYyzQt0k3Pa2cXnO2RwaedPY48aNCueHemg9aogy243
0jHP0WvodQx9mZ9CSQ0IU4Rw74OnT4xVVrceuzz8TTqTa7SdAJUIgTXXpaTdEP5/
MlIGizP5wtYNBu+Z7Fc+xVk8v9lEZYvTIyb9iR2BtRsJGuuksWIrXtRhRl/aKTZ7
x5yELOdXkXoxPHJzLPLvVc1mOK4NmPX1qvtwtBo8T7ly3rS4NFtzAhdD5Xde2IVT
UTgvZTU/GBzcVif3bYXXdgckOQptZJaMu3b2unwPZ7mJ3bv6GJQwae4RgfNd+YAI
/8xSF/DbIsQpdq2Q9Em6BEwcErLEmPIkLUyRO6efaCvsuj5DNEpC48MIavZCsbow
pmW/HZ9GSTh17SKeposjgs6tK/8edqEFsGE+KDFVx6RwDbf+3TlRwJ20L0X4c2RH
kfrxxPgm64Di+/esqRXi9NZZU6w78JD1oCuUhOoRFgRIcWkvPpxiPZ+oC5Q3eO9h
ESCZi6Q/QRIXpm9A7l40bAb7p0SvIaAi5wGEryFIYu1vLprJND9sISXe/+gy29ar
CT8HvwZPwtHOe8tyO/dZKoDt2RkRqq5dGL99nqKAM+5gQxnDEcUQ1QOheQ8/jW7M
B3bPRzcYBfy8vBDQUUVYu4kXWp0SZiySegT+94sS95oIh8vo6DfrRtwMOOQKR5CI
o+RCKcarPIy18TSKP5Kb+aJNQOGoimq2zqjdfezbRFYdrBzzQjkp5u8RmTMScHy9
CedP2vP2vKDk7OsMbazqFTC3H8kXM3hCwSm9JpRO2UWVNeCCaYPQLdyGo3/pOCSY
+X1P8xymlYTMKKEg/8aX9/TgO19Y6a0WWuVKlwMrkML8FTrKGtSjfoeMiTpQAENX
Egs8FHotBUmvgEghhS/bwFcLw2+TK9jJovN2eyXBp3QsE5wKd2BdNMu9iz49qWk4
vU5KngvN7E6ipHJyeEoQkYTMP1+aW6k6coEfFc64sdJog5PqE2fKGsRGQtGjDHVg
07d5jJhIL79WooNXoBmOvxMiig+1RaznZnsm+/wr8OMI0UXGEBCkE0liEfOqN+Qd
8JyWQnvEGbv3aYz81/TtolUsxFHZ39xcqhYrOYYOdhDPZwOYo/U+XEHilDb1hQ7e
if6ZjSWWcixH8Tv3M4L/mDb3ZMdIWnkax46YKevERoOoGqSvHxRu8GSPle08PjKJ
wHK9SIpIIGLvwsKgOl6FHRvCvNTRLNXtxqBgQdS2KDoKFF+SYbIazbr47vNJwsHj
2c1jRIkO5tggRSWUszo67wOKsmZXZA3l6PV3jkfTwIgYPTcfrFS684UlJwAOBsKB
dSX6FZAum7zjmRXd9k1UfEhnXinGR8NZAgiMDgmZicsjOPiFFpsnxFsoSg7gLYN3
Sw01d7E8N29OJiVcyTUiruG+Z0OwxkfoWUYgbHxMjAxMmlSlhIRoA0mSm074l5We
xsopS9yoYGG/S2bkUQsEHgcYqr77MaQAFEJkeBuRIhjkMgH6rxpL/bqYI8RpCzzt
3LqywHloZ8AZ8+bMXHzZ0dE7chER8YR2cTw+IiiJMtH9AQ6d2axnMuqjmy2OG5zL
YRH+FVnPRtLVojofn6jlSJfDO85IRV9swdfOQQX7KHh7Int8eelRgGhT2cLpIZhM
RAc0ABIvi8hPNGgMfucLxICJbfivYZY58oq0+5R6c+3xJ36hKwLqziNz8fimirIN
gyK6yC9slGfdhSyfgcC4+zW9FcdQ2eHI5mqm75sHwxJdRB5roSGSDrlUw9jWRr2H
O9Sm+SwfN9g8F8oe1XYGh4hr9iqd11c9LBTrXJIZ+nVHVXKtfSkbLTLzTIZdd2Ww
3HOThTQu9MS8e04nknIk3jH+u2Vt3CAc6/N3Ya98C52D45TV3qjWiq5eBJ/yWjSD
bbwXUsBj+gMmQc80UaNGt3+KAl5IVYxJTtR7h5nfaloywqk8DlMcN1mCO3LsSaol
NKPrBHZaU9yDD6FMwHIeR4ItsXaRF3oEawKE43vWVyMvoxc17M8c441oHwEyWWKA
7OdTTb+pU+c2eA5gwrFen6VwKbq+CNo7Atp81Xc0VjfT5bV4aM/nsoFJ1vxKcjeH
RPGQSWWZ16hrrG5yKax1Qb4YDPa0bkm2aDyf3G9hgIDKgNA0R/uj42UYWCOzq3yu
MDfTxhBieHaIUTgbTH9VI4tEcMhcMux5rDRFmP4Pu2BgQDvXgku2eG94QSL4hdvF
r3q/OGPRLJ+2+H2jPDju7rPnqXISELQRCrJZFzkrC2wpfnyNB5D5z+f63+Tl15H/
ssYhwHC8GCJKTuwIB6pe8ky44Psn5xhLQ7bl7586hvqco52SaqW/vuud2eow7zyr
26wOYTy+pGnFdsE5lLikoQW159khX0xDL5Zp7d/7aASdrN35GICgBL0vZtswzH36
Ake9vAD1sKAVfrNkkI8k1bUQqflghkMvE2sfcnH/D6YDYvQs5jkzQHE67dOOlKEC
GRmrD67FOJGinyiRHTgT+DiIIEgALThhMc3h75zj2EWQ8MDgPE7QXjqQsccBtdI8
jp5cVtUZceHTJy5U1m8SiSEGiXM0/FoMEu8cueoArVypoDXzQRxGpD8q/tpfJlcV
Cy4fFvak1tD4n4UuK9LQ1vbUcTB3uWNEJDxECW2tSuD15oYWBEznnqj1dmrQJaHX
I4wpOYO9YrXTpVJ6ZB2QoE4QddBICcZWIZtHtb37k6cUEHOJ8NT+pW+me5ZD5m4y
AUzBGW3Jm09sGIcDYDxmZjTqMqpWzXoP6aldHzjtGGJ9W58l+VTOh+krLbFdSg/F
6fpi4wLMofr5Jo9vr4z0mUksGLHodqycugDedZdsxcuaOIyq/6ibMza1FEY86F+k
Gr8j6vSrk4YRQWVII0j6kAroLrD5sFhDpwZk/eW5k6npawJcA0V9hv5jZh/71DIA
vhbh6Aby5KzT56z7pcieBb6r3fsJuTTTXgRQSkmyUMjqMnvcb4eNZdUjKTxDIKwe
E/fHviSD/Elei8rNB1BEj/wC/OUo96INRJK1jDAGqsZd//xeqJuOdi9ZP/cayp1K
9szvoSiV0rv0YJgmo1N2d8S5Aup/I85IHJ/C7j6FX73BHRtVUiaFVgXLcitEqknQ
zjsajoFIEef4EYSGgolEFIcWUnAlFz6z5zv/W3Y/l9iGWPSZaJRcyvk+PJ9lV2iY
WyHa33V/jqY8HKsZ9hthxw504Dm9myXdAdC67Ar9igeBH6wyvIjAwn0fslZs4yeI
h/sqB1kwL3YIPq3zcdgAyEOya+Z4zm8A0FCIGsAIT6tCWm1rZHlKNc3CbOlwEAGP
gljbxyuwodakYO/6x+RzoS3Zd6LgSZkDMiIzDkrOeA1vcr0m475CWjQi5cinW3/T
uxZ5HEi2Op+H5kurEEUluJN/CJtnTBT0A9+j5x7GrkgmIx8al4a8cFjqXiSbzZyE
H20Vu8UjL0hIWX6mkNoTd9EAMwU/dnPhiiKLmhkv2pRZfjQL8U2qUjfU2gS+y3Qa
dcOe+c9zO8L9TZ6ioBAKtWECYaq/fjRfVAR7mOh3ld0juFblM8uEClbnxv4edSzV
qn3sQScKPsXjXIqk5hzFdVQvHMKnRHALDaRast5KFhkguCd2/eW7bnO7nHCc8Gxa
0LFbQ8k9oPWroRRESpWEWxjqrZUdhfUN5i4Za/VtAGArWFIo51XPfzA3FeNIOWnT
ANPlo2xkceglQ1dEKin8N7tmhA2PsGPLh7HdOgzTboFJHOaLlHdiESjazxJ+Pura
fyn1/AyCJIHgI6ZpH+ipJR4kn7sA6hsepSlI2U5bHMZbdMNpnTC736EvgMY4/RkJ
59Tf+5Nx0D6aN1bVBAqHQuqb9nv6HUA4jOQY3rIWCsF9coQN2i8DcFOVY9i9JMM0
4MjCFUShfPqE/iVAV2znj8yAJmpsQPFGNM6ogItn8+veB3SyM9kmR4dcTcJotA3M
tKgTl5I7396ndTvIo/eR84ocp22IYUAaAwNIICIaZHhfUhnXUo2n9zsNQjCz3VuK
rIhU2rtWLUsHPkidFRGbSgYr9gu8+6NoVWLDulnEwU8qnD1UJlv6Xf75myLZW4hg
zG0nF1AOR3dYgMtn9PyXTaM7s7ysfe0uCoLv6LsF4sArAtYg3Uw+i6cKCBpy7GcD
PDxvzky+wKZr60qZBWl7RQANhNFDiCenxtwcl3jzSUxtpTcNaGP/a+vZ4ueENbS6
WOSFTJOIq/4q/DWiBJIAL/s+4FKrBfWXAJvboc9onp81YJR0929AQc/4JnhnHby0
fO4gxjq0MKIw9bSqhnhp8pknd7/Z3jbnhA6MmoFhJSUoJhQ8N2koRQkP/hVk8Fmt
8sskBW7qp5TDAydKVejVCCixYTsXcloA2wEHNJIvyBr2Ct8WPnoLZ5yhIOOpV44X
5EDGLxygV9TfX04odUSDh13AHKQ9u+8ZX0Er3YQ+DD+iUvd9XSFBWBgbpPxJejEp
QDrAon+zWp6O4jolAKOHwcrMdyOghr7wQX5GhRfa2Kj/TIBhRDzQQg14ylAKhLqE
tKFyId4JcK8bdv0YdjABz3PfdmY3EA2fe0biMzZHrTzB35lpiCCoZr6YXS9h6n7m
r+O0u0M4uBp0v55i/zswyO+yqaEc8448vfSEW2t/CARZ2CPlxNgig0NbztA/gA/m
VAWKj0gHiK9UpnQvjZra1HMh2HcydCV5nq3Bjwz13v2zwtYvIwv5rIbT4/54M2Aw
3ePu/6VmnGdMybdwQbFefESreXun9RyY7x089c18u7wkyREsm5M/7f08u27CkIYJ
+Xd3Qhd2tn2/iKIbXYseo+jP5A7DW+WWQ/PBXjduh/2/u47hvxA616/KF5g1ldzq
mjddl0h+q0p5PxrUzZmMUei/5hnHANTVqx3FZyFnyDYACGV8VY6ais26sCDteZkp
O8ULKEiltsZvSdZWEdsaKHcpK3ZCCEZq+XnKpxv9nlpNocVr7HPK2p9XqHRrE7QR
JSAsMGlFMcDJQKqgJNOI2FWumgpfffdOOgT17RlOcY9pb7TzeTtPQCSa/PQWHZsP
sffmBkQ4/PWmcIkye9GS8hjxpS8Tu22VC8+2ZlsvTKnUx/4agUJEwevjT74suibB
kFn6aL6wdj74/LHwloBb6SLSEgWUTXUJ/Nh9RAJ9r5/5llclXjHUIs/DTj+ONHrS
3bFNmvskJSj3+hb5N15iDu/17AkybLjRK3oNTSMthG5hDhr0pCvgDyjc2OxkFAyb
m+WASVnes18eJfYQYn1W6Sgq7+NOiK2dldS//H3kWSBbDKs6jd/s+tLzywTTSGjk
q87yWKMQ2TLmUHFTdb4mT2s3tE7+qOnflU3g2tBhextLC5gPD8QDFaeSFY7nQnep
2UvCZYsfzoxHFR4zzpGhKUzZSSKejVwUkGFNBF/pRAFxZI9GwjzMVXbOmZOQVHco
ThuWv6tYpo3VjoxrttUYL9xwWxxIjav3B6e28rDZHRovm4t1YLB05L0vGxjVNgQf
uC/BofAGkRtir6pEKeellmJ0dD3oAj2LJmYLeuYfi3aLvHhyleebApDx+z8I/uCL
38xOdhUt2ed9+rsFsQT7NY5fjMx/JWBOl2yCIWJAowwH3qw/u0HpB2EN73AMJoC5
6NeeSqOEmNdohr3Bxm5Z9kIRD6pNFXdReLdLcTttE1nzRtRcCvRnuGG0k1v/En1k
Pdy5HvqUPGA8KmInFrmZSLnX9RiQvhJh02qLVs+NcVtUTK1i3UCoplnfw2QlqZXe
tRhQKozORMP+viUqmh0kxpS7mOqwWsdXMjwBH3AlMPIOwosAUAR/w0o1cnpJp0LB
Q/3VIGkvs1h1imSfd35r469S1YIXhwbdnyvfq+cZqn7v1RpQxRdxMS6NmFODkDOe
wk7Lyy5/3aDpmzNGMeJFLbrSsefzyoyrv6mDcyxlg4Kpip+HBWdHKZnydM8TLGSw
zkfj6szgAGzJQ9lY5Exs6mvt3ViY/TJIhgcLlJIpZFpzmZkpf8f/wo0ZHQBT2JwY
dZBCm9ZXCCZylLIcg1pAg9+KP3l74KZPbUSGwMljrZQsVepZQxrPm9/ztpfdPGM7
u58HBa6qhV5NpVNXLC3cWNPQy7leKdDT/TemL3YsT3RO3zEZxgMekoxzW10kUx5M
wERzYo3BLhC6u6FtlnPbNHd+/dsJZyo1u2jf9u3/ymedKDrk1UBgkH0L+4zZJz1r
SpokYiMLn7UnoBqn9L8Bphbs3iDTsKmd0lU1bDh3f1J2hPW7z27IZN67rR1qGVBk
5tFtMa1Vz1lN8XmPWlaXu5guwO3bx9DFJOzgzTPlZy2xnRj01GLhDzi5zCabrnWb
KDM80as3Id5LLJ0sp5lmSD2VqaN2ewJMEKphsRJH95+xLKyrkHtL3C2YcoHNBDr9
c5oqFS7T2z2KA/G/xfDmIT8J5ynG9xgBd5rMMdsTBlHPTxlC0Znu4ZZ+adUDYcAl
AlmzPYKrVk+7EF/pFW358uXj3kbjsvhVAOWY+qcBdE+H2Kcj7ppITJ5XyjW2EsQw
7Pv9pBxEIAhv05fE8ZmDySJXA2AjNJyC0oIdtcmHSzESeWq6/JDI4lgK+6oIcndL
06F289+SC8phbvUZpCJ0V1U83n0MLDlutAXUCdwSB2DSCxU+l3ksYSf8fpeVuo83
XQHR3U+BDlhEk6hbVoeIGEdxTU8l4Vr3bq/8rN2xyfq8ZC+zXE6SMUEyrjEYo+zt
5XQxOZVW/D6oEmGING/G+gdjDyOKKfOZ0LkSUrd6HjmcFaDM8Ez8vOEBb437OLx8
Rn+mrCCOprPLMgmgIrgp3SguTUB0YVihn0QvKGWkirSoVfseBekn0pq2D3JLbE5y
2Nc8zNhygfqdf5Oa9UzGskbp85fCRmkeg+ua6iMJ5qDopL/AQZOfAbvnuGyz/K8S
KySsumnUIdgrUkH9qyF19jq0MLSBw/CZMHMNfosLGxWQxBwziwuRU/kYutzevYtX
ovrwZDIXh4DlnKcHAIy+dEBi2OOgLXZSM/gKy8qdNdL1wgCMCEhYWUVrfcDu9Nln
VtaNJCRTgCv1klBbG1awlB7WyJeBM3Or7tpeLAhw8lpYt+ZoGDMCeTQ6SC6x4wPD
gzi20kxcRbzYBoyLPGq08dzjtBH7tfKNbEEwm2SS0ZB2kbMo6QTCW/FTkYYuTg06
DRTLLkGgVtCk1l7Zv0IEJzpNfXXs6iizlC4sN0P4og/PIOPu9L0SX5QiNe7oolO5
gOKOmkaJgjzC3rrrLXBlTbUOErhTJYFSidJ0hnV7qJ3q/6qoy32VLbOGzB+ZJx7t
ojzsQP13Il3Gzh1jX9jjA5eWePYAdNGcNCA7LogIStXiO4QqW1X3YvxsvaduBsVq
e5r1XDA7JRIswsCfrUZErN7JS6vGuYuVjoKInPVR/p6QAM1qsGQoPStMmxcxXuqK
LkXIWISwF+TXKvcLdchJeOOIWgf1F6FrL5nY6iKM9FUji0pNL+VORSimaAgi3PXG
yatOcMFiet3BZjGIpDGx1/ACF/8zHzPE3jugLBORB2ibtArA4WU2xNGTtWQPWmHu
y+WNj7uml5x2gRz1CmxqSsCQA2pvlzEnT67tqJQQ1/1A6HLrDxHBfjkZc70FHAew
Koc4Bc2G1viHtmNan0QxvQdhC3AtNkZeQzT9DTjbKYDp0Y/h0fjm9TK0VwWEbJU5
EyGwkkMXp5bTR3b6Tyh9GvcN8KaPouf36k0r0EeCapJtQc4ebyZUe+b1J26FB6rE
sd4/+gnE5Xo9IO060KGm0ou22X5C2QeLBFqsujeXU2Jl/WVhfj4M6XTN3UbkmJe8
tNxa96RD49ilXY2m1EAG0v/GftltzCNDfzYALez+civZPvmrOu9DSYxC14yqV8GW
G0ihSjze67bjfQ2ghX9ywSeC+sFCgrjQfDErk90mrI8Tjxkuhml1tmvIgzrJIH9M
Wv0ZMJ8FbIazowe4BLpM/cyB9MuZ7lvBJyfj1G6CMSk016s3DEBxoA4Zt9p7y244
I3H/Q29jrrAJHQVVVBkvnlMY9XhuvQSPG7ivd2EtRzo/CjmgCjIEGy2M6/248nOb
M0J1QnPeG2KtqbyOWr17x4oYqyYd9l4rxLo4kIwv4n+dNnf6jo4lQ0KLSNWdrEwV
REBELSnJuFVG+4M6MMVhL3PX1e1gLv1/Rp76ySITPDKzLtYEUCMF+soSZo4Ow2VC
04PFi2ixWqug+UWbfa74dFW3jXrh6910V1+TOOkrA9jliwOCkJuOzU6P4eCxjetn
vXWismH/SN7k2I/yuEJoSJUOSzWJVQMXNKSzO/ObD/0fJDAv9puV5PU4jGEiZ9nJ
VaVXW8QtNP78Et5athY+jtZgFJAJHq4aPEervwcINRc3qjwr035DHYo5M6lCww3c
xWcd6VPLHJzLciG7o1v0mNa47rXKv6wP4naAdmjm8gOOi86F6BNoGnwMqtNcCFwS
pXc19qf1UvyyLzfGbWbBN3s0NkAW5jHzZ/JqYy6xfbsAjc2Df3oZlXpOYxt4Yt7N
GiSdVOAPNovLJg2TEeudPH9wOptMywNWIO7J+9MBtxTpc4Nrs+Yu6vH2q1MTLx1i
iAqYm3GWLnBBf9PNRUTxhtZRdmf/zhhmDDOg2OAGyPNC08BLl85IlYsFtU8akt23
lOg1X0Sb3BMvKMAbY7adHEa+6yowaUXQVkDW7VupNCHJcaxMKaveI39BT+fUJ3Ya
AP+9roaN36cKCVpfZEJciIgUy4bNIrlIgkAPgvAy981n4KSXhOvTdj1hxkzmsKmG
7PAYrcdRqOORY7zUXi94CRplQ2TLJR2ICPlS2fZLeFHpI47qoMGAX433BkLYK4rR
guJweOW8xUGV9EPWpaN1fnODvn531L7MrO+z1d01wEGxw0rwkbLf+Uwe3bp5AcWQ
kditO37L+sX48koEktoxUotVl3mggAjMMaaHXKPebSQSdDyh95IaLjohD1vhKII/
TgWTDTteNAcU7olLwtdvIxB0kBLgl+j7s46yPI49rYU2Iys2TZQ4G7yJuqghnXzO
ElXIvBmF95LEt257oZRJbqZMrQs58D/yMdqCWWO4Duim/OEdbOkjAPU9z1AIHHfp
Y4q9jPWCFq+y+/RnAPOxx1pK6ZpoxmBuwgUxh7KI2AQNWKd5kjhc/kgNjT9HlQGX
MPHmlO1IFSzYWKCWyUEYgpvhW/msmI4IgM0iKGnleRlXjJbOFtwWTmteUsGO6Emj
dmr2quWing19hMphQFhPPEHM/0vDPrAiuflgcvkCT2WtsUNtSjbA56fNJ4NEgXHH
I69GWhcK/1CfLp90kB8t2pF9IMxLapZPSt2fqXaXNhLb8LfgJ5bW9VCVTPtp5zrc
hIe2oXof9K/vR390/wGgEjvOuybxEmDSgM86uo1uk/u+xHbomrD8L5+pL76wbFBq
W8PpwCUsJ8ecaxtahN3QEtUmTf8YXUMryhRxom4eVrMka1XZnYaQKAlxmCglsQb9
7288IKUCQyATWBujwhvJOe7TdVWORNlsxd/6NPwRlYElAhYEIOU2HOkthxfEQr07
AnbGAUqHJy9dZ5VK+CG7r7uz4GJ7EA8TWeoSTupTy0gzehAbF3hcYYiQYz22hZyK
0i5TdqOxUyZysAEK23VjxjvC32I7j9T8JwYA9O/mUuzanv4e9ZigaYb2+Ck8Jqrj
0Y52jkQDLUCy0N3sAe7q9Al4hQBPAtZFlugDe9Mbsw/Uua0c5vAFdEV6GtSS9hmE
KN31pFsZON/HGKZF2dOQlvLWNlIieW511/e5JI4OJt77AaLHMImwSIpJVViAxOq4
KiaPDesyFeppi9kqZdYDZRoft7N1RjsjgcQHHDZ6WgSrRV76OuxGUgC+zNVPh8ck
pzG2sa1CCxNQSxqNyGrgvcSEmvqll2VwOYXAfIeMr9o5kgIQjTiNrt8W5r/A1n/v
SpTG3HE59sydQ4zI8nzjjGtQIc66cwGD9LhLt2DAOo++hUdiPCmNm4LXgD0/bFJQ
R1mx4s+9LX0X+6UvITuCnemsaigsYV+SrLX/vZuKIeDsgh99k18y5CvTKDlBcZvg
ggdJDCiYBFX/AAm45aOHa5bgZ+Tr/aPxbg6KC20WdBm47JDL96TBzNLUJAhL23Ss
l1IXY55Yl02OMLpsNkTaT++mSa4fSw8rUu8C4AaKeObdpiO4zCHvfE7m8maZTEEe
vuJUj3M4ziHRfZswj3nfkinLY7NVKzAj3DpwkaRNf3Q6VwSAvIuxrSTaJsoFM+FN
S+FVNu3ZQQBMJl8A5gKfs5nDb6d+u4jeI5oyte3Zj4zWFQw3nUOjtBnca0EuswyR
u4XMFfxaNoeILA9HjKLxFfjkBhwLSdkgQXPquxBV6lRNAVs/e7xdVewveyKQko9n
kzpLXwZYIV5Wgr/bWtBmUcdTOUjH5y4chu55GuXELlda8POLNPO0r7aBiWUBlnbi
7UUWwFOh6IiMiInufI+I1azJVtXB8udC+5gp/HQLYnweCB0RwQdB2Ve8kQbYX0lS
Pw3X+vK5wLdkmp12xCBnuGucQXppEPbpYHwJdZQwf50XiA64dvRCkVpen2k4B6qB
TX2wLFteNUm+FQWjdpS8SCKqi5WQQN/uC/IqMxtsV6OKkO9BgiUosiVoPDYyx/35
SXcMkp9K+lkUVhazHLSraZao7KqLArbYEg+4SNDX1F7lxmEuov9bo9HaqDQAco+A
R7M/ljg5+GnCgT8M6fq5xWdPBkbWsPI1Tlpyqtbr567GiFF1ITbFK7avqNEcqxxF
nffKHiMFKA8TZfDa5sAXAGaJowOEAuaI9ZpmdPyR04kvgzxkqtiw9ylAvG5QXa3J
nBm5hKZPE28Se4JaziI7e49VWccnlVVbxaxSkMAYf8oJtka0TM5OF+cltsSNL4Ph
RZTdmcva24G7P8NmoRvZl8tw5AGA4hBlGw+u/E0Pb8atr2KkwLYhXxoHi9BhyD61
GSuhhnLF5R5v6Z+7zCa/Xs9Sutt+VJ59vGlnL89Ih/DJWFGoUHBiCmqOqIIn/zxH
fXKfBFknhiODuuPZHOS2fs1TMUmO5uFDaHc5lXRNR9Hz27v+3YiCHKMzMtUyhzWQ
V0PqpC+30mfZ5MhsUbJAv7+FG0qFHxbXhErU83nUYOcBqMHqaNiYDdXdPhorQxd3
AYbuNBmGaCgYpeX2pNKYVuqWuZqkPStsTsMVHLDS++M9iDZZiN5NThOq6a7Qfsc1
oIrWDhqgt6q4I+c13clHlne2OyvQq65YgMK5bqoFN0njLQyjcPDidauzY2rNQuNS
4WjzumoEDc+3S42sr39frQAGVriYnbst5/8jZLBo/abVKaVxLnCak2/1vBJgEOmY
fZTImPuCFUEhjOw927lSNp7VzFP1Ctqx7eyh1IGkv0r1uOHbwN2700zWm1sGncAn
K3EHuaK0PykCdW0w9/ffdXCmZt4JW2+mOq6WICdjrrDK98ZS+OIjwdhMhJgbHRHQ
u8BDXOceKy4NRZgqB130NjSyF9jsoHmwAu+NSbxK9LKVoB+MHa9gse/zZZykFG9R
qVjZvp3tz2bvuEhv6jYGBDnLMc/HO+gTTRdg97p1wcZcCYhuegRhJ/16okoL/dcy
Xq/GPiRv7/KiiCVNOEEbFMuabUKst2vSCBhD+5fTGIRPBpJ/RUD2lnWdG8OGTXaW
LY+hMOPycOJeYnmLTOaX6tQIgpQQFOS2vzYNggv0V5rv3h1eNlW5mzMV+rboXrnb
14tx2I5LJHmTidWERuhFx1geJTPAwMuuFi6A/yrYMqZEHzopyX4u58SSH+uzNOvf
Vf/yJ+An6uK9DJ193k2FDD66r/i+i67H0fFhxZng2Z1c7Hir+b6EH/VYNVxxfVt3
K9wPbmBVXP1UjdFrJrQi5ch2V0IiJKzD5yueMKXQwS0IeDKV19HDSP1C1xXfKUsF
1YxsYA9ghv01Q3tjAvzjZpvMh0MCqTuZl2IGCcloeOvSfxg2ymRVDGEvdQnlyrgO
OEGASikv86A9b2eCl6kxC1tTaA4HHRm4RkxUDoG9LLl6JSx5CYIHm7x48lIuGRyI
+1JtbJQ2q4JohUalf23v4GWwx0Rk4Oz0Szm1NSYU/PuYW2RmflAJEx41zENa7PAb
ITDGS+H5hMcI9/sNgqQAXRU43kwbQzjtQqDXfn1FCYHBq7cQjZNFK3u3g8/e306M
daTJuuf1iNP5dhylnZCFcW9h8yVriPdTGFrejAj33xumB9SIkSp7+Vst7n9yaF+t
HsMeQ1nnTMOJHSDxx6UNWGTROG2gAdoEMDHctZAjGSYfZ9t4VNlKBu/dL1KxxUCB
HS7yua+93tUS1o8gIHM2yk5c1JqNVbfBOP4fSYb9yM8vKVD/+ckn+RfTdwjktoC8
6gJRHuMhgMSmbihLKC6ZHRfjQ+zOLr96RgADm5M/mGD7ZzJJor50KGsx2sxts/Mn
HuDH0S1Tsim2N/fYYn/KSO9K999aF8uCugooMbBjHpuTjboCpClRFkv/ruj4h1Jg
cXylcwFZuLmWn9Gi6iPkvmA96e8B5kMeKT+ZigD4fZrXhiXcBybKHEU+s8aqrfj6
Xc4cYluBOphUh+OgFsTaDsi0xNOmk6ARZmKVREAjiB79vTmll9PCyCbBuoG3qihA
WTr7FC/3JtAvPZq0bWnkDOwP3ScEvkFHc8Up3CnJYu1d2DJgso7lmBqh+f7Dmqg6
2oKcqL56uA3enw7ZkfGj9rizJfpGb2m6yxkRsen2kcasOoQIczfTF6tGuUWCzqGg
jicRuF6VkyvUTAOSLhrIk/uRV2WChBZ1LIFYDrdeO15LCQXlsvO7iZI6ZqvhA4Sb
OVWLBDCmeHOli0ZWOK812Wh7iNOvNSzrHrqPJEiYGzVZqHMkVoiSZlAA03X9gD51
lY7F3qxzWf+eM4EHSZE/EX51edT8+mP2pp62ZSf7VSQ/s5TQ6aal7+luZXLNZl58
9O7wmPM4XZtP9U0u3QV75XAue1oiA71sqHxMfsTvjHlCdPYCTf+HDzKpx33x8xop
IxAnciiVvoNhDcOumDCJSshSq3NWjnTyke2FWiIiKAP7H9t5vR22KgeL4Ez7z1Pb
R5NRJKVmj1dadxak4+Pw0rxVfYV10rL+K6YkLjDLDqnvPfUYsRiHBbmfpjI4lJDY
Yp04uJP4sbNDKExigYhssgPFJct0T2DmcUUKSdjn7ayBh9nW7AbpKGPGOe18uSXr
kIw0PwzE6Kalwddl9Pby9i8i+r0WnbJyzX+LqOA0pNNM7Nbq1EE76wjC2oxLuCrL
p2XRxOg6cwUYN34lZaGxnzl3aHQJPfeCniK79R9MIq9VBiLZmvRC05mJh07teMCS
XgGpnB59PI/KQkWGHY/KYs9Ny44UrDFMzJ5Qvqr5wWtODmUoJOmvxePWPezKN1ZM
buJTH6F073Ed3d8oQPneehYeKUodWCbP8EtFKuHi/TDpxWe5kg0eL9j9m4+0mVw4
vTU10YIPX3W+IOCKvZSvwCCfgoZthWzxnY8+GNXSv+1+dBjUG7FRbCrJfGPqsSIe
NE7jW6yRtrZ4LD29QNCnT7+UysOZLGESUmcIu/sur43frAj2lP+OohteRKco/pUW
bTsNM4viVlzP6ko0bdV2RfISBsfkldMBn6/6GHidckD/m5/7tXm0h6fYvg2ZjG+r
JhUY9VT10fLkAHANPslzMR//CQ2H93PZWaQcq4DLa6EmSfW1hmt2UKs3zq0BBDH7
v2UyHmfVkZd5OmiRUxEQPfDZihgk60cSSiEhUGuSMIzkJN13bo4z3n+5HUdY8gXS
/GylgP1wQbzcH2nD32TGo90hLFoF7wYz0JgAYPjnqCiA+YUPkyNe1x/Qm6dDkp6f
0cuLLQl8SgrKftuR0g7sKGvJ4a2K7A/lPqRLABJWYxznWP5WP2A3fSbq24F+7EwS
SvelW98srCRuVwbJJV2LqtFMqPOoZ9e14yM4BAailyvAvtRIRxhbaNXEUTy5vrMc
pvwmfJ6CntYDqob0e2Fsyi6c8KBmmyoBZpQVair7+OXPwRd143vct5ybXYUvo4/o
cj3nmqrd5Z9+aYzSSRDQlUZf0uahbJT5Qr7ueWb9k2nkMMMIAS359nN4qa29geCV
z/F07d9AIc7i+pRGyQxJ+RSwE88I3XID+gco9jUZZaxhGZVA2/uNjB3b5BKRKszw
M91/XIBPDeLjX+pHBNTqSPN/++rR4NrhXT4/gI9hTVZexwbgH8P+CxU17UBt37+Z
8cnP5IOorwyIZPJiZttpJlOQ16P+iaFtjVzvdUWMJ7KpnzoX87cf3kXit4hT0+To
YYkcL1v4aH6zTYBwwywVIFNRNbTplmB3jJrfJbh4PePL+BjW9Vb3K10wPHlIDmbr
IxKZZUsEylosrgJP5/HxZgHgwHjDGq/B1JxyuNIifhsaQXjBuJDytdR7som74vG0
NO0KlqCNHg7up6MR26gjuPrGm9w4cnpqTxjwHb9S6iHLqUdpRXZgwD5NFWhdmJMW
VZojDVyTt4e+ki9hj2jzXHZ0UDD4/s2QrPsgUEVjXhd2+c7W0KtoAL4prk57A68W
3+JsyixTXijBRbiT3avh72W24puQKFlq3fME7+Mk6l97c01JIXrIsOiKbePN8jJq
yTshqP9kKvvqUKyBhRUOx/lZXaJaBp3lDeXhco0R5wofxFG26eYmRkm3m6ZZJDtn
496cXVZYPgLgtw/ACTrysu6fEMu8BRff4CiKEXwmsX49mICxln5qTJiFhtP4Ktia
O4ioFfFrJwD2jddtn6LZ2WcGnQJ2jjCD8iD9q1g+r677dtR10PAkmYKdFRyiVC8N
3uU/g39UIpR4R2S/q9DPyesO+RJZ8B7Q/m2NTE9ROIXZg9DeMVMyNJmJvhqkeuOJ
p4FSTxJufvqf9wRNAsVxFqZbw1eILRMXOljJLy0wm6MRN3APHPYLH9urd9dJLOV+
Vq6c3DeRn+3dqblP7xIUNL13kRNgf7bwW8nc1HkS4CKAkIpEqRMC3jnqDNEMtHPU
ocDix61rxP1W1KlfRBRXFlY+ZBHN3Nip/rtv+iWdwGh6fjeJShvxgBPuErZGHQgJ
Ci4ioYH5+b/2bYUgAjq/9yciUO10EIuKe7JflQ1/N2zzpFs/7HJW3URNuygN36UZ
sPK/e3dpOcd+OOmnn+kqMTkf1Fts2bUEKzDPNbLZBvaZZ6FE0nANs4QAh6J1Ov7q
YF0aYLZ0GSCFFFAhrUU0uhR6NEmd1g0nPjg6f+5cgy5TmgIlmdjcS74jF3Ly0a9f
9rzhEZJaDar0xLzQT6b36fk1ywJg68Xocbfwr0VCHGs+lV2/jA1CMJqL5JcyMb0t
cmq2PAvt1Zq4te/ee90I9r8Z1Kezkl/XS4q+QNZ3nr44ieZkcw8Lk8PimHePI0ET
sUZOZABfkgba2zd553WWIVYZkv8iaLB5EO0HNZaD5q5P83ib30V/aZ6xOmq6Z5Hu
0SFTDv3lpZUmk2/TYSOhwA7mUJrnyqPPkDIDE2Phn+J6alKcqgNgUIT3OHRco1Lg
5R3QiOwc2Y6CdhwdSz7+zQBbUGKPlr3obwp0PcaQ8jCMz3wi1kREPXBIYmdwzmzU
qp2Gcg5WZ10Yjk2sJpV5QxqmUI8nVus/vuS4wEPYiKDvJBSIrzI0YahyVv3jnFBg
vhOQAOrV1QNcEuF6mlog4XJdrIIGp8wrEkLNZX6gr8hEvUkvi02ACY5X6wHa4zJ/
ZrP9k7HLTqzIe0hbYnos8/WAfm1J8U8YDE/nIARJerHSZjU/EkTfTOePF/DF7wFq
mutOJ/s8JAywiJ7K7pnq5RXIBIgTfW4RG6UgWEwObo+I3bf0kOXGpsahCQH5605m
W6/Tien/nlrCCkYOhFTuH/cwKXAJRNk4/MdrZ6yNi4/KwB5WrvHy5OCnVE7BjX/F
kt++ZgYrey/cYPI3QhOqz1LWE52JQFU8uWprxrKyYusTNE6gLyzwd7ftvylDyrFV
kam7ngnF13wgpccnWW4RmCMCX0KKcQT/82LkVz3WgPy9t6SQIk1P5Ec+uURWlBqV
K22K1Zec9XsvfuN/x4Tw1Kp+UF2Q3xjae7zJ9uOgj7UtTqGVL3h3QByjOEXLYGN3
fV284nEPnqYcwjWV7qfXUMRHb0kTJsF4fcebG1GiKJui0tJIV2iE5U7HDyezyu4p
jP0hcPL4BWKMBYFF5f3oXanOnaQfFAkZmfpgXLAC5cq5DqWG1VVcgSKgOvUl2jOR
kkz2II9tFAS+cJs8icXjbpumo9/5zePkYyzpVrk+y8nq9hfXpYt/YexTq26bx8y6
12n3L9XCeTbAExsUChDQkLXnp1rd8iy1uUCTpD/+FBNV60Ixv66RVwpgTOlxOxC4
Ngw8ZpxdWv05P8bZOoxsDbQjhgQYyhhhHW9WPhRJy8KapCjpKIoRcBO42+s85VG3
QvN9sYNgmuy69nrswEj+7G2MZgg666ZjXR5F0I2WktkZDH5qjzAn1J6ACon5OHTJ
WHHc0r9Vs12YGU4BHSkUgXMKFHIuohTP9upsOQJnVD9KHi7SnA/sU9vnhi7Kjzst
swhTZgJJbhCPdQqiHcFpljoXGiO9qhZT+y3LBamXUU/yxmx1BOyA4lCdb4I2hg15
YDVaoHOHT2jNO7piYz+K0ioIZJ3jMM+fpvOQbXeKC/NqFDMX90zTUqKnE4MhoMXv
eRs0cOI+JKQNFjA7vhAxTclphIEv7S7oIcn15ME1oV0kUSQOOzC//2dQDpa8NFw9
Ct5I1HQfiBObpE08mAvCf6tkT/624ODN4KFwhZr2qdFRpqTDXSXlUAiLrEWIlWn1
NERyXRVgX8gCp3ifT45oI/jDY4e6dMBRYuCFp8LAVKjmfOdBZ839aGYlzeDcthrl
eFXMh59+X+aHOdr0PP0SY2JmINTnw+nqQRZKbOFX0ZOD20yLYuH9jhjpPyPta9KP
2dXbZlVb6M+2ZS4Q/bKdK0fLnMK6UV1z7wMd1OaZGXH+h3cmtu4tEJagoeiGFrmm
f9WYxxuXl7dCz3J52ySdn1gR2dnQn8w5lRWtJSDXIjk4/k9w8BuS8WvX8EZhTBvY
k6zqs5xrRCX7se0V+PptBBLuKvWQcobkyOsNnQb0S9cMh181pBtPc++gor2p2W1D
1oEMSlJNKg5SGUKs4E3JYyRp8EWNqyfohp4YTGONjaD/kVkeS5tNOJdeJ/9Ylx3z
r8/+W5CxuUvNqKXR3xymY0PvU323Ua+X5sFNu2xEpJ+uFUFTJb9ufQ2tRJQO9p0x
JNGkjj9K/1LWHzE7ZKyGPiGecIkNienOw/vLO2qQ7/47DJ5kRynM9HrPZFsoatV1
0aEsISs5uZU7GXuZyWC3tSW44vGMK3JNvCReqoD3Nn+msXc+Z3zB9rvDpdFsbhcs
P2MIdU2mA9mQeFuAf4Y/HIheCQudbnjabGYGZZEaFvdf8YwcDYzHD7umz/x0MBEl
6waSgsi8RPi9csGHcSNFj5AiCp4R6tsqTb+D3NE0s3JIZH+b8NFhttbvwfuuUlPg
lj3qflgsLmtcwu8vCh7QR4PUpKeWnzg57qBmsMpzWp949TggjsBPdSzXpRG57o3z
p+JKCOFIh3+T4eohFGXiqKZXB+PZCuWFLY0eDHhithG+W8nG2L20t6PxMCeo9EBx
TPvf3H4UGoCxHXh8xtiX5aUebIgbk/h/u+e5lbsz1qmiGd/KsBmBjSurJL3Wxdeg
FD5/blWz31SGzbGbZ0hPDqUPx2YL2CS1/P6JZl8XaBEKCUtSlPyVW6/mk4DkLU96
fFHvGRPTESqcs2c7rMCMjJYOlbK7+uUZHIDxur4FvzgXzW2Ghdhdn9IPFiwyqcN8
nI/hHiCzPhlPHFUclv2kSgSyrHgLdxhh24f4XEUJ7fbSThduxPD4GcVoUbsQhLWl
kQmDS0v6DDZehkDJIfyH7xc5Eyc5awbeCPuea1J+b97amPoqFM5UyVJ4ULSSotEe
ZoKuNeOWoApSNfl67ma2+/jTPSjHhRtbCqRZygfRTGLsIAp7GiM/oOxHRm1bSEst
e84n8xtTQUtAuj5sQHewi5P8yqkeIuogKXkJBmLilOdhY7UFqRFX2uJbKYiBFIEb
DLmb5CF0wLdhnzDWyXKYrg/0m9h87pIIif0W4tgG5+MNV8tRaTeyx98eldCifF+C
6bgTqg9/Eqbze3StlowUUcMOZngSAxeIJ0tq0AR/6x2EUslxcHNm2tIk2lgmBS9p
1Bv3N7zz/MPPtD/28JNLpjsNv2tJz86bZPGMvCkcXGW0Jjtl1OiTXlJR5bKa+ZLD
wKQMUe34UHR9ymFzNMhSRYkNeieOq6Ix4CQ0XiXzaDSm1eDQOVpSO1qFnOmCZv5Y
zh0ByRr4CRO5iHIKFqQ1fFyU1ll32XdT2pBcnkoG3fr91ubvhAxuhiju0S8MiwKm
gZYYDbOdbCisHrvEP3r3GeihQgZj8BFVUEo7T94whI9eJaNoDUxbQVEK6Tj46iT7
26r/g68gula73v2zby7C8MpNWRefzhkug71PGxIzwOyGMzP5JPC8vquGzBaddK7Q
8b686KHfNPXYf6sWWPw9qsfcglvAj7LuXcP+U+DQLIyFLvQIRxXG1kGqhSvFH1OG
bnBrc6YLZ4ITiXIC2hRLMRL00wx5rq+XfO590RemRkqLhcLKGTHhslT9d13HuHCO
FATIDAJWR0kVsrj0AjOnV6HVG1AkRUSIJXqSbuwAsQ1IqOlNdUFrAGKxVc4TjdGc
k37JyNkT0lNlJKXmsBTRucx90bIs/d1+RzikxxH2KawRW6kJgFbu4js/WcY74OSs
VBoxNEzkReV5TTTB8jmew8ox/z++Nf31EGKZbvrPDXf9rdVDbsBvjkKzmh2H6QXA
XXdK65o+NS4XnK/NYlwsoZ5MAYrwWsHcDlCJnzS2iOeMj1JlpB7TOe0pkJn8mFU3
uU9PGhK1c2gcudPrfraCwZjXX7uSeEZSYHb1S90fkBslZ+zJ99clAPo1HuAnJjGx
OhC25DnZKEmhl+sQmH4N2QedKlJmy0/QdgHfuhB/S7t6pBRfpgR+DsL074yjH0ky
nmsRh2X/qAOLGpEOuFfnPp2Z4COD5kbCKaqaLgTGap7PM4Xu/eH7LoqJ8ZJWp0H6
PWVT82D7b6YfZ8w5lMyv4OAWnP57trk891Tbq0RHDEl+amrql0gXSIObYXgvxb3r
ATl/pkBlIbjQAOEkOAmSrmLc9UhnG/T9KU+O/QgCCjG3wmLAXVHAOUTQB0SPwF6u
PZ0Nu+DK73HIhxt3IidIyjvU4MfKfLC7Ix+NptMWJJavqBFmkekzZuvhDTjzxF8r
Dw6cysf/192QUl26gidBgTXwJYMdSnqQsPQqAYuSmm6GfvZ8kcVC7FTPHtGW6gVu
h14WScGa2rKfBpkXq0KbiFMPWBWW6H8NViq7rr+tcxq7irbLAE/F6DqmlyKv9/oa
NE0ItwOAg3eNdlzAP8kqfApBx0+aWHCTtkjtws/PhCGlTIExW58gzA+tzewrYuVH
f322HG047US7KzlOpNRzm4UyGGj6iLG9qF0yjZYbqEV4hMYCXOJbSCd44RtnWurq
GK8dG1uMnaxgvnefJq4CF+/+GvNBriKF8Jy/jCMxI/g23sxJKbxStEneCVbAOny4
qTbNE1i2c8xHf7fFEeFlm+X/tnCI6aHZF8eJGTJwsWHMoIUWpXHPSaM+GNk4rSLL
dcxv033Xw2yrs659fgKwrSY/6z+yfn7SgWc9qL42v29RGfMFuqiQB3LSNwVHeC21
1y8IGt4GvbtKQIOlmKgsVbL5BzqXJ2zkWDshPki07FzI6O8aRjioJLWp60nDxgjl
STiHXm5lY4PFo8eL77Ht+F8c88Ad7JYi2GeGseLoEMYLY0AmmuR6aiNXeOCE8XGL
LEeHLIiaQcRUfL05Q2/sW8tq3vI90Hx5ZliQn5sxoz5BBcWCQLKfSviRKb9zbkWa
H6XsamLVXTaIQSL6ZlC2RxuxcphKNf9UKg1A0/9WLVTEfXE/LARIjVsJDUT1KaRk
gPWLYcowfqv+8DSHOlkoaQzrUNjp4QSF2M20FyrTQwVUNmhFIf/aiJbVOW5UqzKB
xTz7hNgnbtPP2jB1z5lgVjzNAi5Uyfe+iAeyrV6i6hB6N8w25DfLaqycbJMangzx
32hVj1tHspkC0lkdC4LyKqWZ0kcMMU4+5QhcghC86ukvccqnlBkPM+vZLi03dPnH
cmsPYZNaacETqUrm+wiMkWESUsn4DqHH2nnCZsYXnOU4wxgWoIbVzaKnPhwry/Qr
sxaDqUhgQglywGiyqy+pGP/KmpVdx2y9/nMMWFhxBm0HQXgpp4HM+gGcjdz/PRoU
sFPUvagDja/r/i6QYarY1LeFod78lo3k43KqWaowiISTBLPK6NfFHqM7vTbVfwav
rugdManu3r1jIKNFGBbemc6VGJSde3DxJllvin4rOLVzigH3Iozh8245Nk920BNj
WVabqLx6o9eRLYcNp1+WR62QdFOIKsFqLEqeZe53Yk9CnySYJUPNwsaa/l/6Q8n6
F9Kax/UrstO7Rafr6pCzxAb5ADXVOHj9jdRnVxIWqUIa6Ii00PM+rn58oWMTpFZ8
Gsa7qKSU9ZVICJ4vGajYOs4ycSlkd4Jqb5IFB9g8RyPnHA05yw1zcs5qfTL1aT47
nRQFKhIQszEMWwvAGvowq5Yi5NayZg3u+WN6AgaQugvKSmuSFHRZnrtdlkkOxyqo
uAS7phy6E/EppAtmFcYW5wouaFRCFGfFT65iocJSZ9ZjMt/6YlO65lkp8cYjpNMD
Y5RrgOf67sb/OZRKBFo1EsezLqKdQBZ6OXFBIYbXK9f7uzLKjd0MTbNZT7Gex17A
PZtmbvurNaNUa7SgwX5R33ffyMTzMP3ssbarjrG1zfwc3s43ifCiekMAQ8yXnvxM
UBYaoDsRpm5WtT0002rpyt/+UDy1cWP+MWYarT6iCBABc1NnrOa1etIjAitMToE9
3QXVOHf2EWnQRtDThYT2B4SNq1kjTJPBM7/nG261vALLKMjfRHed+9s6e/fy+DxV
TB1dHbq4y6fAZh671J6njdjJKyrAVtes3QIz0x9bLIOUtPQDDMuo1Lkxy+LDViHe
ccBIR5FlQLhp+fvbdBT4jqEzTe0o8HkTeWHTEI9jytgIzgDkYnB+ZzgWKzdVDUOk
MatdOWliP1iAKNP3ZHbhmYt+j8YQEftH/Q6K28TWDW5bUXrj2YfEpkP/5WZ6opC0
yUGtp4qDl+Glew/DdDeztiX2C8jaO0e8y0t5A5wttcqpQe0YXVdVWnt+AhvJgoj+
t7z98sk/KoB932oLqu3vf3QlINaFHPzwGlceRBrrta56dRm7W+NJiPwKrlu3ApQx
WORHh+4E7Dc3zQb6OX+4CV49tpOQOOB/NfZibahJZLSSp7Hf+OTEwxkk8g5RTbfS
X3MTSG+OSUyx9mIipIJ/C/UfmKWJc4MP5NhN6qQCmcIihaq8EsnD1vxHmCppSvtm
j0TP6/dE3BpGhaDk59vIafCQgtJNjdp9RApeaATz8AhmCepNO9c+Er6B4YFcuJ2Q
+TCxJ/QIftmXc1qC/bEhEGj5s349xf/TClAvifYPk8JsdlsZ6xClLjqaJnp0W1nv
3DhElZs5OP7YnwGXA4vZasZ4h/6dW8uUlLcCxzQcW7r6j/lbk7QbQka3z3zQMmng
zzzoaF7I/Jw+khSFBtW2MwGe6XA3dIntuYMSP+koCRUi9EEhM6IPd3+FAuLALYmB
4rzyialB4eZ6cJbxvCfGS7kyMHZDwRuImWLmzNCqbhoqxQjVOKVBsAo8SS/phqoL
ujmF08/5G/kbfRgOZQLjfI+4QhkEDf1+R2uMhvbbb8n6M5It9ZuY7vgop0Z3HBvD
qopjhcEMqcQ3tt7eus4JpCfhWzp4ZRptrKCUxl+uy43cby0F1WczS53U35qhQe/2
bMXocGCzuo/LsYgSb4ljqGcMFA72MToictxb3PNLgte9iu4gF6PzSzMdkJhfMYqa
Lnz9XKAZHbMSDJ/E9H0ZgUSmm8b5fDoAUfWojRHuaRUq0Kr3YLrcfjd4lkF50PBR
QgLqiCla6hWxW8oIJoEBwuIK1e8wKsjwTVoutRPQMGkdK/0T/Ai234H8i0fEODDf
fZOckfFtZXqYQU+d4H5LU7wq8yWtX8eFsc5xpb+qXRoPOKw2zd3DyxppYYetJZiE
khZVjW6bIysEgzGVi72jxWGLQYYRWZhWVZ8mIO0Qn04+cF/sQGypkoepdj6HVGEU
+RiwtfNT9Ho3OfBYbxJ/aZsvGeSLckuG4CNbIp6arFHyPx05pJprr5N2R3izg5kV
27PzifSDZNdQexlglCmWamcxMmJCIWKMk/wdI5Haoomoo9itWpe/AwQf9QLPneHK
XPRNzT/SR/mJ4LmAlUksxqv5vJ3VWrYkejbUhdC6eLkbJg4+OooDy5I/LhyeNwFY
Mswm2osUYjWCdC5kzpYXmK2TGiDVLT6UKSJPME9HIqgxAjhYfts2BmP1c38dJ/Bg
LtNVq9+SpciNiiIbmRDLZbEO1V96LBzmD16I4NVgEYU3ArpyWV4gKzs7FMJP/r+L
gRisIfwRf/xZ8/Wfh0/TLSWO3aHRuhpbaLVtN/zA9ts7jEzHEx3Rc/8HuuUyDk4B
4xv+WrxnkLsHybhWIg0B0pZg3hV39IlqaDhB6Baq/OPXuF7ZvniODDplb9sEnndu
+5i78u/6Y/LYP2iUshTARVPHifZqRoAS6+Uv4PNT07R+H59vEN419cpQ+XsAt/0O
g+K7NH9wGvzEsiU80bRpIewOcfI7d3ZloDLlQmpMvgjcMy+VB8mskdPQVzn9PZ0V
smnf/7d2fWARl3q4Txtvjk748rl9MIrHn4PaSeT5p1Bt+icfcYeUuTpBL8oJU4/4
qkSRAXy9CQy6vKVhv5uahG8+stI77YAiwQYTs8ksKWPqq2s2KJcGi0f37yVPp2Jx
7BeoVK4ZyR/+UoIXlaOY4Sgl3LFdUPlc0jftALHt3GJpKxjJeaznIefnO+wkADpQ
Lac6bLnHVdatXLAIsjzaV2HX/oPG1+Dr1NH822wWF4wYALViLw9pWfYYKGvj/w92
cYYqNWF/voZPj4j51sjrH08cxGTTekBTzED71dvnaNigl4LjrDjGXTaajLqauwSX
0aLX+AA08c6BE0Mf51g0yqGbXgBCVWKUuOpNs/HQa685vLy9ZtCbAFWcbGukbQhq
uCLrVUMYOAbUt9Q+ztX1LDTEFlDmXhSy9VJngd03bm1aWu5NX0ndS7SfREcEyMiG
+DRG8Jj7FuQ5elnQhV72J0//g4wOQub+mtKSGP0TpcniBMYIS6GyJGHOlsT8otvX
wt7RjcU/p3bkvKSWMY1HVMdZSqTOwFU+ofuZPMA8BeXTQxmLJrd4jnzmv7UqrbtB
6jy4IXmVwPgE3/GOKbhP1lFRppdLjHatAcqL3OftTFHbdwCK+BAUPNzzJ/8uTalG
tVMmDEQeQRQbXzdm8wQf5xu7YzmZpn31w7Bkk/CAZp+bvfEVlontGQEWwxWTJtRQ
rqPvoyNevdFsww6VlHY9+5DThSWNiIA8EHLizfJ3vR7dQU0lyr56tFuNHjSJ7PJY
oBsErBM9H2eFx4SJDnhCIt34Am3widzflpAlrvzthSI4O11HeS1L2E/7Vg2rjjEs
Y8NsHtPF9qyOqPmBNrgddbXb3sKP5o/+hKvvG0eLb9LjG6BIRUxUmHIHGkCdjAGm
p8tDsrPNbGUFJSmUCIGX4Z3481dc+vzaR6id6BcFfgdNQ206nl6Djqj3tDX3/eLZ
aHOdwfNDcDtep7X2leDHgMBM0DrOPq4PoANNjhaQP9IX4zLSuIkzgiGgzdemiMlB
IFJHrQ7R9gd5lpnPdqKUvaS6onskhtiT3S3VBWYrBa4u/Am+89/2o4uDUnH7L4xh
ki3ZeiQ266m3mHJIyJ8zEmr1cjnAzwqUtYeP/94Jt8YIcbttN6WkfL8USyw8sh9Y
bDNfkFTIg/TbKauZ/z5C0xkHl02kO4RyCVM6MgXweojr6DR4mTc0sTxpTIRdN7vf
+6+T9/v0fss2IncRpXvAjoU/DpSy5M19NVQpGeq05zxfI4s2BZkMPLTxgo5I7ufh
qKgStKU8yPEjZcxpJlCily8giJ4oNtmUajagUf4To2ZB1cfIpNh6VoowjhwQdGvC
CZIszpcDIfXNOw3WhD8HYnrKeaBlkqiv4NtJc+Yb7ZLaYobzFZmohrD1CNvtjgt6
/E+/e9DI+UihyNzefFKl275lmuW7i5UjTCwOtH4j6+oBEc8YZ3Z1njAx2SVjCFn+
aZa168RyrqyvXjcSspDKqPN+cxETnxObLwHdBrMoKOFBRus07NGwcbRvvlorjmhG
M7AyKLEuempGMRBE3WVrRv51TZVI1KNPuVv6GGSVBC4qEB58VuUjY5gkeuwW0QEM
a+3ooxDd0LQEW7dwvSYThie/965z65AtBm/zKXBrau5wDuNaNcIof6jn+nx6Tu4j
xn+xdvLONLB30too2ZHo8IA1Q5YPRn96Ewneb8MpkywHPLfRImYrwSdEpGYwKYhM
WZprtSTWgXYH+TQXz28NBVNbB260iaf10T14YDOcR63hjtBVAjltT/hB2sbvVEfa
0gkW+qJUl0/hYW9Zx8WbBVtycjzaRLKyDwE4IjNBmUaHQ3v9F9P9BJt1tE1sP77d
3HRJ6owwhezd3+jsvrD6fUdNTjNXnFl01Yj6lvgQ/IM+1yf1RF+XQIOmJjW9h8SF
ya6O+bnqYkn4O48g7qa3VJ52yA6jq0E7uNbU6Ux/YvZBeNlapFF05Bx9s/K+KHnJ
ZIpk1fEC3ZiTzoMFI3kQYeULV+BY7Na5679kX0SmL71he6lHqrTVPHzOcyz7z9/L
ZZR3GLYo74Ct035zjdYCMgUdGc4JiQKk+Rba6YWAnBO4q/DDBWXRr5EMwopUYJWC
d/Y8UKQgP1XyZ8CtY2kseXc3QZqGCHDmdpZ/3R3yc+SRLvn0TSdi+ehosrc70gIo
8pAO3/mSuE5s1Awua+0uScHUR5wBeDeos3sDRcgmwKEDWLvqcilRqrX8iCv/SyGJ
hNdGi46nTR0q8BG8mtVN4f5oWPTD4Eyfnkk1tgbGpoX7DBzY47thC0fOdwvZpwIE
jdpaIdfgH4rkW9XZRZqlVupiNuu1IefaOGfGpKp34re5i/ql7tjVZ1VYo0l656Hd
3AGj8plocOkiMx73BI3vwO5sLCJ0mEcU05RcS9rxjwkAuZbxZJ/PB3LWsis2Q4Fl
Mff6h1kZgw8VIJLMZ9JgPi73gdOd7JfM2n6RafQ3s/G1apFZV4ZZQSa9S+ASoz4E
H/x+6A70KAjDpHiSmjMxspeHFUgzN5sQShuI1dlLlHadK3R6zfsv2EY2i3ojSWYl
PneNq/fAp/bg5ERU0F/kzOLNDia9mDoVtMeqoC3IMoMld2n1opJCuqPPh+faBcHh
KnJ1/sWYW67tNlcYi95IH3tC5wPVEPfSqW5MTanL+7GNmqeTt5XW3p9VykRUk01v
a3QmrbCORWlL373GwP5UYIWXX2oUa3a6e41vi2UGkt4e1YkHfeOGxoi2uvg5idRG
Tm2SIn0bNaBf0NR5WdQNGWfl9qNuPUDPKfBGYGypNyGzapobVEijF5qjVc4vFEf9
p4w8zjmNmaRTIsdxc2xMNHsgltsK7WPmZB+tdlg1j+i++UhcYDFuVFFmDWPJiyWV
b0IUMAffZJ1iJKu3Mkh+2auvhb5JWMIB54H0Nt4S+UHakQnFVF4PjFLi5Az46CFN
qCDe8MZi90Lu/Y5HaDAxrnhpkz/3+SPA0SO6w7OOcPa5BOltiKl88Gd9RcuNmwH0
/XX831AunTA6OxWBPlvIa64aNsY/L5x2GA9aZTxuRQUC6z92w97l1+bJ/80gVAiW
FQEfg5cn6cw1alPzncEqOKkmFHIdgsW742v/oJWWMq+k+T5yX/eAwDWJMtUXzLI2
/cGech8lQVcVj6VRlB6GWVFzv4abua7/UCMHqrMI1nS6rN1kAK8HEp8d5/2vtJRO
TbvZcqQpGtnTbWt1eyaiSezM4dm1s36LqsZjFqVyg6WcXRorLWVhOPLTJjYnuNcE
ZPd0ATF66VwdX12WQzptQYaFKBl32zo5x6UgukI2l8pC4Mvp+i6nHCbruE664lcG
2jfVByO16DkYPsuNnOhzDQg1GNMjAm6dZo+FgT6IILazL52jVehRP2nvYvJrSbtv
0SmEptuI08VYlRLRnVA1lTtKCzdEOaPXJCrzuiWrw4knT11gkBBqv54yH5sKRzK9
Lo8BuDiUrXcxt4gZdMyePCvGs3hFe7C+5NO0X9IENZynw5sDJygM8sopEqbQ26hj
wqapcBWF71JMbyrYZszgm/rgIoutHkdVqRr/Y5jQcu6SFJqo1iU2dDVKaEw/nS/p
TcWVCnx23DrzATCPWsF8oErA7EgUETGMJGiXWRbAtyAKB+Eyj0G/LC5LqPgw0LWT
yAbCjyfx8DLzF1a39YQfAw1KunhK1IInB9v/qsIJ69BNkKMvHrZYrABS8VLOxWk8
s9FeqHK6EyBWwA5XGU9aFbNkASwVKIqko1nWYgZSNWIzDBloMPy47WppGfs7mHkK
VmH0Xg9N+/bOVIjphdvsDohZjDI+y4+x91fPd6zjHkKzS+HjS1eHf1+FThsFvwJl
hm+e1BWP+TQ6OtkwhgDFufeqnUX1WWHn/n5DAySWhzHQfs7D4p4GTNBEZQ69f5xM
l417TwT91jlRigF5aLCJlTkufOh8Mclo8gq0tPemwclZKuIC8bkyVJyCLN99uYQ5
uJ4iQu8sBcFEaMrwrlPv4dunxJdFlToEzMoB+UGYDE2YxhrbCvhnL84A/OvpxW/3
Ck8I9h7rN0Y722rrmvX3R1zpdttOi/+4US815RQFoagcvQgYwvrpY/eDoARvrqhM
7VTQPuGIaaAMS1EykKJZQFltyOdeq/u9okk/Ei+h3bCvMnhsHyfBpTWjTT53V3ZS
BvPuH6/UrDuyJCGyt/Td8DtUnL12bcf87St2RpGw0rSdrH/zk0Oiws3dTp/diEnH
VNQWisUcbPAtTt5PYN3Wl9T2QailGQek+Vo4Gg4JYBHwhv8OmVHz6LcJ2elzBDR1
b11kc9WwoiIuxzcpgBB14jFXa0+I8rJpc8fTTtfhFgAGr7JoT8ownWbuhRv7wCH5
CQ9bX3bdxvm/EtCEQ0lt9q2axptkcEZUwwmfiIMXairPW4lxOPfv6fACubjhA13g
SPK2qe73Gfvk7N8Lhz09BPl7j3Y3xpU3m71QmDPUYf2g16N5GK2lE8T/f8xZ9xJQ
p34kC0Z7vNnWo6K0/XVKFN4e+FSTeaKMftob0pkUtO7RcKQnQZ0+RvKxpA0m86Ja
lbjBB0hLRoc8RRQWRe/yRIuFWBIUjsNjbxrSSjUBMzzqWpcZO5DRcksjj/L5DxHi
uGsYDNFPWPnrlk9byPrFWDFTl6NxOAL0S05QVka4I7lnIbDRkLWsJjQ0PEbs8tFG
kAYDYcgFbImO9jL6cmDI8lrA7jBJ8Q3G5l4hHUXq8N5WYFM7LjKfdOJ+KnFubykV
rjCsif83LrGQ/FyXT7SIrbH9v5VAIggUNUVg3pcrOrNfvcaaR3fmEfKC1NbAa8T9
W+0HuXW8mZ42Ay2/NixSICmOVxsXOYjQLNb4cs7fmSSkZv2+QR/myfIkPe1OIAuK
BqIVHUVTONKaWHvWp4z1zdnOcP9x0LlTIjrBOAB5aeuA2Iv0xg3nlBCyHoNSGHiH
QMuCW9vJhPIOOWcyEW1hNHMnHAkYFCjQje/8MVn+DMOg/eeku7FJM7J79uItQStU
g+Q1Yl5RBjdrKaKUqbNz1IBMq2OLZT6ZXTpwzI15j6CDPOloTFYHpbWGlmGWaQ9U
lBfxivAwzlZfMUyC9fcCzxOHVkT13IpCeI06BYa1Cl6VT24IGVx6AqQ2imGOvHQQ
iygSGLetLmSCC+odUwKhg6SjnpjtkWknYJKjVWoibBxpVBHofq9VpiBizS58Fxij
3PoJvpcvmeQWvEMT0ltWOELODAvK9XZWwxEEsepgkj/3jh2TUcVQdtQg8QHi2D0X
4nrhFJNnosUMUVyC+wUwvrCQjLUTuIAdvtVzRdz3z0pyj3FbUopmKISekhEuk8Zt
Ms7crkIJA0JHu1cSADQNNAORrmMy7zJ++374SCIWm4yJPJVWtpYflvUr20a8cpRf
VUz4tFI7Mv9V3ksdr70APN4NFNNIHhJaovvOraj99xKskaiPr+/6cfuXDVtDa47N
snLiUmihzqkgwTpgbhoWLnl1GQha1ZMDc8TSrU9BUqsZpfv0nrQIXEifGLxzfPy6
YnOFOga1/psObVVoPRGfNiELQRyhwMviTebLvkc9ItjJIg4x1VHqdTxIcF/SkiW4
+cYPApSxkBjFBn+SsDVnR/OVxOLZFtAD2PXZN9lDiBmB4JUCLTA5PZTpRaS6WmyO
w85NqNsNC2tqeVywzo4Fi5oTnBzE6AGgs+FA3eL1C95ayoeQiVmBaLNTOtv5hqkx
S0948k062dD5rSm/d2AD8sBsZHSuzlnfQLWBumHwQarxQDiuHzI2HpaQMHdrRKqD
dVPnVaFIgpHfPNIY8bN9WnaqPLGyBt2jzmB2rXduBsRUKO5Uz4XN43uEMzO0R++I
wcoUfl4vhr+wh3aWAiA4SzI+UlwOr9iE6etk2VAGA9jTvUZQCELYvODlVh6AISms
J/20pPipI5QarOTtceCWLPrKhaOikNQAjDWSBYLTl4N0HZdDHv0izjrMkBQFR2Fs
rIHlh6sZbljOmWSZTvapDKL2FCc+CMGtvjhc5JEnUJ/y2mfsH8QlDeE3fN/7+N4q
Uzv7NIGKw7gMmtlJtqnKt0XeTbzX0+m/Z0lxOSX7sHxdrzF1f3ipwu7hEpQG1AaG
zfFW7uVmwPe51V5ZPkK9Gjgp56BYsUGwuU91/d0eQE3QtI/kpq4KQtUGLp3MbLQn
ZgbbRw3RoPApAUyPEfe53LdIjPIMLMdELvZlNwI/MuuUuZHm4VwJEMhj1x6aK+X9
OjyXxf4N5BThYAStB+mlkiOJq2w1BF1XfqtQ38Zrt+M9JaeFlGTdxGjMmHc2xTmZ
BtHuM9rK0VITJK+/c8U+XsSBgMHAHALQtWyHR9IJOjkb2FmE1EkAYKTKF+IBW4vh
PlXA81BUiAhZ0Pbbnp5Sbz1KpziGcJiuBbHPUxleZjRoPvFQ/rsITvseHp+HNb0S
0pGqCSroK5jm8gSFJylvpRo1t7Avy3lEK4FvfuuErzX69itH+7TZxUS8D0SHKbQ7
fbGnQZL1ld7W0pCUe9Q+MEPnTZpC6sRQIsa1YhiB3KJcc5srrYVv8INkAqcc57zR
yZtVHPAkUZrqsFvpvMifp/hLqHmJt6Dg6U95oc5NZQNKUVm2771fc+U7A5UZhThl
/ZI5pPNoOWNxc8UK4/RhEv8eNE6fe5URJm5zDrI6fvnQhJQ7D7Fgmpkhx7FMLqFz
e+i6UbZB75kdifcNyy1XwlQZeRvy09kyW+gRpMfXfuOoP0SoN8VB7SiXC+cuk/a/
d2LAGIEELT69EBjZMufKzxunSz6HGpi7XW1+JdMu+488yMrVYNo8c8aCStku0hpS
GFMz0bNTmV1jLsqlfnpMFZNfYoHAKZcfaL7eo/Vdq7GVGZVOSeKFP16FJNjWkInH
C4Gvn/VaIVMzG8jtgtQtckb2BQuwTMk9mxl6eR6uI4hFnnSAahoo35OHAMMgtWQE
piHJvIHlvtE+fClch/2X7iRyJnErF9E750CBlFT/cvV8d688FXdT/Sl6EFDWQiOO
5PZUYKBo78HyPK7Ttcr9BKtQW85gMOyrxYrP9wOQNwRDqZqqcHNMbjfwFh6zkrqO
UYOqAf+0vBROvMPkkfrNGnk34e0UgZ/wzj0p+513pn1Pu6iuq0II+cX9VRtuw5VI
4zBdU2UrND0Ts434vmcMRsrfL3j+kkNDa5y7CumzgcpcY3qH2CJfo4IP7dT01qno
EMhVJWIOjBBxmKvnLTSu/mvbb0vkeP9DxRE1vH2Nbd7StPeef0jyyJAL24TYoj08
elsCT1AXSHkG+2a+8WoqnY9j/mod8Ya/fWFj9nwbQp16vIujhltKC2ZLtBMr6JfA
fXtxf+PioJ1EMRwuPtcxwVPWdqMIGzPSHXx9XldiVDhzYT0zHwPF7kc3Ku8f6hsN
AZvWt9DAWLN/dHcdqJcFxdODNWAQecia6XTTfZimmCKHF+Ux0fVrbXscMWxTn13K
oK5zEbaiXG/6UAv4iJfOgzUNmia3xpEID+jV+5nA8SqgoO9o6k6ZMGKlnm9vjVNL
ucx2+hueD8L0jIdLJXXunq8vjpHExoIispi3Xv8hnSdDrXD3416kGCOK39GJyNWE
0GazFkops3yW4of6PKhgvC4zPkt63Zxq6LPzGru027imVaj7Ha5q+FuqtFhzW4H3
qXMN4G77tlSlOMO/YNEDTnNhR65BDclg2DEb7d94SFqjUqNKkUV+mxSKCJ/906ak
H28bZeWE9LXJgNV7X1fmVVaFLnntkoTi5Q/HBID2CG0UrTsABCCL+JPrnSSJQ0c9
XLaY0rCQpFxpqgUMZgJYa0zkbTPx4b4LzzUTnYH9OrDeSQRzEBt/1/HJvZeY5KKF
fWIBS+PFvwK8oqwDvxJc2K5y4hRyMVGjzKflOPfiaerA6+PtqfRI7Q0tBwqN5ITw
PmkLR6huLmR3eKVhyBBfTwhtDy6LpYtlpcRPST53yhHkalrJ2uSGPNSttCdcMGOS
YCgdgho2AfMFJwjsh5kdduGEnc0mGsnLovETALp/NT2Pfy0OgSUdL/kQVMVC6eE9
Lu2xeCDRztQ9ersIGHhLIfRmb3PEM11NiU8vuFRdHAKzGlWkrcv1jynwZZz/xFWG
Fm9udAXipQapJaMBtimJ8Ta8h+m5yJdagmzUyfAOGGa/9tOdcvbxVhK2CyW0rYT0
IT4BZpW2V8he4kf+cHLk+YuPGB1vXWd6FQc4Pp9uxdKcroDE7GvR+VnjDW85KCn5
zvKFApbwpsVgaxv/wr0Px1Yg20ousg3diQBpur5PZGsr3Cq63ibjxtztZcjDFMl5
iZvQBBCgCW5VfIa3S1aNwlOuL2jxs5O0fvAYX6NPkNUlJRwN21yKVB09O/E9ai5Y
7rb9gNL8jsUdZk32+4LhuCUPG6k7MmY3YpJUKAXbOUYfEHDKr7pdx8+ftYA9l8+x
3OBrHhsZnfAlqug9v/I1yNyzK8zbD4txgRAZoerDbtceL1BGJZE2po7oFpHvK0C7
2kKG2QjtY8MIqeyoDRj5NLbO2WRR8NCFhhhHLqGwoUJd1LiKJ/i9yoxwP8tfVuLn
hasxuutttQ0FlYoXCykf0ElLmJiPVOaH2WBdz8r8H0+46Hg6kEChDeimkCoHJzH0
682+sQyhVh9KslpA6sfkXsq1XTYxw/e4SrxBpMLY8R89F17o910X4sBM4dRZOAeD
wpQtYyG252cx3K6fmq6j856Nw0qD2q73lAJPCk5wBOwUGiTCXMglBCfHJgZJuwGo
r+Ros1Vqq4nxSjXtZFzZUsxB1C3DH97VUEArSHCVAaTTJ56RZ86cufmV37YuICNt
nrwgVY0WSmEpyZLOtwx5j08XclWZN0twZnyEqYBIOUah0waJsdyMr301j8y3VCTj
rltKJuQAFMDjy6uGT/xNGM37Glntz3fzyd2i9ia/jM+JEs0vyjecaVGH3UJnD45j
3KlnurjOYZN2CoKvhsiAb6HpY+KOPJi8Otjxo8agzlRrd2w6qAZZBKRN6vPflvyy
ETK1gwTU83lAuenj8qfBVaOm23XQ9+BML/FNB//J+5i5eOYNl2QU0kbOzVXV7gP6
GA3TJiqXfHf+WghmflfpxeuwkmScX546k0qgBj2M4H5otcihsANfz6+Y6xcOpEVo
VCUr+XOVKqgP0R4/VQiQVm7zoBZipTEWRvB5AC7e+SUIvnwUfB+l+BbBp+H+wJFw
jtPWgcNoQvuuSen5jlEXr/pHo/nvjQT3DjaqFe+wXgif3xL6u2KIlTxetWG0M33t
Z4JTspCi/3cve+4/VaV4LrNEl8r6jLseYLS9QRzyRaSg0bq19AbHRCBwqDPyqqrX
zbEV5dCleptk/aUzJ+2s/4yZc8mG6AAPfobockYfodUrW0dkvWwaA2bpGzzgc4iu
it1XFnWAKCbTLbPqmDZr8HpgyRaNUYtTW0vFvFosMkR/UsH9KzxaUwG6t4Z5dg/N
VffQqWFOB4PRs+Fs8hnQzo+lZphfY1S8qSQyKxytKBKQB2/Ftirv5oyOIxY9qxOz
R/+z2zbp5N9uaGpR0nEbR+33GM0o6adU5xDwCjw0VWbQMcLJEbRHGdgVrk+GqDu2
TMYr/U5KqhxvPW8JP9yrfgBV4jQVLRLebzfJT/FcrLDS29XNdRY6/VO17Ggv1HFb
tXN6GyBXB6S3AwkjyNZ59TVEsr75clz1GovhgR3uwaOj3FzRiAC2zIIeV5gR+c+u
KPKYnBSsPHuIZQDW2IF1qlzJoOrHy4TwshEYcR+AchmAm0dcDbbE2O6fkjzEEcNS
P0FYONLfW4ySG38nz+usMqX7CDn8Xx65B71W91whOsLFzWHeoPjT9+cvF4HGWUUq
dWNajSlbxsGhcihYfQz7w0hcjkFiBZLXQH+Hlgfl6GMkbP9YDUQ5rQUD2YLmVArH
KlJGfJkuf9piOJSurE5n+jfXYkayJqwMCMVMHdV/ys5oU/AOP7+fkFzIrXn3fk1k
E12VNU21U83P8V+cEFQozLcsFdoWR7JdwXrIJdNWQ/WsrUKhVVQaX04XxWaNe1DN
8GnYJqR5O8TQAzTJyw3XdlY7llZnjgMXXexSHljY2ANI+EZbNEn2pYpFlFQnP/Ov
avg3/QvnCLmpKnfcD28coLyt/motFWnxu6Ts8gF8KdY+gFb5p6GAwta0Z7dowrxk
xFcJtYa8B3tWfL40wgtGgesikEvASBVBrFdhMyPTtvcP8ULaVBbGzIoZefYCBnyo
tp5vvRlJzG+hvJAz++PHh1lnuSakIVinvq4a++3HtCx3Siwoajc3ahLfI5a06K1v
4FM03o7yjYCCj8xLtTXP2nJl24NetOHU+LusgFv6UIBginXLjWOoNyJPpn1nk45y
6YDvXHWpJZnL6fE0+dkFh7xwhDiRCFasyLaL3WUJ8A5dS2odfLRYkzIoTFXl+275
8pq6JFkG186h17fk8URoq/AmLgQHfLQXjBxpCK1e8YEOE/FYqiTwRZbQ3TruiRKH
rIkZVmwEjHpKltpS7zYmb+pwnKolXitk42pkO4DVwDlu+xuShNV/D9ntXMRkR8cy
aiCfG/b0TK0TQHpCMqJD5Hp1kk8XzJNZQUk+jfFT8nloSygrx7qX9DCfp0HRC2Sq
IbyPqor6fIHu6Sejm4H0JrIFEbpKvlCUi8giVxts0aTlV1UpD51z9jO0vqDWaMDj
qpJfm1epVN5DGo4vIqwY4Y9pKA7Zth6jRQwhjbumldE=
`pragma protect end_protected
