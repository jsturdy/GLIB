// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p60VxY8Ne74HSqB9RWFPZWlNvJ7SRgIG4wAcb6S2N3cnYOqXpeEsVflImL1kKk8O
zdCHVIMJ1IRU+Y/zVCkR6y2o+fd2zwkpaGYekWqsf+sekyeEt2SleVdndKfeEokG
2XK/hNCTccGKziiFn1QxZKHs35iAUNgBLsGfL58ekaQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22864)
eZRK7LXcPRy4YuCv9jNHG7Ai+yIY3yFBNfZNiVLRxkmPbsRz9G2eoq6f9RSdtI3q
7+WVBcNLEq8d6L38Xyo3YSnIlnO4yQEm5ij8i4dm/AvrGUQzeMKWi/kq6sEE4bhR
zMZHAwkw8eEQVP9BmnzRyFHSENwnYiUoVc9Ip/9rtJ8HapCIxA9Slb0LEj96Qqd+
CXF1IWT5OyLgUNGm4brle03ikGU5PRgWrJE/gTFgqlAEbpfDFnS1EJHNKMpCipXF
9gEG2jJax7nqAPeuRrqppHuEO2546r/9iNB5IP0KE7OajmgFCEfIIWESfkPHiGeK
gbhM3Q/GTbCwptnrIh5PrWfj6FVQt43f5aBDA5lOl/+Ch0MX4iERLxCA3r0Ao5B0
vvctTccmNgY02PmGOfmXgZu6ItI00DrWbn/gy+bemAhjcRUSyhOT6JH0FT+poqX2
kxinA44ytC/dQQdcpQ/IhZ0gNwy5U7LFWCsh6edO0P76n37XJsx75F10gE9k9tSw
4hrxPKrbCq+a0TEG5DwzcvMxElIzkT5Ykx5wNnwVVzBmMP+UjtXTanWiyCTmO1gq
5nSJaEb99MMRkC5Dlz8Oioi+MdpQq8xfKygqkmIymDwuaEtkfW4mOfwoib7EM/ly
fhvrFjkd1AgyjrPO+j0qwLkyqhp+v5dg2SuOtX5npHUzop1dVz35fVzcXYW4kk13
bDQnvkVoY3TD/enYj8AzeHrD+0txf8BxHXJ8XitK0MjsJk/ccrM4L6ojVS4+fhSa
ec0gkq15PU44IuVENAL2BxlD27Nf3Ue9Ny0riKbgh7O3wOk57ktcQIBb4bm54aqI
e1Jy2OyXYgurKmt6kOpdCKgRAxj+B3MetgMtxQIHR2oDHFFZNkuQSfAdEHtWJ2rJ
o3TeQ5e6JP2w/UY0yiW8EGHlhdkIVCjaotemftD9KaT71c60HOwaklk1P7DqiAAC
2DGRdvYVS6Kyt+qDcYFv+flYRwDgqckmAakmyP5jjASp7ggOE6RZT1Xg6dkdMet1
g/hrXTlWtXvOH3x9OqpdeFjCT3PcSpIte1BJkM7aqH3QmHI1d3tTgPCXvWKhyJJK
IwxaWp5X0YNo1czsWrXrOkQXgcj0zGtwjcz9HHlrUfvn+NX2zhyS9vp7MHue00jR
fvjF+Iow8Mp2J7B2ndFITSvC0Mu2M/2xyBdtuhEHju4ROO+rcoJyOiB/i2GXQdXK
6tSfmAFcpIkjq54Lts+3ZXRd5YU6QoUxKevOc/bF+ZVVMvLcH1N1W/IAKbbDMQjc
TLyIUVTL438i8abk9sbwrjw2v+cgzc/yyKSp72Vhq+DS4LTROjxYkCvHyRzdk+Tk
YCVChANjH5tT83OW5bLV56O8k2pD4MzJtNJXEMl9oZ66PRGgcGGUmjNYy0+3KuSb
8fIXRcvVZW4fOPKXuitGjD7YdelmEKl7552POBXH9gsyM5VeUh637pfIHLlVfidT
ZVOq+GJJPbnukxTPBFyGiLa33OU9n9jcIYBdQ+FpP30Ggmmw0zun8ktsogMT9Qx2
XZrwetlvFnm1pVTYEj2pfovsKBnD8/q9xOaQa+HlcK8MyYnp4BzvqFlqlOhqIapS
T4GFZvbWC7d3OZp0hOot66vDcRtweP3VILchrobiEOzL/ks28WyMgiPk+1F1ufPn
dacrWKzVNbncFn/bvRzTeprbJr1JO0eOkFdyQlDInzX4huuHVq14nMr1w9UVJblV
qKiIMGQy0UPc4L14NhDdjSY+EnFeLpJTbTCa8x69+e794T6SBcrdKcvvGiOMdlBv
gfGeVhO227I0TgyM5zyfJqB+8lNFdxIVTDQRjQWivb+nkVLzxJxMLN/N/g8wb6vh
9IUkj3qCguv9whTv0wT7SvCYowL4HeJAA5I0saTOYOZpYfN05NjdlPNgKxjDxE0P
dGtukjeOLUtouwU4HAQaIUSMWON72esYrQrzWk2D0Di1YtlJHdGmm8U104teT4pb
t+BzNDsLpA2q2R/nuwrdcafrXUg4c+1gWYATv9F84rkouiZqfQyXTWAeQVWY7CS2
IEW4+7O8P3uXp1PpNTKygFPwdgO8iu+Xidofoc/4UxUYh+OeR3B9GaeE6q3MoLfM
Fq/HLzoN3mDVZogxhLL/AEcaeeX/A7vzwszTdDMUeGcIFyDwdt5K0aJhMfizHHHb
mBrC9VTGNO2JSEXPkWMAZ8NV1Y4uYvGw5sVYE9Qc1nbRzyzw1HrkMhhfVrVH5zYs
0HSExzHGKvaky8XutLUbvhQdi2BWTqOBckq6Qhhb69v1pKy/kLXuSNvN0Ost1iqg
ZUreDsGndoeSdtITTQUnJF5Ls9Dy/mKmoi0vw9mWAMbQkKoOBZsRr0rUBiylhWZI
pJAtmbKlzyecpxi6+nwXX25huSezOIYBnQ/hkNM/oVwBpVBceHl6uhVTK19pNEFn
O0Cx80ir6k0EVmnfzG5d2PM6XvVREWR/AUJ+ulFljHpnWhFc+avw/sehJyoXwSBJ
QDbi3lybbNW2YGHHBMDFfmTzDgV9CgnYT/bSmk8E38JAzmKF9hh0lan36HMlN7zG
15sFbtjGb2wyknXD66jDgnvHNyvo0EJqHRkSjuOL2t2Cd1MGOKZLeZLuLW3iyeao
j7dUnCJZzxf6UQaLfBEgZu6IudP38t0OfA21ksVLfiyKjd4wSisP+cN5VXtIFeEC
pKe7rhXfypGZAenZZd/P8GEGggcd/mfCMknvZbKMqAXbyzuCh4ujHhM3jhG/bymP
BgjQy0iaazDNKk6hUMH3+0PraNLACC3xUXtfnv8zSoLWr4agnDWx+h4E7Clyh7V1
6JTSmRFd8VF32a78mOrI441N1j42moJGqPrAOTeqqKu4AwUQY8tO6N+19lgxpBIs
0s5d25vXKK3ATpV7Qg9isAtNmxluaTMsRC+Oy0kCpSXSROo+ZiRnXRClJWCj3mW/
IKELoKSfo7wYXjBVwdKfhMvq+cCdX9XO0EjvKoyiGQbRNsi9Fn8DhMR6TUINRPXA
+K9rtmVvZOC3KMLsmQcyxY8DPNJrEWPa4qAL3ZdTwBgsU+C8AciYp8ms6J4n+NCu
S9GkawZGzQBkN+GIRL/cJZfPolZOyPHIZ0kcVfmXRdjFveWcSTWXnCfidJgakLAl
k3neNacRxlKeJe4areMI6233eFqMSxAOTFL6rXwdyiXJ/aM2IOmV8DQTYRXMUktZ
iObulx3DjhMHtymZfLR8Snyut/86NanQx+qK/aWOBYFV2PTYX89roqOmgrb0UlKQ
1UJqT+FtoQfc2ArdOhNmGN/pXXC+p3hzkB5N+Ai0unPb1ZkbjRQRtcWvxAd1WKB6
O0EhFcrZyXZBCi3HhvZlZnC7XFADVc39Ekt6j0DlzVMsYZSUPMeZtG39TH3eYzbM
QRx8LGL1qFhpE+vfamSNctxWPZ+Vhxa5VjTpGr9oichofsPUStBnPaDzj95CDJxl
4P5cCH12mMm1quPP7IHKNwAm/FfA1NqSQ2BB38TBjZ3R1rTK/6ILqblVSJScV80U
CVvqF6YN8XAvdwxG3fyhiLAZHyAchx+MX6lQinw+UHRUUvJsxsMrfdPq6hH9Wxmn
Oz/KOxoZhZjFGsuTcU6AxDF9NraRnCP0claRZ62R2qBSmzgXF+ePx9ZwwqbjvMSp
iIIbuKq+eZcYSvtCAD1+Q351Et1myrwGEPsfdb9bJxoDU4vmeGMh9I5O/3KG/Azd
aU+Fkk8hvRk1wo1fsmaCn/hyUG+BSFxGUXsxp+znIsNCuxWHo4oBP6vv0PrRO/X7
HvyAIAdxZJ8tb3t5dv/HJFvuG4E92xKBCmjAmmpuOcVV7xgM6/tp0ZYwT9UaNhS1
rDQUJnZ51O1FxB0Kwm0jhSviMj4VknmogdNrIRVlEAw2VwdnvCx0uCoYfFCSxIlV
N5MkFhPkc6NddrdfmvTLl1aWyzCAFj2Z35f1AuAB5PtuhnVkf3j7n5kMkxua/k8h
2vbOcSN3wE+Qv9KjgRjqeOho3/izU/aSuB0gMFWMbkSH+ob8rXt4AzxZc7Km2WQA
j6r5r0BuTwCt1elcQP2ZG31kfILtpEGsibycDjdr+B6+oN8vIP+/k7O1+V3jIhq1
8XwlX6s72YaAiWDKVATyR/GdeLXcafJa0gYigm64OTmbtcK6nsr+8QY6IXsaOHfW
gOc/6A+5osBnGdTzD5mCx3FB5wYKtQM/feiOvl4JNULhdEHU8uuDIekJyxzvFQSL
/73fskrRNr+2hGoJFOJZ6+DsuiuFW5cd7xVGoTXOkpLYZmFfO88HnP/o8rzutZMA
DhtC84nysommAjrqPXi19pmyVJh+f1ugypLtthmR8NJ56cu9nFz5IArQXIccfiFk
q3A28Qn8/bbnpESO7Tgxmpuv7Yoc8pVIgsTgstvScBzVwcAMjoDWSvEmffbSNe2z
KYLIi0rKFiXtazlfLktrYWHg8sOiJBKuI79gTJcvV3qCjTXq1EYneUn36mlyS459
01bahHt2v4FtgtjsePJRGE10pFonaQkLXDcVz3Yo1xnJuf8MR18BR89unkrl3ocv
aaugW/7Dr1seg+03LIIL2h17D64YXfIWUqZ9yNxJlgHpildY2eHUeooH1t1uq0uK
MrPQudkNaoyoeiuJjc3rmjsP2Rgp8djiDISAxvLdybWA5FtlopWueU/QVUeRQJzH
glhrRUvVU5uQPJwC+mk2ZiL0Ae4GWT7yOVqtT88e68cfzrXej+2zWiWx65jRUNg1
Wey1rIgE7aSU2SMji0dH0T+1wxezB/BlfJ3tSOoXfcIGUmUShmBWbipCFmfg1zYC
7Jsr8BeYou1lQUU20we36KKLpxSGEzxs73Onlpu8LWQN2NdGoV+f6VRxmRRXxU1U
tAPcI6DeYdk/K+XXkmIiR/TBi/xqs5gjKgwuEQfBkfH88wjXkddRBS3bt3mjDGfU
1Q6kocIkgz7jhZlTfTg3H/3nXOeYyYMsRf85ZbEw931JeZp5JOfCjt9fPIt4O6eE
0Iti+A7RC+rGPZkg94WJexZ+/w1Ryi5qSodh7drdM3dl4TWHyKtAllkNMl9GJi/G
r9hXfHZm8Q7jJ8c9Nx9IRbU7y32SxS+2pE4o4GXWt/9qcj6kV0NgcvBn+fGzaUly
t5MiaspU6n7yOtclHnzU4zW+erA0lsny04KSosPuL4ofGsNqcOYH8SrudD0NrgBP
yIzFm/ZE9cUjSQ26+ZNC0+OUrSBhWW/L4HvzBWezSqYxgoMyXUlYoBSL/D/BD+yY
5hNiU0AIGdPzyiQwwBETVQv+PsQfrEPx10bqDl4bQ/fdwRwHuAZu8RfyeQ9t+u7Z
GYRmGf4kJJUJqr6/mtg8zBTJvsoQfJkC4TM6NbYVO9jAYO/TL+iLRxKmwjaFGh9Q
v1kOTR1eht2CuBmU3dgL2h/7+mHwnnI/Q3ZoUj5qE3ry0wyNwhuGf9uooGatpgV0
MDx+qdcHG8tLr9bHFhVyU+4UeO7K2UbaBymmIA61rJpNNy17lkwc/AHM08pYQ5kl
pNfxor8TJFzCTY61XIDrFtKft2rQGtHOneGZQ0zMmE+gTbbnShsqyPSxE5caY6wE
U6LE6nalaHQO7DJdEGGcMNn5cVk6iG66ld15piR8Sge7aeWBA8+Ro6BfQ0ZA51KE
1jGYmGzBUzsOSOzSZYgbymJXmSiU1+csSY4i66XAC8gVGi27/wV3s++s5kOmuICO
OArwgyXsc9cUvBFkI2mu6Ip1i3o8pWiulKbxzfekt/GGJLFPlYQXiVtmWdO3cfp+
XFzDxWura2EFfTBe/eg3qlJVdI6yymRFFNUZvCZ9tyVICMRiw90moJCHtSqfK2IW
QNaWtKTtCsqZ83gEdJPCYNk25O2BNWbENasSawzNswYMOP47BxBqe4dg7DfiEqZr
e1A3m99HdMdHTm4sIkK3H2mTfiCLdwhyxZln4okBSxtxtzc/Ytdq0lcFngw5LV61
1tA3jwrhRYtmJ1G7kJlFvKR+KkYRMNHUT0S5qt8uEB7V43uHmqKaCC97TEXo+zfW
CNL9dBxcMduZ69TyAQ8c7vUCWhwKnFTGn+jkNDGHbjYIKYBC3lK13Zorg9Jv1sIK
mOHWmbSLrGJIuaIHk0loYxQTb05HdfYo4cdb6EgGT1EdUaxJ6NhmpmbXMCa7/FGq
/lyTDiYtavkI8fG6idHCeQtUZ/nNp8CSFjcO3NtvRz/+6J+i/MgbbujnIsdkbDQ9
np8Xw7AayW7QH2GOjStqkM+H1T2y2rBHgArHNEvvm9s/n8M1jwHRfIhDh1kRdVAI
9oYvKafvWQSCFRxG2MaqSMB9NFfXNgO0RLATn5t7L8vxek8IOIVTrNYzwbunEWqm
tlLtY1vs6+ZGfhUo28TPCnsKh2KPjFUEVuMq+7AtcRMD328JbYy8NiwXXdwxevjf
tqy/tFRxe/arZrz5edNQrj8csht30DZQfIMfV/2Io/ZxgVn9YDqacZWom5V4elhI
mdChbnpyd5gmqSDiCQkEhK3eTpwpp6oj1xe7RkHFes5Z5qsdvpU5ydBY++/4EQkW
mdANL+kN6kV1FHNSqKQWGVCmmyu9j72ASPUobrv8JYLxsw74bDzIzezYDKQ16l8l
Wkk8TqKmCdeDVgAD8RE0un2fE/cVNDShVxCM6sp7grmDwcZP68nOEa0W5tTiJ4g0
WoQ9ewe5uaxzkymmpwm+EaCN0s73YbUS19cIXfdBo9YhYtSge3lTCSChQiON9Cii
3NMpt8OpKJkrtB27Rmuny51Clcc9Tgyh5Bjpc/mD/Ax2jWvlPV2yAbcwyvIUk/Jx
Rs/uLz9rIu6rEEv5gsewcd30c7ntQH3y/FiNWPuoAXJxZr0bPvc55hslxL5SrQrg
k4S7pir/T+wiVjWHfueaV33gc8rr8YmpF2dk0EgN/DYnYWI5SaIFDaTfYcW+hCTl
8cwv3XgqY17ssPXylelBrvlAzqH8ppLaZ+MVvQbd6X+K2ET0DorOd1ORx0pKv4jW
FXCUJz71ATVI860ygy+RCPknjRf9OL0BMJTif5zg8IHa+mV1NAbCLXSe6b3I/Qwy
qLKxGEzg11xvF1BRmgffKCVzA5Tj3yn3XBgzJmZDoxVbcLafqeV96Hrmc0eWsG5c
/lf3jsG+CdCCmF2WKAgujclFRKewp32foLOIYUv155KA6ogZt7Vb3QkHrMJCXtUc
JIQKMHOflqSBXP3TFdHmDWO3zWulv3nb6SdMh2FzYSJBMnAahQ6b0MzWfDxSLT/z
QR2qd2O87UZwe9FFwxFzSohzZyf9LYIZgtovJclgMM/AeoWIU+YqmdLOzVwjr6+P
sSfcsz5QKpmyPK66MSP6ZQ7dbyuwx9HQ6OZLCHJXN0bLRfGgZgyx4sMMqnuHcjNp
b1QTvGFXW8EKwCSy+Itpo3wMwLZZlic+rALyfFW7zbTvdCxjiNxdDsXX4n3X+V/b
Oe12xtex6JKJkVCKp4pOL9+vsgBIWZAOmjkTYi40OW0/3Z0Adi4b7j5TLvtktqjY
wu4UDSC0LflRAKj89n5Vhxb0HPv9c67qEzod1fgwvdUlg0kYN0sSumS/4ZBBNqzL
Wtll1zg3Lf/CWVcdX6sHKkk46GwvJ1IBDQsBeOlLEIObLRTSYS0r1F+5Ngex9ytj
eb26Xlkb3QHcjqvySG9WpoVptE89AnCZqRZ9vlk9XaDY+NO8sdvyWixH8VQMfDLN
hH6+HGoWhMhjmTmtUqR6ckzhtiCbIDqToodozSe5On54v2TDb0wOjQM3d5+u0EK6
T+nQXeL3GaqJVqMGeDGUUbccF0MGurV6pUqon4DXe/BrIga/EaJ+6ciL2shDaFhm
ypQYUcmWv1GjBiTiQgo1HWo6sEXenu4OTwEjFSdIfYGZIPafxyxng9X/LZPfWBG+
rQlfWTx0K+7BzlM/HuuTeeE/GBxefKVHRTHhXCZwIw2DVYZJv88P8dOkRdKgiX2Y
Z+qkVlEv/9MZ7ZVrTxVFZYddOG3VejnlVTa/iARHLt1jqZLLQ1JJTzjsUNwCaVYJ
sCvrYtxVf1QTV7SeYW75nSqiOyuqmrt4pxR6k0SgRA4cJ0rwmRMV5wNkARz7JhwB
7wBlhQt03nn7r4NteuRXjSszZfy8BcNpoeIS6XVWCY+xJg6duDBFy2nvJbyOhPa0
j8K0BeILArffUQo977oPIGO/MSAMof1nj/ZfuhRYTIp8qG8Czvr9MUFVZvZjGXhZ
AOS/QWdqrn5YWBDG/2wHbWYK4k0CT//YQTICWtP83POkdSKIKH0Ll/64DY1dc904
Z7oZRkXPgVebqDhNhkp3V1+G8qchl0cgtnosCeQxKdpwQYdL+S5Al9lyxbuJBpZ/
ggQPxE230OPuXuPQx+yL9VzZp1TDgH0EygineePGOLI1s+yFGca1BBiNto3F4ZTP
W9I8UaMtM00BH9nXzfWqiWQ3/ay/WklyF3ZgVvP0CCW4fMvXedAxGcpRmg4x88/0
0C/T21B45BngXgtVqnDSWC5CDxFIzBSIlC0Dh4rBknWVYXMkjKmvDAJaEPOYbr4o
9hSRmVokbxnPW5f0uAZByBZoZtOMGftX4shMAXMzDezzNXmYT7bWKT+rzw7nJSZA
oR9WixNBCZ6WINc36z49UTmfFNpdeQt74vKpdW5762lQOapgtxteY4ZyjIC9faMn
10ErDYpEapJV26L6VM9GqmayeRhk2u2ybeV8bHnhPWbh6XriUxzRwD3uqiqFKbph
kVZUlaCeExvjLFG+7nQu5NLTSqbiWsLf2FLhNsUx6Y6bY6pbr4ojJqRgQ78acHrf
zlHSj8l6+hQex8ixNKnMezp1bkrJVm0TujCTDH7b01XaZG16fRTCptpMJijllhzy
GUiAzvDG34lps/RleC4/doLWk3IDQCqZ5ELJHALxEZvTM4jisOdIDgH0Q5Mt2rvg
dhOpXro0g2vwg/vIN8MjAEfvi1RUWiiKhE/aHG5a6Tgy6wCmzfnh5TN/USp+DqNe
fI+SBkUDPrPXTsw2BGErR3HL3ZpvZNJowehOj2j90Ap0ErKeIskHH4TvsAMirmwN
tXb5tZ7STAIQJjcA6sibfiifrwNpXNh//svPp5oU1Ly14mg+hYfXB90KyVs3m0yo
CfZbVfjUSopsu/2vKIMiQ+TwmYO3Vc1geZGd9i7HmGRDkyo0EgQfhDX9HhOusBFy
tjmyi7pKaaN4JUOyHzmppcO4pgvH4jjqYKURynotL7ElC0pHlOSmErOfFixVCYBU
WLWoKElyaSqXw9CpzGNaQrNjN6qtV5aJinK1TAag3hDVKuTq9Jz13el8bpaJs//g
sMrP/mMbPVukB1PKmV4026sp0hGXMdssSAGChGOnyguz6wxyBV4ei/Lf5qnzUMFW
4IbNXcv1a/M0adIB7pNYjB6nOI5w4nsrIng3gGDSrCTbcWh5hinMd6Ka6fOmrYw0
VfaRE2YQqNZnXuqBWN19i8+HbCbiZTx3U3OCsGCOO+4g0Lx1PIti6bbsHElbd/V0
X6UNCg3kh+QssFWXRg3o8f4cbJgkryOh++jrni/2trfSEPnlIyq017DX+Ou1Y35l
STMQlZHKAtVnb11+/Y6WefweMTPmSUSi2hTkPc0Fohi7fOyUfYw+SWWxhwZQLFeg
lrP4oKf2nfRd/djTTP5UXvIU5/CGUtuFV1sLa0F3Wqb32QaZZNjKtoURzI4ObHsa
ZBQAhRfK/cz608G3VkFcBvAmR4GieHZluD62XXn5BqvsNOF3tjaNK9Unti7Qze47
QL0Yd+q7pX/ty3TopB/UKDGuytsmT/sJNiwZZ+c5LdcYEagz2NIY6IsYXn5pscB9
eyfwWsAcENTQ6DDioFBGPwsLmmObSri167GoKNLCXW9GhfuyL8eOxg5P3uPmojSK
Smc9OwJdNTu6CgG43xVUySmG+zs4FPqMQsJCspWA1EI2wrrQTvdjk2pJSQKjpm7B
FAPI79Dff6QSMjK3MEwi9t6Kb3SIZQS2YYoaxRSbB8jwZAMtBGNArtHuAXAsTt70
LC7qN88KQlv3mKdJO3s1TWLaRBLR53o0n9vY/S6JXEdwjhi2nQYFsJHV0tdyJ1Lh
UHuqZ8gwX3McNN40sHXH+yNTyLFoYfBcWqwPKFR4Bioe275turxwFtjol9o+T1oU
pG+yT5MFr1vkjSsNY4L+Pi2Y/O9NZ+yfhdYLNdfKK0JtAeEvPoMWmztpzO67IdBp
IBnYPMUIPJTP3+fOfhKy/M7S+mqv7DY6fzycsnEhJ5Z4Ng5H2anMEEOv+678XdXH
0ytjkiaP28QTP6+YWnNotph4ALITuvO/v+R8qZZYlwwL9w2cpdVvjbf35iWa+4lj
lyKdU76OzhdpUnapqUz3LLSKDmIAfccsGiSJDLL9E2Qdi63XKoDd8UVAAY5aeBlZ
Ig9rb8QmBtkQyCbHNZoaG5X57aeZhjdW7XLI9u/z0DylA3y9r5Oh/YupPykNDAfU
6bBbl9BXGJPy4553OpnsytN7JDNhwN2QAt4ykXlGKt5c9Fs+ySVpaOZsRPLTy/5j
zkTI+t9zfQvyw9uapVpafSgzzD0+eU113jP6o41fTRyi1H2K9U9jVTcj9wJTcwRO
aRgq+PPfLafVRF/VzamE+b7tixkXhOkRBPc7UPHKgUaz85fZY4zkiqLsOFNT+zSj
MOLIl+VOwKl3qUZef9jVTnbPbvHLk+n23hFFyEkQQchw5PxGwqI5zuRWMuIjkJO9
ftl/JpyqzikFbrjkfhYQ0ceHwbA/qrG4floBd4livKaQy2QRzudxq97pQJgi7MqL
zM6qJMyPGFxTPKBbjadd3M+KtLs20PjS/PUBfuZurqVDuqrdoovm3jj+BukFm2zz
xIicq7GyVZeVuwpp3K8s3IhDw3Z6kTG1H1V3vX82eiZf1SF/Y9RsuWCJhwCt2PGF
HRIJ7U+jElU/eTmq0gdKJNvYr7cEMrUIQ4lItC/zVHTDpvj/sKFuwSxePyghjZPE
LW5BSR2EcqScdVmQELkrpKrQbTVQF+FMtICLfcp81Y07xCyYkRNxGnRbBqFJ72iZ
e1CUVe9OLisMMxNCwq9xC5NQuS/JL0vnDujN/+y18BI9vEC6qeV+61599VlX21ML
GkBiMAlGH1it90+zoYd62jm7DZOY+7P3/In1rjjZaF/qxIXvPoOq72EgjtCvCkrW
mfsVc1dc+iFRy5JwSu9Dfsy3QTfLRs/rKquqLDmN5WSlygJ9u4Im8bwelgnATfhl
ReVtRhH+LbJ4lmreFklp2+Fkbe8FfmFwiCgEL8Q2l1FKnH4A5IDZgzYwM7BHFv/t
CJRF6OhDVUgpIqhv3EN23fnyLlb0yQyOdE4juCFFVjhMditAtpkLOAdkgb54WY0d
ERs7RRYIFDSaByQOo3jsLwgUPFth9wfqJ6DjIq+MAVMsiPw7Np8iVs0e47d5oUqD
IN/XDw6Ja4lcpXXoostmWzE9XIVbikRkH1T55t3/LQKhpzSCuN/FWg6L3ItkB1KF
ucZk/ugoo4ZfjnDuWYYLr+SG61z9sKSqoCq+1Doto3uUjT+54krQPc6vUV8Ing+Q
wIdHSzRijZrhDIrlIyOcUEK1o/ambAQOUTnk3YxJZrcxEd1NgFKy1vt0w+1PaW6I
sA2KA7ZRy4sznZOywV8o3U0E2zK1ZnD5tIGN0nWfH0nuTuto+CP73twCKFIpSjlE
AZqnpZ/j3r4NoMpAEnlyqfMrqvwlGOOyiBFAhbQgEIfgq5Ok4LGlPpI40K0zLKQf
jkpUtrBfRElinP8mfQZYD9iO7S/LvwFISiQv/xqauKULUM1VousF5o6GuMrzp3py
59MtPtNCOMl+/ZMKtlrlJAEQby8jLqFf+610JGqFIvQPiOmKgn7pO1RRNBbcYkGM
zT2HubFV+QpUD8y/fSC3Fih4ldNkDCQYrT4RwaoFqhHYVOmsB4xvxnL+xeQL6qLe
kB9818qyhXL7fTY5ZGgqxoqnxhQSeWg/zetGPxbWdOJBBufSRMb2+G5GGUjgl8rB
AAEsUkIYOjjZqndTtI1Bdm5/AKnff4Z4KYmTghrmg9lQt2LrPdkQtTJSTqG/hRiN
qAo2gYOi9rax51G+8yC/jFXqsjwNHnzxNufyECCtiV55tPfo/iVA024dtGOuM3PL
+QCj/AQ46PmL35krpYMCK6n37T8O+/Vqsksrw30zRvDr2qrmHl739SMBnyxRkRH8
K5zx/zNXdkPxVbd48/kVtlLJzAp01m6xKadWl12f3KJDSSP0sO+PDbS0VQH4IOSn
V7yGROAcHM3wnGbhOdbBwSkqbT7AmwWfOxiI7wvAM1z1IWAKl0dI0Nk2Rvjr/Geq
TNznBwoE60E7uiyPX6A2tM70Wctuc86cpcesFRMd2PIc9OxbJUSf/J42PumPD5yC
eRshgrQnhHvGYJ8SLjODi4KP9W35cbqhqP40hHKq3mAPEEa70Usg/PZxSO7EUhdT
1cYJdcje6vd2vPd3qSSNQqd8dUfl2NmZYDSHGaLldJlVS6vbzx7QFx1Mmtk4k8ry
TwzAh5IK8PSomQx8GIWc6Oqdpvlk3YJdLOg6NP8y1DqB5Jx37lNi8DxJkoE/VE/c
tM+Gkb8I/I+JdH58sjXlew/+E+KwxhfTqJpz3GIDDnEuxUKoM+5XNy0CbfVXHTUZ
dTlE+Mx3d1GeMMo6Exrs0p6CyjIsQc0QzKcCpNs+RtW6Hqr9RUJGeATk50Wni0KH
qEF+clh2OezU7UizqCR2yk7PbiF0sTUoZNFWcipSmP0RxTN7zMeBnbg6LF0FWI39
DdQP1Fp2Ybr4WAkloY7qHZJaRbSdw44BauUQCxkENW/dYB4Uc1b1xjS0GaW4angX
gq+ZnrZsW8IdF7uWx6SGhGs0M2RGUz9vF6tLlaGBVDa81+Eg8IDIB7VQlaRrDP7M
XqmzRducfEvE/sAHCp3K/6PB9Ip05nd8FlQt8XlMM6miVLtJs/QpCF8Mrmvq2Tkv
ip0Is3sl8ViJW3zeGViAh7yhu3AZIOHmiPXnboWKROswnPDaAA4xfXOrZORRT+e5
pgnT8ee6/VARP6MX5uNNLfV2tcKsKq/PpK6Jwbhfqch2xX2J1UVOeHMun9u3RUH/
5bX8ZDCCevS4SgXyS1/E4NyycenLZS2dTdRxLav+7nsL0ohEHcPkCtFz7fufxpsy
Ulqe5P0Zs7qo06W5ujHxPihDOBsKm90Eb4NSCjvFZO4U64Tg42vTADBYysDKX3NB
Usc4glaQQQ8pm+PpI7eQ8NBCT2XKFTBrYIFYXiZg8uZq1MIJkG61sMdCR1ZrkFML
ZjVfBeuWzU4WN7h337gZCexi9/0vVXFSX1HIl7QatkxOaCPhgZpmWQuT6bYfs9HZ
IGkU9I3qoPXO8nySjpJpbkqMjReawebOQgDvGE5/pcbBIZl8lbL+EB2rFegCaCxv
kV5mDwnIxM2pkQ82pKydKU/A6m3RIoX04HUTJ/LzJ8yZdYaokuPZ8G8WKMx6FkJm
u9XBn1tbJwkywsEaAsWpfuFkLFoSFcF0TShE1tR0DsfJh/pHG4VnhjtQqSGkWD4y
wP/YHUD+JpdaqsGhYNDONj5M7bLo0lcESnGDM9KvF94BGgxLj3+gJM1HNHsjEe9C
PQxpd5v6KeFLQJpDllbIGF/jF3lEZ/J3phBX5z/CwAOcjOJfaYt3WVqQt7MJmOk6
aUlFKFbBcRVS8z+BGqg4m42oAmjyWMezDjL2+qr7A83QQShkOdvz483T8Bs1cTuQ
LF0LKd3/+ms6ppJ8yWXLr4AYCQKceXrOxr449gT5YX6zQNxK6ugD2rI3sdA8vm5N
lM4CeTsODCnE3Uy5iYOTSuJ2ZmCNHGS9IhCeNfXsap81qUHFX27s4Ke88PP2p+NL
KN77VfictAjA64VChf1i/1pK0WrVXLRK7IKgbFNNPoP4+lLhOP+Y3yb77WcEB6w6
pWSepAaXbcliPE1Ojpc77u60Y7YzEQyeSPbby8ZhdP8X6P9hpZtrXBR1RV7sQt+R
pSZ7I8SY3XgETzBNDBAXsIc+BagIAL7/Os2QWsEVj3uoFrHyxCNNjG8lF7egOdQ1
VVU3u++YVCuCjoY/iiYogehtE/l92WHtYjWVNEKW/A1JNoX3OIA8lbs7mL6ccjKG
9vtnridrKtIMUpfwzvw1LjL8z6LTqOS6Pf6MgsgkrtANMGi7ti7TbhgTCVdTeetu
x/uZ1+Ge4I68vm8O4RvnApUuZFsGa2IEH6HgDtChTU7AWh7is/G7CK8q8GvJcKLt
E4uN92zgT7uOD01gAWrYq7gVkzjkuXopNt6PcYNtaQvAPt6TrOHRai8uJC8knQLR
O5xRtvfOLQPsfRerPnvvm6elClbokE8jzfI1AyvLHjLQ8CLgv6DGiNsy5cSAhAKT
bR0ybtEU9Gsdj6A3SZoTH9dAW2y0UWhL4hLmbFdEBqmB+zQW00R1OASsiTWhrMJI
ymsylE1oi0cMBk/9/r4RUdiiXMridQSmcuDCUwYq47oAVGg7y0x2O8xjgkQdGdkX
EVjMyEYvAPhRSm2zwzRaJl67BqcKx6CDrER2oq3zv0J9GHTzthZdaPL8SF9R9Zl4
b18jkTryfP2xrPmLKmhc16sq80THTuR0jfdX3dD0VSLjkCW8RINDFoRzhjHjG+TI
C9vftvaLdIYVPzdhp7Es4aP16Gbx5xW+x7cT4vIIP59jSr75l/4/wniaJmow6MuD
8E4PLpatt/8xwFti6KG2bBSUkTgAZ6FObgWA67wBKDLSRgDBF+qSXA0TmebTp+fG
lMQ3GB7yTJXeGufl/hYLUOvmPVXJOK5igZFlmhUH8Gef1bmOA+7XOiLPEcZE4C9G
QfHYVb1JzLXS/KdPnFITnCeVQVatObEemiDEu9VkJDbwtZ8Da9q/fdx1VYT8VzJb
oyc3+Fqa4QhwkTbmVfxiPDr+TSTUy3ubxlEQ+rwFUGEekWH63g3X+xIMZfLFDH3H
wE744kIGU7P/zSM6xT5yhZyDmh1yrurGvtzqb7Mkl4+vdheOTFYDilm/Qp/VqILe
ZPHAN47YoUBUwc6u4u2EefY87gVdfXXLHvHwZtaDs28EsSexCYy/gfzBJJ5MQxs7
GGUWRS/oPxWxQJm4d7upd6CuBZOi0xDAPJlzsco2vVuHY0MIppKfX5EztjSirXhF
PPEPC7Psdz0IGo7Cf8nkqwstKYxTlMUgT+sVfZf8rKXZxfdK8W7jY6blK9iZpqzL
u+Waml03v0xSYws6u1W/p0nYbpjmZEbBstFDiJFUyHXTi1NmvPDFICrfZ8KScZ1h
q3wA14PKnowaobpl+Z3Pcqfzh+Kqi258+o6XTMM7E4k4WJa3zB0E/SJ+9DAaYy6V
etLpcawHjdS1EoPHTdGA1OIJ2XKrB19JtLcBdayD+V7u28xrexiSc/Y3poGvqHYy
yNsl2oZ7NkYY4kr6twlGvphWIe/67VhO00toeX5iD4PuZLrTrWKZ8/M+2Pvcrdjv
N15snHx8NDBpyKZoM+F2j3yZj1KoYJvv64RRBqSAW/q3fhHtzGEdezv8G6abTc4o
PWbrddAqzqXGVv3udylDjqX6fooB6/dZGRP49VfJ1EUymI7KDAoFxQzo25q34/55
74Qqnig59j7oYkq18iSYYJrWcNHrC3gnmkk7XzGsppXCC4ql9Wph6IWJkQk1D1VW
DTXuSjq5AI1fQtszYR01gC+6arUVQfH/XszvMKcYYRDjVINP5h2Ub3EA0IRfzN0R
FZ76V8evApVnA1XTQyg/Oyf9wpVAsG1pANRPacQbahLAykTXXuUsqq2coD6Hf7lD
sDOdiFaMaEv4qIGIqOQJe16x059/9Feqk7adyH5oZJsu2YKJz8+Au9gMHmWdaE5J
F+RImDnp3YXoT8WDgKx58woh+ArYktw/BJccEc0tetWAtj25DTLAaV+TqepFrXmx
0SQX1ABKKZp/8IeOEOIrBxiMwGxpb8JbxZ83Ibhf0B51IawsqgDY9P/OjOKf2scc
olUzSk764NdfSDbSiwybO3lm6yR0Wh1SL4KgNmzgA2w6KcDYQMVsrzl/sOefPzap
YAaLF3A/jF5+LIzlGyre4rR/1u7aJNPobdEPFs7goDV1p3B0ZkUKQONv6XeQ3N46
jDaVc2QxXm92JjkfDJTQ72DyMCGZCSC0vEGo6465ffE/1Bvvh5cYzjwLlC7pp5jd
YS3DlvzrnPEx8NXOS9tOajLgSGqFHqAc4ocyq7JO18DWpWxyZV4RN4scc+N1q7f0
+E2T3z2lgDvLI9CPPm+0qpLKKydIkni0wbZSg4kgZFCyAtuS5L1nj9GxgeMt9BHM
lWzBpv297IhGwubmawJOz2VpN9d+5wUaGjCEOtG5ZTU6bJBlylpPftvrOOFP911a
LSKugJKI3dkSJg++KtO762eCI1TLg2ESbwuK14PNSpBCyz/0tT9hmPGhExwijuCv
lcsfe2tbsti8we//z4IuKLoicte50ydGSC9OJGJ9irHJ+V+qp2QiEyLT2fKdY9Fu
L48LiQ0567SxtSYb4N+Y2mM9n8qzMSSroXHBNOMgkbWF4VI9/W8AmZaQTqxwune3
oiVYe9AgFV4wtkLQuSzzI7RDymOCs8HXODzA3jzik0rmJ9UqQOprjKUUtfsuGD+e
qvJ1rapx9PzdhsHJuUYqkmEa6cwueZk5dO3BXKJUHPRYYKygkhhTie+4DgTcFgWF
v1OKwHDlONVGw2qF0xILlg9XaPkPJOvD1oGe3GUdADTuYQ3BRkanb0pyi37eBY/v
d5kfg5Pbc4OO852+GwRxnNWk+ei6xrR47HxHhWAUOy/eyLWGuB6XV9Dm/NhM7dL5
mrDkGU0p9xS21mEsUn6ZW7otGSHTfYpZ9SHnHV2mdlE0ft4vBb2UXrZKGfbZ6zUe
IM7LUp0MkjMzg1hsowMKLb1P2vISOUkxp87Sb/k8ox3b4inunVd8u11lkZvnORyJ
lmYYXy5U90TO2yws5MloR7mAnE+ZJcbzvUhHoLCMcNvWb88f8iYNpetyBRDH204j
PZUjVtXJPVeZ6dAY4ZUTU2Rj9QXP3APpFmNgKum2v2ZuQFd3F2c7vZFxMlm6qBPV
omVM+6UvKR7brv1l0MwmUj5zJyi6W46G4U48XQr7xNxuqt/hXWrI9rXDmF58zPqi
F2mf+rFo5LjLhGHZjUVWTU85DPb1HIIsMdo27RR9YDP90kyg8Hr7AGt09Ea+PYAK
64aXUBl+VWz0457OjLlEbWZEIUFmkapz8hEIn1Eq7tDwJZuU6/22QC8AlPgKvE8L
sRCs0VVyGfA8l4z6Z0y0WFslpDiRX6HN1Uf4DGc9mzrnVIJ9/jOscHO281Du8XT4
A9u4FwTWQFkJO6I06+8iHyTSbesDmdFgqeCvGzSqT/RsfgkPFP6hP12s7lA3IdbB
HYgA8sYfrkYHh8Ic4aiTAYFICEBrOBkIfqTvUCXGME9tPM/J5xEX5yPH5xT5G7/y
4A37LhM07kkhNVR2UA+ouIWsEggbvHmkq6lbiIrZXw2PEHvEfJ8/XVbQP29YRY7w
L4O+i76buSDZ+GCz0aLO6HvBWe0jMx57D3FYZ0qwEt+8SyAQEmNV6P4PnRtSbKo/
ls2q9k6Dojs+DfBciS6SdGkg08VlFTFrLodWJv9WAy8tl3WhTc0oUzF1JT9soMVt
sEmDbEmjtJW2izLFrQCazIgmp178mRVWX2WCHwTGVziTH0bmM39YVjb/d+g2VUew
egK0Wz4hcfmqum5gcZeARsFGzrs+RBurnqakMtZEXC26ZlzvPw336bQO6KhBdr7a
XQOwcGoWhwwOnxSCDpJhiErodjsDU6leH5zMvgz9f+zDU65TE1yZtYst18W+KomI
TQvXmU86ykkltR4vV7XCUPQMC49lxmL1nppyr1CN4+U038Sj1LAW8co95JitzZi8
M3Ypf8m02j15etiyqVzY8nMvTOV1FlniO1f5sg2TPNEo8C+8Ew/RhdEpPTZm+Wey
qSfwF6asAQycI5CNImETex0NPedrzvzbKZdWAbef0i0XUBJk4nPKfMyBi2Pb9bWu
xO3+mek/IcFY/0TUVT+GR4YZTomO72VL9Ca+VnmX6OAEIoIPXHMC94VDuoQ+HMat
ewMRmsxn69jPrPbnPWRkO3sfY7EnRk1f36RZAmMHJEn36O8CPfZQLnt3hvoJdOgO
w/qEWNXbLG6M5W42rE0WgcwZ2B3yPCbjbn3gcEYPJthL0oXu3GbMjgzUxK+aBPOd
BUpbH+U6tP50KjIx0ODkbsTjkNaFlE1z6cBjwYLkxfPql8hCqwES9Q9euNtYjgTt
8Wv6Z7H9R4pBwyQDndCv370MKITFstflHqxKDU92OG32Us68KdJurhfjVvS+G6Im
SqNKpLCMZjVert7rsogSnHCq03NliqRZUo3eflS3kkR8GVN0wa9jWdTpWLvrDuFn
2+sbRfdRNSCPgS5V2K3K4xfA74S5pIpUdqUf7DZ0MX8Ln/8o5vP8JHEoB1FUMIq3
3LaVQihr2e/iRE7SHFfWCkKc5CFptqB9RPj4h8FhUHv6Zl0gjtZpvtg+aYvsx9eM
QrpIVBt2nYGB1TMhTHYejNvvORDznvX56/xxM4oq+MLRUVVwUgLtFj/VYeRoCpzD
vY1cooPvIVsIKdA4inCuevg3vI+Lh4zBpznf+trIPByyngIfZ56ZVlOnG9gE2mfa
noWxUQrHqZONpJCRTE/FtiCxyu9ImGhUSBgiWTX9rDnrnqnl46ryAuS4IcWumggE
K6wz4QDAS0QZJnd76UvIGnXkaY/ghKAc3XEyqcvHKmf3ZFPQuNMzzWNp0FlmP3vN
8djYrFAnSo0NbcjT0IXlXrq0+3yAwN32i+zsMUZPFrIe8hdRnVYT98DZve/WHCIZ
bI7+U8lsyxqjr8fVN6L2/qIhgr2e1lKL3XLmIb3LdxIg4gqS4bdWCabCnjWo6/Wm
EUMOIFhdNwQIKBln7oo3hY+JQVI5Pl53OEcAM9y/+0luBY9nS9k2/51bXIk+4N7T
3vGCRz0us8auZr+sCRKovcUSa8qoNWUcqvq08n8cL7bmPSQ7yGb1UkoZSRa0vxA1
UO7u3x3mcxQK26fNz2l7U/rIVXU0vgZmEh2hB8qc0lyH3ScJf1Dju14ZHrDq8Ciq
5scbE4ZICdLx5cAdhpFib5a2HvmBaRmb/temaowUi4Mqd3CoHAHgkdVunJxfDYb3
8meVrDLGHais16aGBWJDrb9TG17NS+okOfLUuxhk48TYC/ekrL5B05i1ZMP1YtDi
uZSZ223C8WOsWBvb38CUeSxZksnxdrLFcl6YfVtqHjcro63UuAYjEUMs/UfEj+0A
fkQdNdKjeGTJoo625ZzA6Nhd2zKdvS6NCKFknscP4WiyKYU9akjFkMzIyBPgvrLa
k02ezsbe2Pwaib52ZA2ZPLrPiYfCnn1EdTlAdqOoNtIozhrv9ZSNFRt1uLuoiqu6
V+YIIJhA79lW2dPsn08q6w92K3ar35zVY3elnqL+lfJ2/M82grxtWdid/vRpkgpU
uZ2G00FIOp6m5o+KQCDgLHoB74DvhboNxJKqCdvmR7M9Qb0TLFz1caST/HM9Ol2S
BeUwEc13kYKczT5QRPGb5rmmdAXU99inAxVG3UN+MVz9v5jL2rxVZPol4KCPLSaD
sx+1OQ0ENY7epJ+wvQaXiGsPPC9WbTg7z+kT4XSd2Ijx9VmXewefHqJVV+WIzpNy
dbbpJo6rBoh7jNA9tab0sLgQ4LV0XkwX5+3J9ROk82QxE0pjic182YX5miANPUtN
3z6nvplX3+gUZxfkjf1wWyFyf+YM4sIRZ1ct3GkroB0ojoQ7octVahycqWBcz0vF
VuSQNK7UhI68wXQLiCsmGpCc73LPeRM0tztTyy2T8izWsEmWPQcEuZgDTH/pF7O6
zi+LRxyCdPOju8Pt/+5o5ytqzzuVu9hDvP61AJhHBAfnAmogx9ZyxF/DT41bJ72v
BLLQYz1jMAr0LirbWCxoAYxlYqaswOo8Ru3VZa1z8z6jQLyHq9OqQFUL2EvV3V2t
ogWdvpfO2JrTW/KlfnQGAEbRw5dnsdaLSZegJe06xPMYjCkqXNFkr1301zWidMKt
uLfX9mh3OO1d1wKWPm6f9BgtJN0X731rdJBT5egIWSNYIPO7Olfj3FCySvVSWHHf
oV8Tn67B9Ksq3Pe9ZYGBovJaWYUrzscMojTcJcLsFARhMs5N3csJN34wJXc7vnzu
mT5PtFSdfbt0tXoGUYeRLYzluKDqZ9nyTB8OyesE7FVuV+Vmo4wBRuqp4/nc9bUi
c9IP83lPOvsY3fkoA0ObQfRa7HheTRsXyB3HV3PlpTtdAAgU4JEuPSmCaq9hV/6C
ZvaCLVt/j1RfHd/T7pm/qoR8TVaxAa3BfOZNDs5gIyUv1qvUdyLWSSY8dyqoRxuD
VLz3yQqLTV1sddSD1ArE0VJhYsrejPL7rXqd+QQZENaRiKAAeowK26G1CVE7trY+
kHjD68SIqKHCTyJFqw8SgQGRkhdmUS6m5YTWMcWQqOM+xeCbFM0gES44/A/KgJw+
LN29yspUg2b0RPrEKvKWRTdTacSpEIpLsM4kfZYO8UyjU8Jc6VVghKqEf4ejhf4O
JYfp+B8Z+KPGpE+kjbgU3BP3whd+jYN2ZSjp4oqvPajEKy5JbcziWxR9cJoxNf2s
8sfmQZlDXzdd5XVMfRhIYV8TnhGPWM5LjsRvhbUrEMEFupDsHXo3byJPFbpXOmqt
3uxoWPf02rFCjoeJfGSo5sUgFmX/JKdVOiTpw8xEIaawRX/X2kyAa0UjzYOVj5aE
OZ3DCkO/n4ON/e1ibRETGn0coBgxHshoIZJCJhajKZ0w96vguJdVGsIeKhHJbO4L
pkfQftu36V1SVn+hGfrp9kKi3/M1/IoxRhvcpbwW/F2VViLLxlOWs7OlvpZz872i
7EpoWvnkO6KXL4Y60k6AOL9qleY9pAFilIY2q2wSg1U3JmcnDQBY8BoScqCTe8kS
AnRWIOj7yRhHhh0EyK7+K5J/+TIqtTzufGvVLGdeDGlL5K6tFdgE4mxMOaihuOor
f3XrBS9UVMYX6/IZS8CjmWeM3tHOh+hRalIJ4nODxL9MsvjtUjc4f3WOF/h5wJWD
xmrX61vTj/sE3G8MdXZGdUt8pX/lKpX+NqwsX8el6yMoxgG9Y+/yYtqjr24AwrIB
PZ0UpnpEN1gPBTCamVQd8Nf3XWvZ9IQ+Z1PMZOl/XJBJuWS/CCIB3gWsEZBJ0rgy
6G/eMyQgAR1fT1j7GfkTi5WWB7emeL/tbbohYt+lTtkGIZ4aV+4Fi/DD7ar/1Yph
JAzIhoV8hdxk4IP/gl2KbqiJWnahNR2FGzSTL9rl8gzoBBaNGx250YjBeOwQDgkL
rKniVSwHnLTOOJYPtFQhvU6BEkxVLDT6GWiwkr9mBLhhe8eSkIZxQdWVIRmYsLKP
0vCJq6cw518kWt6DWKYAvwUJKZN+3riRIMiubNmqOkIPDL9b9nSjKkDK3oe2zs6g
fcLR0W8AZLGq0mOyaOhsaiOwm/T+s+uvdtCyaMN/YpTq4zSbotrVNRjjQ/3W/3+b
Fu6isnhbVivFuidpXwOGzaJPVXpvlfTmLeKQpXP0iQVYhZqpdsqaiAROKod0iGJq
YLtzXMiEDusteBAaRLQe+uw85XNM7zYMrQCCYlAfsNYkdWEy+09mj1jZIayn+ihG
Ec3P6Cln0vVZEPAY02eLUkTeAO+7xX4szfQZhrh3mCXST/gqsDc5Lo3uYHWvDAJN
TgUN9CwdQ4On9tiy6vqhr20jRCpOqaauySfwphteaixbg7rjvv8Obha+wiwvpCJ+
E9xDDY2BRh7c/+ff/7YVVnzYbBk3JMBx9nkQX/yuufPAvXR3+U7cyxLMK95jlq53
qmJZJRpFYFg8BiZwiI2cX7XUycd/43TnXt2r6/uZxIOBbQPXXCmILhFDqTD7/9na
SyapUHxOUriSn6xV8ycyWRFltlGFLrRjqCiNN2NJMSPlVHY1NZkC51hM0EsiDsdo
FRfDAllqyRBSSz/wkAhrHHsULpMtsARc+XkmHWgw5u1+8fnU8v58h+aD8RxHzSjW
IY5uhjY3Bdriw+wFV/w0SEDL9CqYcn0GuEdEH6wJgy+MigYppVBMwqkyUpd4ASTl
PxiwmU+fXgtYFa42WmAGOuGYuN+Od8+i6w/i9OSoynHUHSVCu/1cjeZ13+u7DC1o
0euqEBxrJZXRDyFk1DGYRccEnlK1lMjGQ6JNmNccbU4kLJzp/p0ZLSw70COnAzDj
ca8+//99YvySzTzYX/k70LmAsK2wWQX9hd0UIA1Dc8Sq3SguHGzDrzvCRtX6IMJO
bld3FhvFVnG0P5tNdr8apbOuhFMckmThN9p6Uk7R+oEmMi2z2u9Fnuyf0FGYfrbB
8d8ew6ln7sbMdTySalYOgtMqx0VEErfVqEL0CIn5yVY71r57ErKkeCS5Qvaadqf0
EgdIfqIBxGT6EJmEkI//ARwP0SKFd3GnEaxOyzYRZU60IyUMclwGQXgEPm6yUulq
fJ6empmdCzGxt814ESpNCt0t195FpzV8ecq+4mHxX+stty5zy9lsYLzzklaGejkq
ES+NEqxw+yDV/rVNEcq4o72xJ/63yNYnxLDoeaOG6eZGixFzLwU+jMIRFWD+Ierm
s58avO+SFENuYm6YdPD/MqT3NVb0D7RZGf9WpPSzcM6rrbHB+Ypkqr3dkIab9T0C
/q3FYqmzjgJ5yvGFJp7SQrf5hg7iPy2eehMzjD+qS9ie+Z6Z9tsC+p+G22BJ/Ye7
l6OcsjacSxJdxkQrAyRocl0uSel+d5QUnjZIznNOYulbH6VuYDuOS9bW+He8Vokm
OKjV38etxurlUmI5FQazhqqg5pv/FiMQTnaMzZt7OxK4lZWF0y5DxkETRwelXRkG
DA/wwKdXiIR/Z2m+88EzGy4knhMxzBWBvkJuE12OrmVB38XmSYu5AxPE2AtRV1z1
wy5oisgCR1g7B6C/QOQgHAb3sypRXKL46tTew2bQ/NJeJ/rD5566xzmf18ZfDNUp
yFShsM79bC1ltqZgkVK71BcYvzQC7Z+LsIanUprqNExygf8C2v0TonLGPdbTdTTJ
9tCx/UtjZ7TPg7arFb7b0YhPK5b7eY4zIRTnR7Xe2ZO9sEmwWwnMahxMOBhuYbaV
h7P9Qb3rciQyw/x8ebQ//3oUhJmZxpgeKGyRNFgZi46nLj0MPn6Q6BkL5Ni1061f
eCV7e8SkgU5EUWHctVvVXD8mYChPfG6OPwtX5owMS7x7nSIsIj/h0/IkyEYrAJfN
UXs40RDUbYGtC0aAJ/10JusRNThk1RSaQGndKAK7C8NoVG/sTRKBlYpdRnrI2Fbn
mdjTd8++i/Jol2Prjt9KXaKrEkMVN1h9cMjY+r0+zHYLMum5M3P0IvsnoIsN/f1u
abDzWovn/q0vKe2PHmAIjWVb5+5YQS4FKcyMro8bfxAE66ACT444p8VwcqlF/gKP
6DtgHE1WXclKgonB3Qhkb1xYUWb95f2wH4tL3hyGQL7uFKpV8KsLXblcPNgMoX6N
0jvfVoGKCZIHVvN6y8DmcEYGsjHA4IUYUbC3Fm/SPZSoTJkaW+Izdf5YWZS7IQvz
b3AbmwrR9lONZklv8wk90uUzz4g9ikOTZxTh6YF32DylJjiXoPtAvBgoSO17wJl2
CAtGQsk+m6lfM2WOzovLo0XBn1hH+mImrKnKGtZmcjj4tnBb16tqs9reDqJpR2dY
LAluCbv5C4i4B7sTKr0EnwZrcGtu4qL47HdUbOfD/5rW4XCTAcR2V+hH7jYL7Rrk
FrHwUEY0MDvUkLgESXLIcQKfwnHkH7RvzQ6p/IkwYrmkzBW40kmNSncNg0Pb4THj
YsjdGQwMQVFzmX5xRhYy66xorCrUJk8OiDlGsYOL3iUwxZk2zxDpY3/IVfVeJxaL
mM6/BtDQiwswkbpxtOPSmzW0FDSE9hwy0ZLHsz66TSZKMXyGV9E7Rsz2yPeD6lNc
efJkxiiD4g/f82+hjQb+K4ZT7D4ZC0sLnCT6gYd5H7w/g2odS954eAxWZgMduZ52
DpkTyHWOnZydnXJiYjbMuqT7Xf64XXnRUuOu3pGEqrQd5WOzcdMr5ZnbZgwl0GuY
He9C06eYXvFAP5Im6/hKJfc+PP0EW9P0mKEkQRbWrHL5X5CUBIzPuDdWAUYsKCEk
4cY4bZrSfm9O6ZkMks2rQeiMgzurEZ9oerhqszYFrSN3i2qW/iBDjgsnl/h9rn5b
YrUs+/sCgsg6pZPQDvj24WH0h+hG3XOKxO+NUpoW65CCX0VuTAW+ZqQF1aq3/42U
/hLeSqE9QJucOYXw3VNtAhObU734eh+bXnw4m6Z5Ik3q8xTQHZ8cZIHrk9cB6/8i
ZVq60CvBuwNzKkC6xrRL6/ZKTXtjOyhYeatjMQiTC/DmkC4AYCeqwlde/LcrzlS3
O3yAnC1m4ejdUeIRmJjjvvJWoylIZQPdXgFMNRMykUgUYeqr/OnsvS8Lxq8+ul08
1CmtvSsgChXY9kjme1tWgTKzZFZx39jpbh+ty+0kFZLR9CtnHRXuzSqwMiexTK1n
H6vfVJKI1JpvtHawdrIrONW15l7TE3YVVAhfgi1CacrcUtyrozSUXnnFPpjKrfcM
3Y/nAeYmMbp4pjj2ME/w+JM7W601xNM+3BPa3+U/+v1UXi3vN479i6ingvLq3fVG
U1MaR4l/dN/VlYUMjwkt8K3pOIloW6FmpiZzvXaSm1FfMBrd3HAzX4sfZbmvBp9r
g8Vw/YbhgdF+h5P9sbsQnnFzOipPaN7UgjFArrppt75hfZaICpgFHN/AEq0p3ox8
QRDz9Bvq4z6Vpdpf4SLZNin+fZ32MY0H9w2xgG6sHLfdUvVXjPVzIynNy6so1Huo
p2vA6NmFE08k1YV1e9+D9TtezZIdBCFDsLlIsNPEhM9vlkkLBshNVxfYb8eaIsag
N0heuLnPBcaK/SjpyA2D9V7MYHpJSJXBNA0CC1ldhowaoMLMyt3d9Iq2gPlFZ8IJ
LplchlZF0czkXIPJkHmW/ILzBUAB/JHZW3B7qczaGCQhGdJ44p2fbUl1Qr3SxR3X
iQ7ErdX61QzQjSfs7AX/UoPYF68dX2glVfx8FiGFSpOmrmQwqK+S5Vue0JobvdGY
MHfylTq5ZtMeUi6ZokyeEyTH/k5pQj3GOV+BnH2xumSDLL+SFLR1ybWzhVsp8sxK
DLVebDQQmy9ccfxLR5nSXdWYoYod/izcrLjAAjztuMcB1xZ6yQ/9iQOWu2rZxCUB
yoqyrIoOhTMjRidRez0prYCZtqFtTGHgzr9lO0TICvpu+sWqbmkBxzmsT1Xyoa5X
iNwxYo24iRbQLRIeQX60kaBvRGn5gElTs0IA5OynP6JncWXty+wawVexQgtkEOkD
/S9NIVYp47f5taEELvZfNUdnp2l4usr3ncbvmYf+tugDTd61rwdi1uGdci3mLpxG
FHlpdM0sXkzU5He8DnKhmAnbw52UGNEY4tE1JRj/CZDtNOfsbRpqpiSS6KusNpT3
1NhIOPn756YcEz2WLUpmcxlZtEljXYj5i9t8JsOS62g4S7ak6xTNLao4KFc3/Vnt
GtjlaApm4b2xMRSlqFChE0/gkyw2PInfYn53zlYUBxHJOZBYo2/1zMRvHyVU3Z6m
a7LE3m2/6NZguYwvJlM+82PNt5PJB/rUtCxjVjP/SsJygIN69Sp62Ac5c4sOs852
OqExNwfaQOG9aZ1xFu/5+GMoniqTGoFJposcJmgR0EkpK/93wrGiukWnW/nZeX4d
7+STo6CNLkBi4DXy4PnVB574PPkXXQpMcjX6QJmoH9200m0tIOpklTcZkh2OAci0
kKiYvRdHCr1ed3dYc/MilX8i9UPlNtVFB4hj+fYfUqyQge2ObG+keS6P5cBRSNIA
XRuGW6g1v4mNqK4gV+q8Y0WtSv359hnccqLRVbWFzy8yjEhGFBIX1iquKEXm36vZ
8iu6ImoDwAhX2kbGwww9Tc/4j8gL7DT5+ThmL2Vd4k7UVj1CkIbHVbhAxVG6AuSY
gQ6CW14akIhQcwP+4XBbdCsH8D8jJBBTdC/u/zUtHE0e3amS5tvTGF1x86UmG9N1
ZUe5sfMarZT3RciRiZ3pdyeXwnY5uGPJKrYHkIQBar24KZVeaeFTOI4FsGd7EbSn
c+mqVy91tIPd/yIed5Li/Lo/oehsqKwjXx1CGhuPZfyLdSXWj8SUFmFU5R6R/bD8
9vPiOq+Mp8Y8a/41ABaXDZT7ZGtoiB+cK6PQyIqC8pfvGiyry1vuYd70f7gtfJ66
jDkkm1zOxfAhLgX+FxS11zl1bG5oXzzfamz5m2LRsfI/0eff+hJUt12m9+YQU9Zv
K8zEFJpUAaa3hNTk2fl6z6qQ5JCBrz5s9BnfmyDhiGRq0DEUWo9zxbMj+B2BImdJ
tHe18/CZfl7DQ74NnjH8xo2MrxJliQRjCuj3vzvdovad/eTNPCzTvgGCKRb3ja+i
DeRdLxQhLYUTR/1zbUhROlKZ157WWYPFzIfIfX9R5zWirTecOPLkHBUxcVwnMF8Z
zuLY6fH3Os5pq9aU0UCAn7Oe2O7YiKcpAfZVZ/tUsCUiuPldYxWaGV+eZbXzbr1X
/rA0c67TLwtGi6kFG3TbPuHTwFwrBZZjF8h7xCEprdj8BmAKLaCwb3TOxZBrQSaX
Q3c5pxBsPj+6i7zAwRWEKa2CIicgCggWU9CTYUhqiXZiIXM3lF3Gug7UBbUAni41
ZH3YMlAjv4FW4rSTuuLoZcFrdulYVhECXY4SgUEUZUrxJjI09K5uCKZ/5N+GzuOD
L7khjPz4wpm7OseGbMX5cEn/eG0cZBPxhRSTlECspnKzWpZnm3qoRdYb9DNENief
jy4xJ/4cc2iZa0MJZeiLFe4Iq4KSxcJLPZh+Z1yTMo7Mj+ol+n8uID4kLiXtrEd3
ptevIi7WoDs4avv7Cjdz+8U0kC1z0YYK8QwdfVgDtSir/oJmdWeDYonMScnLSBum
+4U++GmADz7zL/pYjTD/KuKaoN5Hx1QrlYLtIHnc6VSco/9Qcy+ZpZH3lV6KWtDV
P0Q05OiHfunySRxFnRKy3I8Ur4uCrLgo0TUZl9jLcR54xLsnuK5jbdhnErehYdMB
0YLm6VRh+/JdhWROlP303YajUE1l/LK0oEBmnyaB0FE0n3P1D0D55oECTZct35BD
d3yGLQjwEJuPPQY1IOhnT0y+xu7o8y7nRpuMwvux6pS/d2+rPrDxJ48LlDH6Rxhc
9BDoIUq7+kX2rlBd+YQ+UhqGeLVZUoP5m2u6xGDBYmuqK76mFOdZcMyDwjlVWIN5
1hLBkWrox0GWFvFDBTmPtreH9jRhMmU/xNjZ4cVPNUHWEDtfmu4MuDxRGdCx710D
85kKRfXrR0PsFGBByahG0Su25ytgyWrJpt2/3tdVjCCI0whr61w/1AdRluj6fLNu
4gK3uWv6qjeqA0ct5ReouqkYeRRoeH7qKo4Q5WvBtOk/FGuTHQYpHQSkkoiuhTq5
Fv73SC57hfLLbjS3X1q0K9XCFiJOowB+l924sI4YtncRRohNUGMVh+3Z9bcvcSMK
J6ARgs38ArFDwv3iWvO9i1nI6LnK+5MaVSf2bAfHEma/5eu+kz/TL3Q4aupke96g
FJwkr9QVg8uE4Vn53+2N+uvfvq7w7tz55WXz4wOq7Y47PSdEr0GT1bvHh0fuhyyn
FGrunXVk+lrqN1X1nFzRHN6Ycu1NUgoiyEhZoXSA0niGGNGqebGI/VuOytK2i0DC
DKvELfgCyfYamSjWVSkR4yXoT3AfCpECJjhHgfOnkee63V/CcPt/WVDW7rO5kHVB
6pcvaG0rtp6JrSXXJ+xLUZw2/7se7NZCb8rCY7w9C0tTTHIP2aaAdd4VTLrj6d0G
r8B5P0IkzsXJwE1CWMRimelOXbWBdQheE6B+ZrZ3mgo8AzedJVvlz0Pe7eNgXAVD
vl0mdRltT90+dDSI5nMtlhlgjVNDU3G0z5cP97iDReuHF5+W5OLhPrOpyL40BN/H
f11GVaKK9mV2lWX/Ph9eWqc5cOJdtG+MYIFmbDpLw2dWRPyYc/fsxgaw8MWyq4nV
Mdv8zfAAF0bq3a9+hrMCrvho6CyI0xIsbmgYJxQzxcaAZUXL4ODiMAO0bgId43mE
yU0qayjG2q2NUPb+mGvBlrzxPU0TiZTyQEZ1c+FdOerDgBN91KWGQpzn0B+AjbOO
BL7U+pvKysd9V2hvECmASX0kdRKM/r6CqSQ0l4CX927uRO+I7zuqA29RBe9VU6/C
rx+TDI254IIZ/S0QJyiMY0KFt8xYn2TddgQ+1roOB1hNwQfl8HlyouA2ZiA/kbLZ
jhlDdXKG+RiIQB1vh1eCXMz551oDhY/bU266c0ApI632BpURkk7vEB87s1m1qHge
Nk4kcB5eY2mkr4kwogHRv8UC4J3TTkKYQ18xpSnLEZkTFZ4pQ86lomHohANJqsBr
WZeogXNiJfTTq4/hvKt+15mN5v6feVlO+CxMBkP0yCuk/rhQGXo8z9v+qsD9UUyI
hSooUZpErZpNKSpVFzoJXpLsWYTWLbhka7cTf5rzdg0JOlxuUxG4fznlsoa6bad2
bqCNHwxLY3v6ZG90AQQkKmslzVkkg0fWUsbIbdAvqff+kdAcwAqmfrv+YaQgVm7x
MiEMoKhAOujPyckDbxqtBgLEMb0Ct9QoJgESQhOY3LGhobR/6BsR68uiJ4iMB5wW
0drToa284rGKE2UgTC5RokBa/2g4NRVtSte6zBW+D7eFScTJlpvYeaNexaL9XXMM
gIxQ6tjR9Ebg7HV0nn3fR/hrhKuBeMYOUEfoO9y9+fp88PJsvF5sw52jWyJUB4iZ
NgJDRNldYVWuM9w6TIs9udKQk5JKi91oDtGG8W9jJf/EWBDwkRlgSQRR2d4GRbwR
0B8KL9F4V4my6IGrRndzXTcVxy12a8GHSBWMIN19kX6BAjgUK8SZKogqEBeo4+GW
xypnqktdusWuP/HchsbGvoFovBavacX8dBmva/QRiLBB5F1G/GR5ZJ2lcXn9Od0f
TiCGIkvaJdAPi169n/0uKfCw+GUHGkzhH67y2T+TH8KYBQEwuOo6xIv5927fsNka
i0p7p0lh/aghYnzpW7Gr5iX5YuigSlYpzRlAJwVQ5bzv/8ezfVfh55EjbhMSo+a3
CBEtIq5IYG/rhxc0f89LET20mrDOg4akl7eWNUYC+qul9LOAEKlAvZOBMblYofu8
dy6AQjfNSNE4UgjwUxeXs0pnuM68i7C1vawn6vcVC0rhBbxKH+3JRZAtutQ4HHws
a2EyJIPEfVHzMBqbHQBYI4N8tPdYRtB1GMGqsqyJCmKVeM7JiYXEMJIiUmQuc3hk
oTpb7llJjTQpSf/hK/kIJNiFHnRcYs8HDsPqEaJlqqALT3MT2rMbHtroeVselrZd
7gW8VbzRcnj5pVQ1FN+1XP2QMJyIsAG3FTcDA6Cy4EJWMUtKO+FUkMeKh8cPpJTN
ZtzGhUOpwwLXNnpDlSfDRz9r8D582spqdfecuT/tD7818/D2JhRMYwhCA+w20KJ+
7PSYDSh7RQKrdEip7VIMoP72qIAwz8aoJvtG9kzFDBORXp6/nLgj9uo5mM9lD3w5
PNLUXTmULBiQhSH5KZr7p5nr4jCipO4O9y36cu0kJcno6X93h5SDstoTpuCseTc0
t9KVwhOd/h/YpTf4ZnTqTgh80pJHGxt8LAY4WD8FYjix/dDOJN8N4d0jumCTn4Hg
+lxtAzOhRCCM5rczH9M5Lr9Irx2g21X5EkvONOEqnYRH4HUOePtxw/AWBZUz63l+
IzyFX3lsILhtDgAgnVe06HAw74S9t+58qukFmhFeeGPz4IniABVb31YETpHAZw2e
O4BFfFmiFA+H2OYXiRwT6887/OIivOjl2St4Dgy3wbcPhYXCc4zBbyLVf098Xdi0
UnoAguMUQhKMyTE9/bGq0LsA2eKlmuKFY6ok7aNMlDd1p0aBRjB5AqXO8xHqVeQp
hVrSpfxzFCI8rzGf2MWnQQU4lE7om52zb0GjBpAqxnldRPkhcFXZktjxHdeTYj68
aVa8DBtPVwVrl0EIWpriRXuLnheOxjPAIAWhJbvtM1kTX4kOz2fMDKJg9xobI5OM
rNQq0FNu3G9wFWoiOSc/q/W/Zu1Mvr8+JBZF2Q/U5utqCOrVHGLmNDAdsdd5eAB4
ypqMgGxuJzTl5BsCUQMwdY6QCxiy6khS4dKB/Bf9MJIRkhPLahsB/Ij98Ucpp1Th
+odjb6bsehRF/qB1/49NA1sUXi4CsjS4qzSKHLZHCQens/sYirg3HUOeLnej2fTG
iyuuCbIXdwh3iPQ3OulckEAmruPDIUuLiSRYPCflDOlbdQ/xxpnWlRWaxtFjctMM
guI3QZEc43PqtAiBPORsmF7TbvS4flu6Cmt26chHGqiPSRh3jBblXFcR1BJN/J9n
ce/UJ4clWw1GHJ45zTnUFHDvc8PDO14LP5x9QEwp8xyUzd0hRzbDfL64Ix1xAwqM
L19SZ9FMfTRXyjHMOeUhuw==
`pragma protect end_protected
