// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:07 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H8vXzxeJy/3jNyvKAaNHLg5ffsqCipDgAYRzk/xMc2ganHE1Dzg8MAMBVgT/tfr0
N8GqP0kpzsdOExMyC+vArFT3qx7o6V7OxRTlGt8R3m1d6gYekD8ajVtFuwSWdEps
Olt/dvay9CiEfrrZVq6yYuU7NSA+q4lDbcF72V2uxCg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29216)
6CNYmPo0prGgeA+ihBYdjWR9B7HZjVK5kohNhKr8JSPNoMQVVhXHLj9wmdzyihG/
VETZR0JkgiCgPbjrNf4lgi0/dZMbiHFwe4jOyPpiPz7i6yNDULLBhOHFFqFiDGpQ
a7uNpmbLk9nV045IDSVcTQvcABPmymIe4rFcF0IcdhouVj4Wn7BFKcCipn2AU7yQ
JuJTjdO3Bnld2h2FC+mS2Zkmpmrunr1+eMNdWcT+FF9FJjMM1Bzf83/OgbZ2IWnE
okWSfcJgFSCy18N9S8hMuqjgG/BY2t+ruuS+zetcCEC/Nw0X7pHdhinFzl2UiYKo
8H/oGk+zJbgPW84HbOgabr2ZOmu+KYPoNodsksXfd1kXICjt62OH3wSCxQILp3GP
jb8LWCrYa2Hup22YXGVDov34jeXACWAX2wOSA9otZ7I63mkOqqmJIj6olAd4Kaob
ZVhPbDg6FQTyuQHoIcj89lyKiaqLMN3bCf+xubCUv3bliOj8O2pBq+hZ9SIMqG0+
T62C/Zd4GjFBq2kL1oATywMYyejrp1tFCDSudmRHGvBEshfnXQUNYcF2X//8Jzgj
lgmbsTZBIIXN0tKIa32ctDiMMHwSK7RZLnTnQhL6C4eEPZjF1CDUBfZI33NtqF7t
jNvU/LUr/FWt4+W6onzZErbNjlIef2pjb4n5KXOV1yMOFG/xTM8Y853ikmtf8hZt
NoY6EJdQkFoOivm7iQ8ISomHoqUwuOqT1r1aN4zu9vqS7qJj0ecSWYRoIMsVSFH9
34Qm2VBEVwFK1EVmfw1Lp1YJ7duoiPsmP1y6/t3unQ7TsHV1HbYL+8HGBMs92O/i
+EJrdzu7YOgvAEFRcBX0o4QPT4f/3ItSzZeR3xNC6+A+6eiqYaeOmRfb6poGS1Kr
DT3sBM195sZkigGCB9UGUqlWl9SaO8jwCCHIWi3V3xVOSkhTCWfEhNImGX9HzXoX
K0gbGB0/8e+XLxgY2wjUm/e4360bkQAgTxVvBnWhIdOb6OmD5wk1fVYEE93CJFjN
k0fW4rC8k9IaE+LNsYjgai6O5JPXOjPPCuNu5DImlIKQOIZcOU9YxYD4mcQERuYQ
EsDlCr6W2X5WBf2z05Xiw9Ez22+O05vZcplUBTCzr5kNpZTSoYrssueGqz94Mt1M
Mjbx1fNd/8rUznWbwmmXK7bQ95BtlpPIzuk8k6heBpcebt9qfm64OZdhZWv8dl9g
oewf3DysjeTmybJ6SnceWnUn9dilNgciAr+rk4Dwo3CHnERjXuN00hGoGdVH+em3
nDk8zqR1Zk3EtM+lOmMNwt8scTtIX5UqQXEAiAJ13T195qLigEJOKSAuJln7pllL
wvfYjnhkfbCyYQ6/wsK2V6fAg0cqq7jwvIGg+XhfOq3onsuoXJKxqXHJPWYCkWun
WGN99+0AMtCQjQoDuXmFGjVTrU/MTOP2dLm+Ov+a9jxP7gNi7nVwTCTYQaPYXsJN
tK2ebTaKnMH+rxzzkRhoDTD7i8KlJAFXNTXaQCU6O5O32uIWpyAS0El6ljIqzz1j
Ly0EzDbV++TspvYn8oTabGb0npPZ6rAQaZDtebXEC+FXA9EIByS3kGDNCux9JddZ
wIRFBNkVlPVHCXIN5zTf0Zx7MAObjkEUImDdvoeSmpJjcYprPSsg///18IORPd+M
sSIMuEvcyH9WxE2XACMB/WO7jWL/OGQzRdNZQDKfmOAjfT9umtqjK5uZZHdPp7F+
Bfedr27/olBJi/WlDbkwvIzLelb2KOfCO4ApXI9skr7Gyqdk3a0VVROfe2X14Y7k
Vx3QjDF1CZjyBasz/EvCIlcDw7Htt2DaGTiNVCntuyM+SZDa/jr2Oq5rSSejz5yN
SnONhYYcYbNSp0qqR/smbK00PzBEbO/Rj8hGCgdFSl2Jqwj+lyZ2CO+mMpwHb4wW
S34pACOFATscpsv/LgM8g+M0gLruRvaAvqRRkU+ul+J42gWa5PuW89af7hAY+ad2
Sd8w2E9rBUQA1fHfYYi88QU1lTy9gHJt87KIqjziY32eGs9hX1MJ5fxpjRnjqVll
5vtrEfpKsRYPFe0gUDKpqUsLhBY/AVtMI86orI871lxJUM74P2Gesz8wqJuYKPXK
NKz74O2O6HYcjjBFzECs/e/IMRY57zeRbZyHPinvzgFXsvp64R7ZFmC0LkLEJAV/
VDX1aRSDd/Uk5zLC9H3TGplquMR3C65MqpXTCicodMTDWkPFNywnHBl/ICMNnypF
IvWWVwYIE8LdMpmfPcrLq4Ztjd0dxosID1wO6sePIDQca3D+i10UyBLKS79NXP1s
r2bE1aeVD93ufgcyW22XSOSFGn8JwBfRNE8gt5SQB1OioISLEf+iXRwLrMjE3bdZ
1p4z2SCZym3GmWcKJ5F58n/VgF3BKptRvVMDpqJ+O6vQvkF9FtNT5/XSv6lhwpku
AsQ+PIV+4BiWwSiUvFjvaD0XRfZY3WtNQv1Mo0fQaDDy3wjHNrQMItV4K8XLVxas
fnkKeFh1afXKAx2NpQvVXCIVeGv9qk99z1Y8OvTUGXuCXGz8Uwh9klk7quZE+7ZL
C3CkttX4rK+DGFPBMEM1O3whQ5thTx4upFdIrymGv2/nXOC63AGXb0OjGtbTkPx8
SHwzi3zfz2TjF0DM3MUQwvC68svn+vPFQiNgf0meRduPvNnHWF9zcAVGZ7frkhZ6
dKkK1HANpxl/2eZX11PR679ntAfGckDsdN3SJ8KPgbEiUZtMrT1D4vP2nr3X10l9
TCGCdyb7vGnEE64ae2k4JJvq3PdlxgbaYe/Lt0mzAq1gRNsGD7eBlrAAzl2naDXv
n+PwKZL72qC4fFtEjRyQiUVybpCFOi8dUYx4PcGHtHCOtkLIdlp1omdHBkrnjMWZ
2h+8EQrVcmNhtZk4Dh1IYDyEWAI4W6cSmV6+gy59YTl+mNEFj2D08kZUSeUxvqZZ
MND9DD+MnVb5/Ff2SyRAucXYHvBPs6QJyWStE0bBU6emk0z9GGpkjiJ4F0n+LEvs
f9A63nok6FXe4mdA1p2MWzvBTMLfkoFk6FGS/VEvJeSqOcgD6qa2Vqu6pmuIntQa
qZ9yuEyG4AGJrgLP9fDqQpJAont1oEnQhT95TsgGgav0cynWjYHZLA4cdEqOuZlY
EGypUR4JXVZyhRXqp/wdXghJaVUlw9w3cllc1+cNFDKIcVskkjc3++R+OAGuZSKj
sY5h+voqRR0ak5izfTG0cxNZbxEhfT3cryUef0JHmXDG2PJFLyh+1Q05Yw6gXGav
HVyiVZYtgG+TAgVztbMZJuuj7BQL9v2o+RpnmKtyeqLn5y9k6EsGN3b4kTMXzEIG
bhU8U0vp3/81txo63tB2sYLL4VVBPcNdgvbKptBQaN89oF88ass27dRy/Te1Xstb
tI0wutSx+IU4Z6QJ7aofztJi5a2rNNjegqvqyVbyE8+vHcLQZNxx+nJAItSFSIjN
T93lZX71Jh6oOGUQShwZhG4iUY+R+N7z4s4Vb2OKOuy7R1qAdADsBvfr5mQKijOQ
P6PV2JZli1sI87N9fynzvkcrJES9hXX/jRoVHgQmw+hD+N12QrNhws71aFyoq3/S
ScOD7biMqbuG9obSqxUmbF1/hfDrJswpmLkDtRtWVR/irZxyPFoHaxJ9AowAy9aG
H8qMHo6YZFN0crJMVv6gb4yRnt8shV6mp4kuiJu2S5RJzxWCDLqObKIYPlctArER
WYm9Dt7jhgyYBC3E5Zoma9g3wMGnGUA59zUpC16NlIifLk9PFGBbk43V72ui9/4w
k/eUc+vFuoZZeBXHC1fDhJbLWTY/qOs0/S0KIYTf9YiQcb/Y926p3ii8aGMZ2FGs
NTaUl7j/rTDbP3oFqLrpbuvnJhQEnx2xmUs77KBG0o7uX707Xb3rnbIShMBzRMJH
SlbhL9fiZGQdIXxajBX4K3oW3loKkw7XIVVSLnnnaZRKda2iHLpDxGHVuIspc59N
QPTT3sJw2zsEbyWqlSa/mhGFoj0xR3pBQC1zD7NBPLCv0B6nMy8J1rBc0V+3vmGC
9+QO1OQaZF22JL6ne3nN0w+uog2jTZdQsN27HodEpqx6osFdF+qtT3k5IldLwIkg
th9zeV4qO5znb9o5u/bYoF2opO2VWtIuCEqLEK8k1ttO25FWfpSmzF4Bmr0re8rK
YhK22Dnfv/ul52wNmqeKsApYj4WnI2nzN1HEEUcGQW6unM9B2Jx4XWrDHOwx33B5
Gs1MwSmQNbb/1YETlWT5Nn1ycATRWTv8yoS+pSm8oO7uAaSklEuz65icQhQ4hKB6
H5mzf6nNPTcDVeLXzEG62Dl5yZoXH/8XQcwjYkB/sZaYtAu9jcWYTbNquqSXi0aT
IIaP/Kr9CPtfAg/nSkwNX1z04bykHtwQZCt9YO7tJc/0mtI1pgj8/JchwmhF87Tt
NltMc9kWC355s1uuoRP89dDB6+H94L1sn2ItPev8hgws5ML+iKf07b9uA1PC8tBQ
i+FKXa0aYnNwiIUgrv6j+Xju+7l2YXrPwV0D9XRuzqzL8bZM++qtR3aakxnzGMnK
d5Vwi95ITqixPhCZie0cDSCeNX2EyMSMkMtd1yvO1b/Y1Dl3QSTT7jmwZwYIyR2f
5EYfPVgptiuITFHl6bjlMU7cWx8c9ozJrQg2In0yfOrvtsX9Th0nc7ImFDMJGFji
UrUk2XKWRTvLjltNqKFSseTtVgo1H4ptIHMhpWE7Mqc3GAfIdyXhFYxRmiWqFG3p
PaCBu3c6h8lgFJhP/f0EK7MPv5yba2XNNhFNmUDI3MMpsHYemeJZepRWgkNWC4nc
BlXQVy9jwLwZGATDx+NoTA9jDQt+VaWbrbhPk3iRbWtUIvyiyFkjFDKIjgdzIvpG
afIW+m5kZ37fif95e/pKMiX3JyDFfhL1njG8gnRQlYvPCvjM6x+rsVPtBDMtbB0+
TsDHBZY1/dSefLwAN2wPK7Ik0h0t68oyhe64howyHt456Z2jPupKnsQTGnDhGE2K
QT/slCl9osW3Ah5LD4b6Ycq8ukYAPnrkOK9mT20DJcHeyTCC77DGvWaQADEHPseS
LP4ffMoVE0IMdy1m2R8pVNFB8vhILQOBlh+Vbjtkxw9TC688BVPgtxBppG/wmwAX
cZRJjMwE6oY1P5EdkqTPD7j7qIGb/Vu6bYKI81dA+XjNQ0jesQ5OYWUnvcnCoKet
UsA9RRK82ox7PkJIbV8kzkvnMMiEZcSwuInclYVcBclVbT8i37TKYsYLshwOxKMh
BxVcJXU5wZ6MPKdEvU5r6lq8Xptnnj9wMUhxwmfCyJsMfjzVRU9OwIMXForT4hBH
x/jle/YrAj1Av/y32Cu/+gnK7lpX4AnQ0w1Hcc+4lpJFSyOr+jBoMeJqyF1KSa8E
Noax/P7NuyRDfDE/cPRfOfgCsOpWONQvtSUSBTgKhsLDwhVeOAMs55LswDK5W3kI
P0juBS0mwDfBXgoxEl7ULnChu4vdfseJMVyELGW86A3bdbQTBjjPhujYll8TH5kK
AdEmjddzCoosRJ0RQwheQXiXFPp8a/vxT56m2MJXxlR5xNkQiepwLIVtskyIFd8v
f99W11T4XC+KS99Ljum91J060Xc3UcaPuS3q8Ot380O/mMWk0+6mpl8f4vJBxixe
a1dvK6iwvza4dqRRITizic/+8toW9IUDnmghnD2aGAMx3lmg1G/qit/4MnQF2oPY
mHiM4eKEHo8uoEKAZZ6E6GCiY7382LGTEGEQQrgPC3/3Od8OuHyxZJMOnORTJjU9
icRbe4NDzhwNFshr6CN9pDSZgbJ8GlLbnZHRv986sszJ4bhjR3bncz5cmb8JSJw8
gNWA8cbYVzgVELs96lSu5BPMa9qfdboj3ZymXa6cDS9HxiAAs4+Sg3TJrU+eN+4I
quGfPFPQfJLG5irliEaWc2ibypxCTONmo2UdrKbWmCLp1x27mCx/8UzcBG3fGgqV
G/lcoJreyaWAALzaKWLxoIqOPJjaaPqqPkpeX+1dc1EjKO6w8XwMk8xVWJniuKKT
PxcBjYjcsVnlqW9itegr8yKcM3lB+pN8AWZnKDp7NKpwgDnL+b3wodO/OUTW8LYr
9sxdZW4g1c6UAMOr0Yd5Jaf/HfvW/F+qgMXWseup3V+fbrCpw3YI0OaZ4hN/+rg0
DtNfdimKQZyXF4/EvscijNyLiNxstHyi0EZjchlSTDbAvX8a5VEZMhBx4j+Bl1BA
/M5J30tH6wPZSMtcuZyd0s8DAEQbn6KaNfJ2oXNCsiImFCUz2epSDh56iBmyFlR3
Q0iCPVJUiB/Ea/dLWtxN7YhAjLhHHwaLxbtBqY07Ix7QWrohlYpaWUVpnfrCIJNP
y0BtyIrHzfYs44dnRtTwG/sVz+mrm5OMgD+1+E8tAeCjZ/MZU4WCL4KaCZ2/HWjz
2Qy5L7EFJhW/wr2dpeyaolcGngIbwnteFCmWfhkC3P+ERimyBuR/7QbI/g+UUyIJ
cFLJc03fpEHzeWS7x3lOxezX9+o9TQC22T/7csKYpPkXuUiOxSnuySlre8TMLoZT
vLxFNlTBQFQoMKH6wke0haw2h4ISBBb9ZoZMZgYmvxMadixXPDyR6tetEDBV2qrv
ppWd08GFIvgMjpW/JsW+h1NL+t3Cuq7UkfZrQVDSa4+J3t/SBWjFLrJbpA8+5dm4
xef6xrVFwdSLI+OYcV7bnbTiWbGVj+XidPGE2iVKZs5ACybkWRI7xk/k4+2+UXKB
NHcESxrovNdxsgyB5F+rQaF4SSqW8OE96K9D5mNQdK3C9Um4Gk7uoTYKt1r7pVMX
AZHL5PoBULK0u3YkALlwRjBfE4ovTi7smze29ybVjpNeusVTHEs6B+xDir8mesUm
7XDcvTBzWBJu0dOUhh1QLfMJ9mh34gITkIEdc2dl9JhtNIyruCmdT6hwgpBHABgt
gKBo0h/Aj9GAoFChtG4i01grETR4DN1rVTKJkHEtwNUh78PvLOv9vN1GHusWclyg
OJGboqa2/qXowI7mtLElPDhO+DDKPwcDVpPPdPZNEHrymWbiKSYOH7THKHMHwPSR
MLTLzUJU3OPeaTMmxD+8Eolw5ZBKUQz65EEqRoOMQTXcNTfXy4I+NdV4N5ABCUv5
+IG5dCibfoUX+EVMG1oFF39MdbT+zsGzhpIb0la1QIHecsI6W6ciF8NkoFSmEyco
XP9UEqE4vwWHrcXmQ372hZg89h9OZGrK/jM8ulrloLIzLFo/1soyYeVgFIIjl4RQ
TwEWFsXlPvzewLTEa6XaPHmuFkkG875FlVyM/BCC919BCcZRi9ulpsuMtBWMMFPK
EtFyMRpi0tWxNNmsu6x+3+Vvpt+UHurXsfSl5I705yDfBaF/9z9NhuvkCizxd+0b
odQWyLysW5uaEFhHDpri7i+Xb3Pvx0oVveUNUtlL0eYO9Jd4VNgBdxjE6P2m+cuT
yVOUOWpdBt6ZuhmSvL2UO86/6V6n8QnfwPWtqxjErf+xBKoZL0K/rItlqq2efk5X
w8QiTfThawaXZ+wGZjZuqia1DIw/uJlQsGes+CVXbqtTWK5ikNrUDeJkQ1DddGAP
RRcfynDf2EeV9f3Nzfd55Y8awpXH320tfgODrJ+gVxuy7vcN2wdC5wiEZ5F6ecaQ
aL8H7yd02X32qtbA+Z46VXosZZ/Uo1uo9GecUj9cOmyLOxaHxA8BBO2ACaY1Zynj
WgGZbiA/MtsKKNmART+4yw4OwMOrWshaPhdNYq2fdCTlKLBBwnh/mnrXJgV3TQ1U
ml6PHTEG7X/aAqL4YLdR+TGal97W3Rz+GCDWbvmcBZbNIPJ5+N3H5kjdlkIbuUMS
dp7lU32o5HAKoqgpyBDcEIrs7abbWfpJ1ELd3LGZsYf5ggKWnTpHIfHbDr8RtVU4
oreSY9fmBuJU57vDIX8FouFGiKwKyiMFTwb068Q0kUpNgP48jyTE0E7Du4gwyTqr
TE6z9/1w+EhY1x6jKAMnA5GOdCph1YgWwXTMMpxhaawhk6ssxaLOCNUmwPZi+9z8
6zeByw2jnZry+RTnSdypCkmI4/1Dax4lxXPYEMLl4Ylc6eyN/YwWn1IupSTR5B4v
vcG6cuHUtrDHE1oylwAVxwkTqbfk+xg7wSMilXiKdXP8a/c40yA0AwNQZQgU3PNc
SSYinqM//YqeiAQtfazD2s9GE0ciZzWvqMazJrIPtRTFlGcDy+1fFSgFwdafPHdy
UK38GzcTbzb8n9p26sFJUjRqjQTlXv2aQ5ZLhGvv9p4lSPQw3QgoXRxIdB4bCdlH
0sQTB6hNbrTfH7DUWaXqkuwRT81WF8mya2SsAoJePPXOYc/1jfCGa4Q31FYVGJu/
1rjHkJn0ZQlURIDZwsN7CQ3I1WcqN7nsPZI0y/cXBjn4MTXX/cvVAe9WdURHUgLt
S0cRpaSoIGcOC8Xg7/VOaIyEo/kUq56WWAidBAB1b+F6D3XksEjvvX/xuBHHNSTC
p87Xjsfnjoi06VW0gRxniCAJ9jTHYp6ZoA88mjDRcP0hJqOG9DbGMK5FEqfgadJ1
dJucOCTacqGr1yoyl9sp1TGFMd8T4nMsdR7CxDWpbqHDzELTekXEZfUHFYPFsssR
aTpvkdnTdNEwcUX/UaqprZDUDhgYmopGOe8yh2RoZRI8xIVk/ssyw1Wa2u8c7a3N
QO8OWvuRqTK66Zl0QwGuSZzZAdSZSGFLC8msnHtXdC6fVikp6bYqCT6QQVdj4iwI
04VkhnrhuoH+eCWgaOZ//sV6I/LNQvNn+W2DhBzLBYL2K+S2h8I45E8aDUoM7u2Y
vIuQzKwp0bOCeszsVpCmKohj7PXNKt9MtLoLarT5b+RrwIMZOHYExvPlzPT4Hlxt
HWt5RTzr4JIoQdg1B2ExtoIe4zB6f3WqnU07u0lwB2CcAVwArh/2U65pFK/55DoG
GxjU5pWGHkw5k/ixMntm12crw3l5OHGMz8OydIV/Ix780Xjpt+uGSjCndpF2Ild/
ah5l1HWZCvHBHLtS+gDZ0/jW/+eL4+Sy4BLuvCVJcEttlCyb/Bqel5DkSvbdW5Q4
scFIX2OqPX0zQ1x7eJi+vM+vsuvxxIBnbVbDUw/AWFNs1tACiQ10vgHyJcE11YUF
maLKL2D6OJRTqFm53mhYnGapvvZdP6fD8YWUDu6MqkJF0jkEQcDRoDuo+4pfSdug
hP8pMUHfjGCuFg6cMAhCuO0+5yuvATimt3ym277voX/SdJ4Pe6YcnL1merwGiG6Q
IyGLsJ1WMC9sRb9+++vhaEBDyNevRYz4TcoCuaPIiOKaXZwVqcxn/531Nssr7lq/
RtOx/QMHmvxLbE8O/K0RU+IMu4fTOpw7V7qdZOdPmTmvXtNWIqd++ucm2l4PzHpk
xU31XP351UJ+n+afaLuhaWYEN12W8Wq7VWeKVaGm3/p+RMU+CcvBcLRxf7sz45Rf
3YHoUmVT/QAjnd7E6Jpk7FitPFIi7BmqmHqaX8wYIdOr7quygw+dpFj8xOlqDMRf
9KiS5xiPOzNZfiNjIGR4WnhNxzk4LhKS2okydYcXFCH07XwexBQnn+m73xNUujE9
Ntg1b/iSYSnv5ZOp/meAk0OPYNHb3dil39cvMo0CKNWdXUOlENFv3X7mUt2FfHD7
91+r0b34j9LYqXxMEJuGHWl66VoUu86K9wrFSsXDhaXWYVq245IjirQlmGT3BE5/
uL7EGQyQysI6y1jLW566YAHTasHJQYyF+eYHId4x2hpmvRKUXLQNAtl0ihrVYoqJ
2r+KQO6fwHvLIBDqZaQKnZ/Q7RI1NyGCBSP0bW7+rOLhjmTqRryv9eY8eh4CSkkZ
VvrdthUQHSanTI4u6KW/tZ/hiMTomaESXbsVx9SK/2H+tfq5HEU5hih742bfXjUA
aeAj6QwLGwgzjxYaWpXvjBSAiJEtBFKijw5XLJJubr3ZMN9eZZKNYpKdPgpCNR9O
HFjzQIjIHQIKBBdk7q3Xv8B09/w4zkaB5TBGnIwRSkvU8TfS9fzmsWAEILDlznqi
qv2VlX0WngTMSj5umCNnxtbI13exgfIDgRKI0HsQTfZiJNW7VpFBf6xjD0UNwKC9
K+zyeZxnPmavB8vd3tOd2joZt3GTFu1ukJx9nVZqvalL9qGf3FonGztXg2OReYib
XNsr6g5cMjHoC5/71bK8Is84IE2/1OBCDoxJVVSHtobyKJCSf7M/uwQMX9DGzoq+
A0NSMimTB4snNzgGgn6fFhM1l9YgFXmocFTsTpIg5SP4lZ8dA8+TkmzheXBbNLSz
sgq5zbrWflD5PoOt0xLpyjsyoT12MD+xIzRY4DUOmxgjWgukL22CkAk2kslTWRhD
PZ22FVQb//wm1RXlfrs2b5WOwcqtHswwjIMG1gaOIJK/g9hbwXXTAclL+hA7nx2y
msxjS7MKuZgpryod4O/poBPkYIn233GSbZhl0Qe3A+JG44dQNDk9wyMkYcU8cCWU
VTa/0Tv3Y9mPkuPWmqxO4GMvcG/dca37h8OuN3dTG17R/7vfwbCcL4HBtdlTdstD
7+0O/s3+FnVyM1y/fBdJhhRP7T/hieV/tVY34EyosUjzacmgvHS7lci4j/zEGBPC
aN+bp4nfxdVzChIZ/nQrL7YsWvSXYwVlOXP9XLKuCEfwCuXVUWnPTqLOnX24Vnl1
mN3vn6eYcMOoAE6bMG8u8i/1PHTWPNYUgrOqg7HAUdpyzhYEKamxnAE0F6l7+oSW
m7pRlEorBDkPe2JkyeD5bECk2j02uSsUmTWfQ67V47Ug0dbBB4IpsDxvCtt+Jj9z
oREkcqH+8W7MfZp+KnGGYHT/6LmtnTDADiDooOpV0qIkotA8nOjfP7ttiWN1srQf
nm1r4FqyNFvWQZ4Z9950OIsirMV35FnIxjGKJk7lD+n/h2j3Kv8sy5Yfh7XSqc63
A5R0kK2C8vXq8olmYe5smfy9s5KAvVOFLLtY5efJNdhMzg9jcPjM4c/8OuKyqhoa
0YhTX2OgKfW3Fuc650s8ggCkZQ0hS/IXvlr+fipcg9JcjR6z0XKXd+tvi8a4W9Q2
ktvI/7JJn6bYmQ67I94VJLoPVEfjRx4K+O8Rozr310Gbm7CgjBWhKUAWFrvTCMdQ
xVH/uGEdluxnNeUAIg9IzrvR7GZD26IdBenyTAwpXIkkPmOcmnFB4uVIpe877RG6
YWkWVvRM3gse2fwXuTECqOxhojWCTzfeB9Rre7UPsL2/DSdJ0rZI+KxMnDvPKCLL
g593Pr2Od4eDsljvvZZlmwI7sytiYDooTJynscLtrLY5CyaqNCwAJXOSlwfFN3EI
FMZldjdod5rP9osQBXaZLKoqXBwZNaLV1xITvNhpmq5j8fq8OzsQSx6FIEYLfnGY
Gj/SQJIlxhZKrChnCSV2/M/DDTHtpkW9IkL6aXlE4aOmXDvYZwM1tR3ZYtet2Ew0
tXSt3DeCJqcf8MRnWbyieSMUi9qYl92XSS/j1FdMwIPpOBoUIrvJjMHbEu/QLn4n
dNTQxMmVzacOZ/hPD22c+yEwxKXHsOZWkrhNVQ1Tk2N+QQ0kaEvQ5/XDBK7krpMZ
7VpLNonUQN49Jjxl8BqzPnCfJvRnFVF2RZdGvlqNEzCBk9xaJdQdoyu22hN2RY0U
4L+YWOBkG7eIowVdz99+vnxtteGtPqa1N9+YQvuOaRQzmGEMhE23zRFZMXLtklC1
1GUrSS3AnE1do3eKVTIWDRzkn9K8KvQs7WIpByi+z0zIsE6ig1jOTrhpc1Dx9bh3
GPb211CawESAErDO6cKGSvCI2+2etDoQcjYF2yhO9IUKzH0Q9frMQsFI/rlZb2bG
sr94btg+YcqVRh2hO/5zFY4i8Bw6qXcTDVQGPNjqGe1XJXIsvTuZQzFdldJOuQgP
SRoxPmVzjKESmUXWWgIP//m8SJ5Xb0M2NqQrSiDG5jTHjEcstn5nG13ePT4OtMd4
e+SRavekeQU4A0cU127GBnUcvH3YTm8vx24Ovjb+PUAGhUpBxAbU6PLrccZRnTT5
9zub/LJjnPpopQcnaAMiBaZtfld+JWVX5qWDJZbKigPHhRu2txDW253FFpMFvjbx
ofbz07SLIhc9BOVYbU418hIag73wqQuAAl5zjjJwM4NEeMSUlt2IDVcghdmIkuU4
GCJu1ByprImkAj4QDHwp0mfwBcdF/pXCAaJLrj0DPzNAnNqWYIzEAbpRZYBORshM
vrsPPjzxv0hL720c9QKNJ+hWFIQydUJOz305WcdUf+IjwDusS5BHTRtHg71G6cNF
K7NB0LP67cMxAlMS3xBDRxQDkXdMJPBwTbEe5aVuFvF0UFKnBm1tyAJh6Ldo4wGH
yIxK0oodSAb4KF99+PGZsIZk49nUvl8JvdYHt+wtO5woNGbZvCuouCYk3XRv1YBj
fl/bgx96tY9X4Am+SwnjOEKC/hi+jz0QmFbQblhe+X6+rNHiWL78Z8vzhfZZLMuk
maeUjcZzGxumf0nzUKEMoKWPVbqRh5aqsQgtZiVv/uKa+spYBWoV2k9vcoEU9lh8
fDfxz5YbdKm1Qj3Hrm0rl3VkDbRD8YE03kfutvDnYIPso0Ug/m0STtIeyY94iopl
pb7jCtxL2CupFUV6Ziq8gESpb47i9uf2Lls22OWZwxrj4RkDut9WSMosCHSeesbR
AFxWUQjRWjdkgxqEXwlx5YzUcmEXNexKVz7D8UVS8WH+Ga1hZ3aFxd8/sMjhKfhl
23lraM3Rf2Jw/MYH4lEfU8A6wD9s2420L7kHSl6BVzI4iiLwT8P/67X6sj+Et+f7
8uEyv2xISubuFYKOmQFXoSO+/R1lTfVQg1N4yc9ME4acsAxQMvOC8N9Cs+mr5M8g
N6hccsupo6nDFuw7NDrT23eZzrIsLsgRXMkC2N8tjAPOXbHZxYImwLqg6+pKOYdT
MEIRykJXDh32e3XWwQhN325JE3oYnBS9WzXBJ4ruIp+n7RUIrVnMg8qIjz+rqaSr
FfpNjXi9E1aedtjdsWE7aDcMBNY1Pv5S6OzHzYLowBlma7kNdIFyQ7xIhbLMYSHp
gcwpKapU5ljeLQ/z7vH6/WSFoH2iZUhRdcNpcOpMNjnGMJVmOZS/kpcQU5YtYeja
MI2AUqdPfotQE5jgCn1yTqyq7spZ9Uhe0KKHBoEnGksy8Jp1JxCGzwgAzV9aYdky
BpdufUnL7CtdMka7IueYLgyAsUoHPPE/Dphff37e6fA/scUOlQhJ1DryZIo2qyWP
4WwVo2NitSYPbjnC1n8xQB4IMLtx8h34nOePSabIVD38pTiNNF2Iz36Cx350vjWa
CH4zbvDxN3RX3VuJEbj27xxY8EeE/k9VRB2YKRCBJkfH4Z8aJQmH6UXAROyjJQY3
ucEeXtmR5yklnktuSVjzh4RAt4q2pC/yI9dwhL6Em/N4gitmuzH8RnTPgyCumDCS
+H7UWx3hG9nwfZTgZazlqyGZrOReN8lowL57tRtRrfcqEUFjBe/XWaC+eiUs6Biq
1r2GMAzj5lk1xmguKvq4zGr73qDHYxhEXQ9W46BE81u85WnHg+h0H0FoDjlhlyS+
wxcP3jLz69Ljksd4N4viWFIb/i3L1UOA7yX3vrPzGUVOIPaRH9laZIhFBqVVHkjs
EOxVyxsKAmuxNWWIUoRzO8HokOzVGEWygPg9f+6/P35Xxh4DSzkuiCMdtEM6WCkw
mpvFenRIaD/au4O+dl4sYi4ntmafhsQ9+bie5c4hM6YvcN7wl0KsqsVVJO4/JYXh
95Ie7T1CmTNYU29x3fBMfRXsuzQdOVIfEnVsUsECsp4nTZ14XKVOJDrViDGFcCQz
vnt2QIb0j75o9nBi4g/OY8QjAUvn1cQC8Mwort5VTeXGT9M7J9nc7PAhVy9GByDC
qXeocBlJSBxfdI2RbhOp2T1QOQvj1cwy8ijDH+Kl4bqtHB8A6hSjJDSs3h9dEmnj
K2b0Q9NwQvnbNd2z3rVgJRh5zbyLeFiVXsJ26I0MG6pCVZNRkGlWy+V338rEghsK
quuPM0O9lh20CTWrF2tpzze6+1gJ9SLmjL62nSDXWIz76isjYm93Czc0Q6yCqYJx
uhM/M8pBwJ5Neh7sWDgG/5kPwEIqcAVAGMtXltEggZK28rX+4ZEzPYtZezgOMiH/
A20t101a93WnOsTIFXuP83+glaTZ+wrGkuV9+S6nWdn+qQCNaL7V+bpg0oIUUIMb
uaN/hzUAYbtaEmAV8SoH9McDJMIowdgKcj24AtxUQJAIli7R6Mj8aUaR+CGd7/61
kIVb+Erz5Zh0pH7Rq8zhOPaqlWaZKflTg4g+u3GUmcyKQQYdXRCOIAWBOQvyy6il
H6ASpCjCnBp0VS02UMN8v0WLZCn5XRzYms3oEPKofcxv7I7q3iaZUDFM/EtwQLMg
qP+5qq9/u/RxfGoZIvmE5Br9HdkNgFJRa51nXw5ssqWkkjJt18MO/JzR/QIU5nxK
A/YojPMfsetRfv8oX8EVwqJeZaLebRIDi0WmXlCpEH0tv6rZ2JE40zzap56LWRk7
G2wu+edGfrKFdyTl5Yr74EgnA90IgJF9iFg84ofqX0Nu+7kfmjT+yCE++IhQEPGc
VF0xJF/SG6goDGanud+M5Jael7BMqk0JMNJHZnxWH6ukljAVP2QU1EErxULEdtMj
p4TuZzg49dP4BhSHL5Ot+Ktcp1bHpMnHGgy9G8/iCu6DE9Qelf/jpirqTEGD5RHP
IhCWC4lmc2wuoUgEWH+6fevCAVV7RyJc0xTEN6N1aL+Sd+TAnUerZpGqxApAmL7f
wEJziyKwWAb8oO6AaZAzGGckSAXRxjAieK09ijy8pwoVzYPy7ahA/GImwCyY3alu
6dK3uiioH5AoittIKjXYkNZDxXJNPG00eow3GP5L3JCfY+NuPjAfXIgSmqbad4A+
wq+Kfr3DDMG6Vg7BzzaO8bGdzfYAV7c5R2hvidR7JcEJO1yXyAA9rrQuE+H8rxHK
oFKaL4MDwuObvphSmMsphxdEVx5zj/kglgOslOZ7AyZaLf4aGW0m4lsXB5V2bKhi
rPXf9ZtTL+nURAwau7WBiTHCpAmLwozu/wz2z0jQ4CxIRfgtQCjcnSlmsXxmHEUX
rPI9BVggXd4geNIXOJLagLcN62bSXIQ2kf7BZTk7xJMcBDaaZZuaQQDHzaizXNQJ
gWGMXTTwTvdsRTZCff/fdTP4UsH1s5vvgevjVvxk0FZ6kbetL2Y8a22wxKbV5tQM
SFtcBuqzaONbUJ40izuiBkBgy5KjYUwkHnXb/dd06Gtvi/CC21DDBKUHHDf7XPj/
01rYiDupmMtwnqEFZVvh3oqZ/JzCNoSKFRtVOdgZHbORgdaqsOAPSct9THA5UPJI
Wvy/oUqDmNeeOSr1Yy9XjWkn+HakNSjQvoqavBbhsaAV0Oem+i2n69HYwJ7Ehe4I
8qVhxTUucwXHz4nvvrHz5elloD9WwDESxoGA2pOGJ5wCRXStOjryvOw/OT0aPoBZ
ZiDd4aqOS3hPbQPFOfDe7MkVvgpCuXQHpURzPjB5HKZjSo1l1WSr1rjwhNjiVyRd
dQI7sTb/cRsfgH2TtQ9Wkze+0t0X4ilEjZyQ6U8HHx5mbOu3iH5ItXhbbW0P+bAJ
zOvQZk+eP2OpvCDJRw1W3fxDJYK8/ORlgGZ09Z3Ysd9IZwAzkNt8J8LZAgWK/cjE
FpKzsGaECUztqxo191qdt9OiHkZef43ovy0So5MgRuozDcA4UlhqYL6qWZ1dKz85
XDWVOv6lCEaqhLBjXY0f8Y591nVK0FPafdErOkWSwX4Lpq/BgM68pEu3DuwcC/nz
4wgVZqkNcA8qXKnNUjFKRFGkgcWXz0mdRtBvh2WOUYNnxcwzcDnR5erJ+/7CgU/T
TMpE004EvSVQ5LsaeDSEtXJfke3KIgiSvoDb3v+B4ZRtX9b9AmuTM9yPlQoAuu2F
KSv2cckB2Jh6qo2QBmFG3xnIuwC1yiVt8D36sUUNi4FWOFRQlAV+YOUg0iDVYcQM
MvSJXwTXpCo3mj7wzHO9Pfhi0aCDewtLSiaomAMN+DsRKUuIhZKTb41mKKGbDF+T
G4NbvbSMRcf0DdnQUeCPvlmfz86pnibTDB05nT52J/bLAAH2Baq7OHxBZvzZzDea
TXG41lTxH0wU5oPOe3Aa/ZBOYIBTO/Jln9RwzVudMzhl1wloSD0jZF2HxmnmA8JE
Hyh2ahvVLyfj/1QsugRMc6NIT9uymdV3P34r2Ky+euJ6aAUEmJs2nGpIu84V4sZU
5mPpsZE1y6HjkM+Oqu6wZ+qnkT08YQhSpfyYke8l4Vcxg0jl0dasjRe56veXuHLk
SXJ4bYSHFraMjiXP5x725fw3ajdHu8P8K6y3dQiLEXJaQErkkcQ4T/BglcdL3BYN
f9trYYc4rciamSH4+/ghYL7AJQbOzWMN5N8rqo7YV/BV8sS0IsG+KO2l4nxFoxz/
ZbGtwQWRikvHJvH6lrNnBH1iY5sXR3zdf5u0gDyRuMxssK3UwUqU7Y5H9O4hniCk
hh9Io98UCpnwsCHdqU1QfyuKp6ZT1vQSCXRf1pXxgoTKGfGdi54FLdOtpC/VoSLx
cPlcAsBGmCCIFYhKMC4mT256kBmh8nUprnU4wsAzbziKaUTDgKJ6ul3u57x4kTMA
wkfOgYswMDBLsPSle7/AMO2YT0YAnR1rbP9TD1n6GYyehRLIw98hr3oLR2fLyPJj
XPC/sK74cq1zSkanzMT1jL5hdJBfYmq0zgYmn5whL28djDQSOO5gaf9UYpU3yzOP
Zk+1wygW85XDoqDIqGaZ8U+shcXJBWK4Whq+ydiKaXgFnqsIzN7MOzzr/Vrq/xza
2tkHSd//bAliUlED0kxJIZQNRhvlMsyd7NyXp1XIalwcL1iXiJYrNB+0GsJocO5W
odYTN2d2Cm6EOmBbN8gmRHasRyb7PZibhkZ+ZFMsIbwfChsxVyr9QioVcV5/b1r7
qeOPEysTl/UkVQDietm+67yZgc/p/jGJd5rxm09uhiEVSSeLlDX7VxdZsuIZ8AO6
xlUtzmdayjl4oOW9LZWV9BBVJsJevMG+QFIzkA9emsWgTM8ZQ/c188i4Q1WSqDmT
6OOPJjUUYrACL1/4qvplNo7DoUow9+uITL2WglYgj3se8aygY5FSBsoui/G97KM7
w6CzJrjtzSMvmPvH8vVNwXAWVpO5rwUuCK9VbASpVPl0ybQ4PSq6SBfc0RumUVqx
WgRZykrHSmv+uSh2WsSRza0nGm7A4kRGTOqVIdD3JOcmyZWcRaazyNU6mIbPd2kF
hRPKMGueqd8CaMBZ+wOV+rKIyi/S0qUfSLb177c0NllKOA5wNZXOhm/qaV3vp/iu
VQyqsXDYMhP+/UkwOpoBFyLZx6UlphO+0ujabHZM0MtaSMzXHXAQ6xOia2aMdbDj
WtcHsf5UUqEDyIAj5CegSlfK4re6zTbKZaz4Rmu5cZm6c7fWgBc61exrXX3bxdWU
D5zj1ZlIidSSd0+0OVyWSJNqht/1nnP3Vqj771ZT0+Ohva4gTEwEK7P/2sQQQAcj
WYD0BQY+6nsiVc6J2uMwY6bSHzMRmIFQRqqiZGgykpPwxlsSHU6qgQrf4rc3E70Y
+P3S7S0UTL8POugO/iT0AHlmitnvcK7rpsvQI9DXSrXW0YavbITgHPykMTDmi92q
yvRNRhB3HCrmuCRPgliIPRAV4Znms+IwuZ6JsbnWiq+VJ7LFzPBihNsuy83Ya75S
HEm4VdYZsWxugFfo+YXlpgTc6JNtjQBJzonEdGnsjqZ2YBmB3VkFEZVEA7PAEFNf
oxsuUlbm4zSJcJfrH89wDr9b3nNvhRk2qp2nXvL55xyk/YFJMd/EFAD6i4PB6G4E
xxJHmffQ6r9I3ZMDsNaa1dUK2cvKg9/pXvzqtQhpakk8jPbs+iCCqQjgGS/ELB9R
gphPzrW6BpK1s50nwB2n94EvTDellvFnXu/taBoigf/lASMRrAGrSgbaqFaXVugG
ChIn1pudY+zOokcoogCP/KQMl/u1pjNbQhs3MtYMOZKMMf9Bkft4s0clJv20CU6D
bNKKSSuFRBJIzKv0Eh4MXisDPIg/zq1plvtQs6KoMRLjqC5NpX5iGa1R55QyNBMg
0D5qStPignE6MbZEVWRAtMUe6s/HG0EHzUKdHwHLYHjjYEASznfyn3zg8mKTfNHE
jiGipyk2cYvIAVZ3iAEXlgfSBnoX1jBVv8exR9pyF35WZzCQtYIRcsZdSZOA8e1c
ZTPbppqkreclDA8Zxc8aQtRu53N85RKR9Kp/bBSfJiuTjFtqRiTmVZRStMdLzmmF
Ss1yXGGgpAD9YlySFMtfVCs++1gR/U08Z2YYur29pz6JH+ChxF+q2TUv4tTd0KaI
k9Q9eJ/+qfP11O9E4s9TuGM8ljwDxS5AQSklViDKxdgvytD6SCpvjExO+rg/oD//
CkB+BrLd0eWCm1ks69Q/jFB+st440Y8RkMZlhchOHSpesN2EleFMTRD/X2fXtgN4
7clfYME4Sjxwak6UuezrDnwasGndkJAQo5S48vk1G0cUsNjGOF2dxFkkB6NcZzIc
vho5x5u8s3VYAuWGFqsuG/cTBwmWLrqkpnzRFYC0cOt3VPujoM+WzxER7ZOI5PO5
WveUDpnThAmP5DX7r8MOsxNAEksBYK5g0qxv3h1gjpqd6ew5eZ9wNJtRGQ3iFiPu
/4wbsbRPHEX4ZN4dO2fNg6+BI9cjoJdKNZapmn5Y//+2SYnfGMneObjgMDpXJWFr
AtH9Vf78f6+/zHRuqW5jT13SPF+a1v3a/4pKrDaJmZNrSDDFukVTKZODMZnnJhVQ
yWNRCA12+loiAjLjYO2wO2aUM2PoJExtzhV/zoeH0qEqiGj580xtz2C2jZ2ywLeI
OOMZI4Httqu6oQ1eRw2pj9312qXrWaSsfg4Uxn+a+Gx0xO9qMTpgd8aIvqYfsXPn
NafcIQz2mmqxagWv+lNfp+B67rv0FvyJ5DBzGDq+X3y11Ow2cf0oN7n4CFYjSeU6
nRBQ98kRxuNIq97q3TEf9Y+mEGbZfGqJ/KLRhlpJTgZgMIeZbIqg6ko4ybOw2XlD
9D/2SffR/F1ECmbaRZrUwPy46utYt2iGKH5yvpRJ2HbK9Kk3mzG9OkMMtJumJDRY
HOcTVuG3KiHjpYhvFBe+vz+p4lRrckEmUrUY1/o6Wwe1hG8ThODced+ZrZ1MXWTb
0Xo5PEBROLlY9a4tDoAjOFPQSnvNLs+o5vnP8fhxX2/1ySAm3QtTMnHXHqesuSZ2
m1DKvvvZL9IW1kttcuYC1VThIHoqTDiLURWcHZV6rwIqvfNZYR7CR3/5HuEFVB3v
MPakyWu4mXTe31zBgOLQtKJmiS/aIh6qwDLvMDAmfnAaw5gLkLoViFEllVRb++3g
Ttje1y9qhOf6y/HbZ9Agk3U4KtikC8pLSKZbiCou8IT29Ahl1/gSUSCAh2C7lsQp
qqxw3QL1hRuG6XYOEdo7cSjqfpxviwWyiM5oFk+L2aCkEfpkMQPDO9WsQKsHDIDp
JM07ITc+PlK0t8leEIjFzcpzSIFJ2tenV7KuT24NxuKXpEVlNc2ir/KeSTiJkT5t
6qZ9bsnLyS90EfSxiP5QGRcFu833GK56CcqMZGgM+72AtHgFkQN9FuQrhR0ZEM1j
LpVPDnOfHtdl/TzbifG+gRM7eeJCl6HFm6dfFuTFri0fLfeEvzE+8Q6tDAUpUgch
QxZb1oDfSooIFuqNM7mg32nS4tMPgSGUviCA/y/D3yJ7BLN8fI4CIXlv8oq2cZN4
QZJpQVhyl/z7faTit9wbG1oCmeU+MhdD+DHRc+sM8G7mDQcMQ5XfaAN1CizFxLDW
ATIC/JBWotdQeE9pkg5MhZixTE4Rl3I6mgBtJgbQ0HPDBkDd4V2jNVk+wxkqnLbV
kDhuaDsnPkxV3BDNRWa75uAD2/JUSBRdsIkbASODei+GfhSEkSUI5cyrREpSVbXt
GQHRuQiD/xhirCCXqmhSOSPNJsHx8lNtsDReakG7Dw6vA2BYwH4R1CQOPWZmqjJ2
LJcgm3KLXfZt/R/nmcBk2AovIj0MbG2BoaZBmbUNamhdXEGXCYg+zY60s6ngLu8P
vYKsrpN6oFpL28YegNeg5uulzKjtPLLkR0gTJhj801BbxcNtYmPc/1i8hDM2lkkV
0qOF9AZ/lqJAiGN6LB7VOvhHvIwuu28X1NKlGqyq5pGG26+ljvGR9TYpCrBi9jDN
RKcj2LCxViHouM52dG7cAELbcXODhPO2B4Fg0jNbmYOSANZqasJ3TUt+5F2qg32h
PzfQlXqh6GX2XmB4v/GjdhS/zjaTejv/GF1FLxFh6YdPD+Mfw3/qowMDXW0f7f72
n86nTE+d/S8HRGg2Ms/bWKmVH+ZMv0tjnFxwHzIkxHlYobTxer0tPCr2V5kFydS/
rwRx7yo7NnbEzaZ9F6mGSISL/G1GsPdP4ik+rQgRVp/kNr5g6lKL1izlWu5wKXJU
mBGJhnHrutDgtDsTueByA1d95XJgal5bv8JnXyJV8B3uGhuLdzrqm93LwxpffXne
hHz/9JUmPCWss36vc1XBMxbbeDBXpICIXViSQN8Ql9xj/osisNJa/W4yE+DxlCVX
hFy2EDi/ap58dNNufUWbcg2DSuAExshgmHyAoqnAaoMomyjw2k5E9/g4Ja78Ownu
yBInmSNtOb7DJnO3FAE9/TYUHHU5YtB/LzfWJtvrmzrfm5jxdOdPSHj6K43orWIF
SPaXVOpgrPD7nNUJM1xntEmIbeI7CJAJl1BD/eLu3mlLQxmKQI21v50Onrg+6k47
Z6mRLNnut96vg7v7j20S+LyPMRpugPdF6MF+DlvwkWx7bom/3+mGep0p3+XPmFsa
I3c/AKOMBbUBxx6FyZUAo+rvK2Tsmetmoh1NGnCfmpnMrg3NrzkdzAzrbk3+j/VG
5crda/kb0YnJNjElmPYGlJAToc2ehQvrSO7ijSpVhpmNKWxrFq96LOBNHT6mgy8v
CHGrcrciT3Cdru/uWXu+4nYt+U46XUaKHQfzuJQOIUmivHy7/OV9GVVoUUtR4crp
M0T69NW9GVXRcF2UhrdllysylAukO0HPl57J5DVo7ld9FqLmZVpm/9iOkVsehicA
Oa3UHZ3+zjeYsRKc3z56HbBggXsrzhAtdaOYWRa2OEr2RrsRijvwyHrmmkdbYVjX
XnXgu4amN3ymdSxrMGX+rZVu+UPWWGcE8MPhiLD7B+1bdl128K1WonuieuKk/SAh
MeCHwkURS/vOvrj4A67g+TDGQubSHlhansWy1jbkzt1pITgsfKnSFCTY5ahXT8mM
PGkeYAuCCKFWtCQIBrPlBjeQc66FY47yCUEz7b6Fa/KMuqJmowjK6mT+IhE1m/A7
MbQtXOirm36rnwDDQZ3ErTixiPqa3D+p1naLAgd5IORU86lZZZferkTvEFMreKtR
Fsl7fChx6i/XvqqkDXKQs8cbc6ZGsqasT8RM959CqQoqqxoxwjjyZfEClZoc8DWI
qhcUVzZ/k0nda+1M2MSzyxnFgk1YrDDL5YMbIt0xCgzV3GsggfMs2g1/FJldSw8u
uzxu2zgpiQFqD7qC621E6UhaUzgv7mVPem9Cmfbn3paD8wKOBZVgOd0D1ZElXBY6
n9fgCdedf3YEmOAV+XfyQzRzB9+TuiCle1H3eTElP0GvStXYMhyxfYXdfg7sgj0T
2G13cLAd4S2mZ2reLS8hWLfaYuKacBNlb8Z3keNFa9mttB6CwyqLU4+qIEp5WcUp
6kG8fz4jkU1RpWpw1QdercOE/bv4QfVm3bFuiGpxkS+tyZcp/7yLqm+fAT8mVKax
QzirjYBEYJx2CqkLC3V+GWmxKpwiK/yjwvNMEL7mZ5brSgUq1y63msb08gZHQapX
wUEKkRd3Oagl2R5HJ/n86SDF/rIRDs2fH/YxIF7rj91Xn6vSPyx/wrvihaF1IcJQ
F8cDIN1s2ZprJeeQoZQM3Tpu3Js6fn1bcX9cwNs78tsRnlJqso/En/ZelekP+Iyw
xVTK17DQPANqUm42g+GO5oYLFOy3LaAmhjf0qr2VPqV7YUQZOFbrFuyfdSljYKZq
G0CdOF+nuadqkMueo+ofnVFjKU4TdUr8CvBgGZtGzFouLGPnYqt5I7drnmtlMXE6
i2upemWVveAR6tWHYPpEJOqnSBa1TaMV+w24Qhc+DcQe9r87SK0ve2bLuuwT2TfV
HKTZHvRAuq8jFw9+N53+N6PClWDYDN8yJXJep6NE2KTtj5DxvbeuuirEBy6mv81O
B/tjz59ijWIxFshOt2YvgQDWpeUMLrVK82dKtgrGlvSrDJtvTeUt9JCo2AHH4xEu
qNRu/Y/thJIgd7HPIjd4x6Wpc8o8VhueMwx8t1lSJzGTDKrcMxQeis4wmqcwmvRX
cjqZd5VNHNutHh6U5wRigqZ1HCnMwnqkE0QpzEt3iOPvehdpg5rxFbRarbtpGE7v
wMo2/1yh8ByXYwK5NoSZ0kEb5HMaAC3nHjK1FUH2nIqGKuK3ShGBvESP/QchIFin
1TUFAIU2UGNTT/z89jTbv155frews07LHT8rP+nX9liEGijxW7X0RIB3mMb90lPQ
LNOGzbMm+CfVqXbgoKH5ZyKvVMBmY6ef6Z+qe6BsBmz69kkbXtZ9tkil3056zwTL
Nm4YlvulHhAGWCt7FLWobhQkyUT7sl5ox2OLE9wuZZSPnZ72vEIwIxx1195Rf0CT
Hs1v9UiI1GKENivkjvo2Bg8zF/6lPMg7bSiH0c+Y2GIjAh7RHrmi1x47X4wazIFu
1K/G21j1iQxqndIqoo7fvEVZ2OS7iKoa+XjwLbbXUo7usu3UDrjazn3DIk4pNDRV
u4ilekwxrD5mQW9x2WFs+CRwynlbcTw1iC16N+huwcV0zb5KCPXP1trDDsQ8HHrF
ofggOapCqLzncEDdIr60eQLUd73/qFoRpFEDQSoweJTWDWyIWchKlwtLg4qTI60v
v5DobE0nDCJj7Xg3W9uGnLd6STcD/KHx3nZva2M6hZ9Nw4aRo/sIByq1iq02j4wj
DkVeEA6E6WVuREh9+5p5PYOxx0ct590awnRr80MTyZcP0r03anZppt6waztJcnTb
hd9s+OBcTS6NpnINSp94VZ1PBkhBo+ZYiAaN0t9FKyfgBS2xNgzN7yO3p4UgTNb6
qe3AZ+n2flwTaX2l1abnLjjew9trVfci4+wQr8j3HRMUgLVQWt4pbu+eu/YqCrOA
gup++lj90S6c4deFgokkHcB7awuE4L00OweNY3NTcuY2EFfgzh/3eAIjoKqGd15r
PoVvO8v+TmO3roTTrRSElW78NKl5llAIE6rVAk6A4Dud3SWIuThGNNar9+yjNqfC
cm+bumjq4tCC4XxKco0omjE7uoCXx3deR2S5+yLq4T4smhIST5sIa+gQW24jZ9OB
CiwPt7lPjtWtlRhoYCL9LAVIg/G3axUo9ca2pjXIDL7prAi+OhJVdPwHgkaX/JQ3
iSHqezm8ukNpu5CqQBktSmKjfcUtoJowthjneolWZ8++iDlNQIa/XVjajrmqrAr6
dFJDNqHZAmnsbR95Uvn4ulmWW6TeZxQ6xDgHDj6zewNRBKujo8PMRQAHSInpHyc8
tWohqTSI4FKAif8QR8ZHITgCtZNCgP0h+zmXK76Gdx6JowTXAZ1fb+kUYgGn6R48
ucto7kq7Jdx4gVUapYQlxgZIVfMSAx3/c9MIUkWUiFpPfwyMTKPUYntwP41OVQP8
sLFpEkimlRHn5o8mzGYOpfuSjK2hI8sqez6SNr/JQsM7h17IICBrdVR/HHjkyrFm
BYbuVskflZnCOns/hyOvY56UuMIPn94B9O9HGxpFxulSyljMw3KwwwScNzC7smoV
bblW9b+A2HoHQY8jwkTRfPtS+2xKri11uusSkRWSqq8TgjDfRYDtYhrJoTaQtfZF
KACTu/X4KdIM2OreChGrMvVBYjOP5uO6zpCqdvp/sQqVwdK/dcmPtRfRtF1K1h3b
E39rYrWVZUrqm1SwgqKzWQEteiJKPO/Mx36otuLyPJmBDaKBkGcK2Xu6g4y6i89a
ladEWgne0iQg/z8LjXNOQB/JfWzfatNkcPnaSiwd7jIvSFEHow/PVyDx9JjRbKsc
y5OUvUxZ2XCEKck0UiklzU46tuBniX6wbDZ104APv9/a2QOLRrE0m+3n+RaEmynQ
JV/Wt1nYyMwptvOJ4Wd4nBi4s1IoTNAEpytW/dASWctps9sDG3xzlW9Tbru8WXnT
n0n4itNBwUGXPzDgPzItqitFG7BkdQy+BcPxn620kDi7KXXAcfSMbb6ZhYWuXZ/Q
relwRlUF12xEOihzJTpEyKtX0kHHmMwHMQmlPhkJx3zkC6QbwGApE1VZByaCuKbU
WlyybRcduXDFBzWLNJGkMWtvQK+/BXTkJZB9uOs1k35aNoeX/G2Gx1vMtXtVFDJt
pxx8YyPOlqkDwLrnLjEip3pCvqQvnld8vfsVnbHvJHeN17Um905Nj86XbEq+WG6U
O6825zDqVTDGKxHzVwsDp+Tyy9B+UHVJsDJNJeYQojY1bF7Qzo7UtX9dt3bbZTCh
wW0XzUNO0priRxSanlsm7jfiTnO5sZ/RCeS9mzgYPIDH17+yKVmNVQkYU1Fhxr05
feWto3x2D2aWMwpGzdOjrxCWirHiGG4Gxxzdc5AaTLyuXwSCuJ40Tqq5+37TLx3K
0r4HewIL2n8uxbA7H1o3InGcecLnx6v1ZZgODnLDaZc4YOQ1NZcvhkLy1dsyL/8f
UOPa6TaDgfCrbR49GMaXmvwXniAzINNMrlTiv2EWdreWztLGcn4yrY+BWO69yTwZ
e8qXVshrGQhwTl2Pk3TezpX4iTYYsqD+1JmEkLX2h6ZPK8aU9bg4kpqO2O7YkCZc
iOLiEPMWQYfsnin3qfjxwSbhaLtub5LnjeSPfr/IBuQr08VuLgi67+9s/HN0P8m4
vlDBhY7g2u7qT9fmlN+TydXpldRNBp1DmGVCF7j1P8w6KLYrQ6ghNoHDKdNsLg00
W44zwSvG3AnKx++bbf5z5+j50ZjpUmXsyDrB6sppS7LVAsnbGaVpgnED9PXRQ/8B
vVkudnPJVpdR4V6lsZyszFEs+K0+4+mcZtfkSGWAKUUEgwAvF/n06PwudYJpqliA
/6F+q8rUYJnA/O7JWwPL/s1vm2y4AIye8biYKI9NREWKTUMhpSeKPqRfCsU5GQlp
m561hBT/wU8Tp2j1nP0GGCjgnhhf+y1R0DmnhitmwshbTsxdrCt4gd+yLIerl4Kx
6MKobh3x+awJr9JBv/v2C4KtSA/sM3MlfdV93+ubNBXucO2X/6orct6WI1SALzwP
9MYW7vovpI8eIm2Qw4jj53I81tpFx4IonLCHZHSrmSjLHh/FlkeYiabMevb4B9Pk
B65FXiwN0EKNKpx2FAoEPEnGF37O5MSe+e1L24wSukvt/Xaly9+7gj9xUoWmZyJV
8KgBNtTqvJcVlfHKB26zRLx8YZyal+BKVHgHhknwHouce0+dTNsFQn7djk4DZW/r
Okfdo6akC8XjgGxUFtEizrjAd/8nXn6BsjJtr5oS+OKZILsn9vmBEOHxpCvqAfg2
zYIHfXB07MNG02ZydRuIzr8gNFw7VUqaeOs2sQRZhCtDHETlkpQZLbwaA8wrygJf
xSvTnrxpLBFGvQh4hY85IZcdBUmW/zG4YJl5o/2vcBKOI7zv7EiJU2cOK+XEXEqX
228stLqRoyglUUDAQI6xqGIIp4DcVY8JMZh3amB6fZO/lMmvMYEUxnM++tpFd7OY
RkYgUIc1PSBIha0OthOu3VmC86vEIgxeRJKmlLQeE+ScF8zoBPtyedMe1TDPg7Cf
0xH3Blh0bQYuc+TbGzmpqP8Rcs2N2SRtISvsNImnoWRzAAQQPvqEf7YXGbx3KEoO
m4DVsCjqMQGN8xKq9p+midTAtLsgYg1Zn1TbWIVb8iEA9q13ix0ULwUcLrghNDvD
lQUdY/B9xbcIVhrPNksDKoJRSaJTOWYw64IVEx1aEZLS3jOYAchcH0rKxJkJ471G
0Xfx4fJgAYSi4CB9B92Atkin4i4PklwmxGIp+6aX8S7l5Rizfj0RpsDqMslqZj6p
+OH31vOmPqTw+xaGimrGB3JO9/DSGig2VPxkCHaVkmwzZ7xKebKuSxmaFUv4VLYh
RaIk3VJuRsPC+1z8g6D5OOOgIjIVsntxOd5epdX26cO4TyTQvfLE+GrZWMacBqyi
viAfv2j9uHF3TgMoZ5iwEdiYFDYHfRuZR3aERki9Mij4vIte0/7PgY1W3FQHkOq/
p/zIRx4D0AHQlCpHeHNfVcJowj8iiKMh2goJSOTjo4AbPTYv7xnoTOg6S3GfEDEp
9pIo53uZbeqDIeAPGq7XhCp+OXazgNHYcZx6gvo5KFGbaQtxowkHmk/87hToin+I
nSJOBqdjaL2zGeRuGr9QZInAtNcTskPEVLi/cEg28VXhTDQst5IbimlEqY9kocYP
udU3Moo14iBd7VfJwmjo0gTSSs/WlGUSmglczx0PdtTDog5l6+pThpdZIy1LQrre
CRamzZ3GoNmyVHpOvSZK46NwfOciveu3RmP8nYm1XA082U2QZHSd+407Mau8R4Uj
fYgpGfyt7xP47BFojZFCwk02qMAjqJb6CNKS/mI3mdDUC1RdTbT4EyE6lPkjMHsG
ATgPYGhc7paqnjGWFu/xQFpGaCL5i0Qpd7mCFJy1vonzEiBwcS0pyXkZIePhN15u
R3aK1hcXp1RahBSCoXZEjW2cdySaeokIFr8Jhs2pxFmflU333OH6Tk7LufZm3gkc
Um9Ro0YY4t4/s+xJrIZPlO8um25OdxouCqbtrHo6rDOnZpuD++2MepGojCFGTbDa
rvPVWqpTjc1HsX2tqt9uvA6z8TdNIwQiHkBeIthcq5ecwgBLTZfeL2Ku7Oq1FKz2
vJ5/jNeRCEwjePNBMqu2/wPC6yeY6pmc9QbCimfLu4Y7+K+WtGN3DZxLMH4n76C3
XPjyvtl3NIJC/qF/fbJu6O1wkVmZRZgeQVEqduYTahiTENxr8HxJsG14l7fYJd5q
GIFgN57ZtaRLzW3qYPiJfZbsQayyik/bUNZH3v0Iw9xnY6HjMT7C+07YQAfd4ZxM
bQOM03GgePiKL8+TbOIfx/oZHj0jC9IO23R2QW1DZrMYCg76nHJkdeGPJyYo7QhM
g4CS0977BUEYr7cgrMeCRll5Dc9a0dkTjbaXGMskKs3v44rnQ3x4S5mEZ1Rs5iG+
xVICjyqi3fLz221R5UCy66xLq9zKqWrUAFCeMN0Q5b3NCHvPOf8rUt3k1DQDXbxk
hmHKkBv+JnQu75APqt1fOM37q82J+NQnRhcpQqIqEnv+lpRMV1ChKfvhi3Xrx75p
mnJkDI1NhQtn3+j37QllpdfLFflUOxzbuJHJpGQcrvsQ6OUWskGeN43RTPSTshOQ
gRgakK/YOmdxJmZlxa7BrDbTlx9vyc8RSQ9XVtgXYJVfbWrhzFn7qSXQbfdorZap
0l6+kMIeNOXxn2GfNxHCmr6S5M7J2kS/8c2CgaXs2ZCfAB+ydJcX6AFQ6q/Dmz7f
2VdpdVaXM6gL7kTe+m0T12GJxs85D75bUKHeaiY6Y6RvrQe5agWRhIF7yw1KyDyz
QRZQiVHkUnFvsDKKSYDhMF9t1W68hFwY0LZLUsTOZNAi/Z3p2khZCIsKqOn5IpWY
hj4JkyXxP8UA9bswtFbjub4cPWjow4bVWOx1kNAgAtagx5YtRHTToi1eMeUtuqP0
JuG/QbopMXn14fqCk22w1rX8xyNvXbAgwJ128U4RWP+QZtE7Nd7OSiWipyw3alNO
tv4ndbMPJjcQuWoZbbP/kCbLgFJ0VLJAwVcUsQ1K49QCzk9993JcWOv7T771pjSC
UQrS1ZeD4OkBABBP7/ZLVxPxgFg/57AKCsyyfCwYF0HMloVVcMFokaRR6Fowxnf2
yC65W7zci27XuDHTmuy/nqqx6MpQvROJoWwoWm/tF6ukQjSOOd51BRTuqNR3v9El
ccKK2YbEBeeDzBjNfxClOwh4bf7spF1/u2os4tTxFxHCJqqInMM6WxUKhsn5q6pt
+fcWyaqdfoVEtlXeg5ahdO6YroX2Y/uWKbNPnY0Xe+vD21nmU75hOtYzxjj1rchZ
39Tz5KCGJIdethhAiqYlKvJTrdw5ol/FNB/7jzSDxXS/5VYWma6B8khZdB8BeMZc
k+yIo5yWeyIw59NrYJl7TPawGSsAHDY7w0jFJZELJYpFWZ+EDbNf1N2B1NMgLgCR
XqnFXnEm0Tx3O787lWc3x8w7fk2PxXXqdwz3MQUUojyvIOa6uc/jAhDpi3/yRU4a
BTtjRUT0C7rErSTX2mpgIC9b/2f9rtNZb/qnwhGAPYquyxe04KxukfKICyPCKtm8
6Mz+/YzGN+rlVQtfoXR9n+AJ9zrs3hZhTMV6pzFXGAOzJHwIZfkFu2cRoyOBhs6u
i4MnH0qEeUEy56wY4IesauEyaRFxIHOY/pPXGOttoBY+xJxWiACNYFPy01CCNV+T
GBbtwxF0H4fhtFJ9CXbX9fCL7iEBUCJwJ+kZDxqFbt2WuRGSOpRdUeuUf8Lb1zj3
PuQk76QOn/RGG49koj7A04HS9/6CqLDyrEsb814T+l3wVHtR7jMcHdeXhdnteygH
VLAqD92FCVj8468CFe+HKhIRApFfz2NougMvos/WAWg9127b405z5LO2/tWP/7EN
ycAEN6Ag7Q22SapHx8BOcK6sdJInw7iRPh3lpd6QHzqM1dgIZ23D4FOCdphZxMeB
nEJu0t/A8ULVMPMBJ8s+855TWncItGahedmtIxu5xVK+N83/N8szICGiZMm10EfQ
Xgfon2w2nf+6cMHG9E2VnySdJwVZtM4Z+DYN+0gUSmfuRoJPKz8I3nMduYdjtaL/
BdbvMALiUXN9FAlisaQzStFduqJB72QZZHF/xmBPLllQp4qfmK3FdxUGv9me5A74
OnN6OsnTqkPrDjgJdXYvgbPO2FjiKgeaRf4EJHXvHwPDV6C2sq7Yr/QwEoOz7Pi3
nJ1qp58OVz1cNUZyvivvbOmbKy/BZrLQ9ocy6nPib5nyWLlWzHpgt6sB/5zc/HX2
U9FGZYH2p0tkK5l+fo5ynahgLbE98lWBh+87Xy9dKevMnTaJ+5jDddBN0k5TGqu8
YOFVqqadb+VTpjeUCiEAWH6aFNlGDmquzzTqA4aH7PTxOE/cxr6jF2HrnhRSD7qK
QieoZQJWsJvhK5nhv59wSKEJNCmrtZDutQ7T149MlMhGGSFdAXFx9wHi7k01496H
7vY7CS2Ny7xe2+e+LB41blQ3J3mpZYObyKc5h+ffLDjV+yUkxqqtBywhttnG4P8b
bCIiK/xPzWOxnQEHjZ4CMFCTwnBvxIJDDarBBk49Ej1arG0V4Akm763N8cLQ3ILR
0maM3YJFkYyfn3UtCuJBWcdvJnHavffy3Nj0pPcPjecyT+YMAy50HB0CIeKQk5B/
YGOmUvk6IIuhImkzqbK8SOXAvxZ2+DmScF75hJME1E+4qEKkjAACE88HIf7RqxGv
txtLU9uGdOPwPtG6itjw6BuHwuj12j+5+p9EDFpI/EfS3xHn2ikIjHLQAevvyDP+
Vj0vpQ+RahnLCSIcozyBl1wH6TUdhBbwJMkKoDEBduGiHCNADCUBkg6hIh/JCLXV
LBmAQcfiSJS+lnClD9+RN703W/lMy9sb0D5qAhVAfLR+ws2PXLj3PSA7wTtrTmJR
92ZCIlfG2Qdl5MltDVXDVDh8gzjOf05HmyC4S0iZJVUGBjHGMq6a8HS9geJ/THYc
jLtjFA0rSYppeG2qaoaViD4BWImg7TkmEHI44YAf2GZeTXxYtM5KU2qXxtPXm9y2
cOGkJNMFEOG/HvSrBhvs2b38IxecBQm9kuiv2Aig3xbID0O2V3KkRwfvqhuZsMuM
7YAEz1tWvHRJ/LMLmPIsBDVyBQJfl0V+2J5cq1dzkUXnSQkBl3nwQWOr2jJaJKVY
y5gMTCWZCTH2R9wi28lBc7tOHTnqBt16Qj+xqvBPqvfHP1QUZfsIBZqsQ6LL7IOH
9iqA1mtBxcFIkQXumCSXIHjclZPaNtML3K/vXo/GEZzYFiyfIKw78+SaZTZxtwwF
nI0B2j3xqZj42AdGVkhQtNzaxVvNuYWyhCPNFhNKRz5qabGXzY2ye0kGS9w28ndj
WBVE8y60RHDkJL81hf5qAtckXoFdek47uhFlBsI8qA9C+JeTpt2YnTMWGVGBvCJv
OpsQ+XgOKVPh/th0BZMyRke9CrifsNqpqc38jOwlyWA2+8ON3qpg5JZYqEinr8c4
SqGXB3cPFX8w0SxNSULBUfhFjOXZg/Dc6WG9xuWZmRSAgBvBZlN5gs8cVhZT2aIm
1CG/0QNv2LZsT4Dd8xLFWCVDwgA7Fl85kHko71NlRRJcvMcGtzLae1BvZ/HQFYqr
i5Ovb6AuuDl+5B3ZgauMn+GPx6+10QwtCxjmL9bKBHYJwVIr5HDWlJlp3RP273Ff
BbLD/qnr+Jn6zplLXHktDZ7oKo04Kx2KeHAxt4AQ831/NvMc0xi4Z/hkDqOtaVEL
bEFs6/CBQp1COHKuKu4wn2Q4kBoVqEpzMp+5oN2xHKL5rTdQIsQKyrI5fyj0BScj
VF0UeMwJec0lCHoODM3BZUek+9BavorPUeTrm8rWABp10WaVoHN/q2mUTaI6Ysnq
zywi4vl9Fmh6y3EMezgqNlNPavBYDLDm3wfo22RnCLbf3w10XlXPJaA0EbWYHeSK
1auI6vPfzgfMqEmjFns8zj1Ou7/qqb1z2Eco/KACw2hzZSJFm0SfHFVVu2hv2N0N
gsjrelyY1wwm1nI7jPRrgBbdqNLiriELoWBOp9DtUgjwIFpi44WgEH5+J2/FNjTJ
Dj4wbEILFHihCfvnodqPoAmLZkeKoAYzRWbOfeasZft77k9e8bVDMMwm8huuXu5i
LLxjTLiCaw3/SZd5Azmu6U/76pXNqzHl0N3D0PFGmKT8V0QmFeairuBreknb0J3i
+OBI/5SkGvvR5KeRGZ5xBUMdzifdZJRzDoGtEq2GqJ15Ed4Wb7LcYT0WcfpyNuBP
kg0U1aaS0dgehs24qDQ72S+2rh99qGVeCirxd2uJJ1QL57wQFu3Xom3NhoiLxAma
bOrNF9WdYlZHh9+vAv3PMA84fCgkoWqYRvq9XcMp1UGSczjs8ztNNCqOvw0aXR1Z
FgUmi4gWpVvZZ+mOyZnFAssW4b87TQrx79a99gXhezeFvzOPQptQrN0nOv9Rd469
I5j7j5ZRfAeoddeQh0j6fgVvQT7zYfIxmVpuCMeIcdXa84Ht8jUA7M1qJODfVsEm
ZC1gfszaNpEzHuCl5XX1yy8dxKBiMJ83DeO7n1sUkW7AGCVntXD5qZPZ6iY3u6ta
fymalbsdtuXQDnszUUaGE0NQ7TEeRhS77oIPh3h2GzmxwhlpwAQunRQ5be8WPFSc
bmN8Khqwmip2QvRHqYJ9JzM3CItqzKwnS7kyCTAL4u9pw++4XaIREIuHOPZQcCGW
edP4ZzgGx0qgaKA3SVz+9DtuPCDeFUioGe4t8kO0Crq2SMRn/L7uMxInuiCcy6cc
K5Ahsy6NgsE48q0tYSbcEmlbez4q87PKSu6P5sdVOdfJFyflljpxj2baPLOc0/kn
fW1hvlWZG6H4jHI1OmBdWlZd32gQBXznzxaw0gJFgIHzgUlUdSQuqt0f9UlCZFx+
CU0jlf3q5/NUKL1GD95K5XBQBM5f4mn6Rk863J5XzDc/q+eYcIkEqgoPHt1C6CXm
m7jH7ootezs04cFw8wz0tUjSbGwL1IpRUuJgIYLdwv5ms8+ldLUXdoGaJTlWPrHu
AXM/g00JRVvVlxh4MR+1nqmUmR+SGDdlbO5psnafquuQ95My/Ia/D/ejWTfkBdQI
D9SN4O1JVmjzjC76IiFovHvp7Ib+0SNKACnqD37QIMT05v6zCl3KzQJV7Guz7PwI
wI3OiIGHXPvJrDjFjKLoLXcCKCxDWnyiZ4NBljXLtrYiNfNtOA48ByKAX+85oBqo
h/RiXsrO2zby39V7o8TK7tc11kMuKO612HPW7pC2WamSdMxlqKe5T4NYPrREAiGE
KX6q6D4tlH3KHu2rMsZhAD3hLGcocJa75DdTpXz7kcdgQDOGPfO6AC+miLZS7WFW
73KjcSW4eyiX1jqourZ6Ak+7r93JZNVtW2+KF+bIu57K5TAc+rFFZdCAtN2miYJl
ysu3PZmWXB/rR9ReNBOWPe/8F81ocLAMoVYHbgEoKGgkU8//sbp6Pqu7+pqpPyNv
YuoiiKGqpxvsNISj3pYlDfR1WjI7ATN5V6npVEN9BTXFJ6CPssVniCkYhudV5PFM
dh4YwF/1PK8u5GFgG3Fxq9SK4moJ6dr7a6kpwCoeoZ+9VCIlOhUz2rNO7lW+etl9
nWYWlrcumg6v1GFdsOKgYC8Q8ECGT5amp8u7i9yP6kuNoIQxKN0Ai2z6oncYze7v
E2Of7IeO69FArvMkJv12cFpufeOegKsh/Stop7T9vSqndQZuQkHK8GTP5fnPs6Su
9JHTIjTymqTXe4Dx9iJPjXiqqV68jp74778djkL7IPPwiT7hWksAFn6dLNiucpG8
Ryz9BFOl+I9l3lDqxjFmb08fwq0v/W9lp4RpCPR+0PjwoxvFdXoi75mO8To8WEyE
FmTcncr1HBS/5wHmlK5YXmiIFxRPSoemBAuGUBpWJUn0XX5KoZ475zx5Umo1xQ5U
uckTKtHLbIrQn8okFTvmd+aO57Guxmc6EoRJ7DgapSmhRsBcMxnqY0Dkc9BGZ6MZ
IJpHnUdtovctB3d1/OP2JIqrcZuO7q4TnMhWKGcBMM/RKPht/kgqa/H8f2PePH29
E1W82NavF8oxMnRs0m7EELwDNKyBVUhDlnq+saVSqXLLbUz/TtVy2590yVfkLfX8
hLeNA3qeBCi/pWytyCwuNRKE+tqcx9vee2RIs2jQ5DJlk4Cw008J8NbyBDa/BM6k
T1/IJXuJ5xP8k5E9xFXEqj+RK4yhOYtfiNPQ67YGFvLRk8/AwzXE0oy6QS5gEyDK
utyKOEznqZGlsS0JJJIoWVuOQeejLmoSP5CTY3/Fjzf6keeywSzwYVa3e+Qsu/pV
TcTiwaap5POUl1i9ZoyfhRmAIrHQAgOJD5hYFBoMWq9UnNknEa+AHYptbOiku2my
m9M6cc/xBYgX/tb18ou9bh+JnwjPFtPt25/Ln0npqbCWMMzV+J+O65rhlUcpk6iG
XBVopyfr0SLHExop6rYBm6hOMHTy+qYQpMOA3bTBuGjnWElMGzitj/OGVvaAO9yL
x1Kty+mZFLaUfyuw+3yIMPfGeq8+/SU8G/ZG+Ua3PM+kxTUfUTAUxI6b0ft/eM2U
kQ/OAT6X/AwOTh5O/1H/73wEWkqYk3z1aKBKmFESSzWJSKFCd5P9l0WSJHRUWzEd
luUltXO61I6hmPNAldeS8E0cLKNvIsbjOrR7xD8NQEirtCWSmdHectKtqTXLlgIv
lzidjn7HBDb0SZAl03C7iDKatx+IWXsR3JbIKOP1EojLik/4/3INOaitYS5fSxCr
884LIpstPWs6ARn0w2ByjuAEdQ7MP3LJAegHW9safAKevOrXz7AEfDPGFP51lCUi
Ys2YhtuoA4gVUXwsbaLFCRXiogn+Z0fDoj1/X/kYMNunEnzH0jKnH7lhkGW/xPKT
ZSAUk8fXoMUi7kOtLRnL+nAxWWBIRhqB/USVZWKJaNVvs5deiD1uRdEWGaRwBIsj
IbtznIC/JalW904Qw38cFO2d+N/tfDkYF8RAu8xm3xe2x90hshJLPUdIW9nCKnyj
QYwUceNLCMnPq6SQiPoGujjrYTRw+pnDgAjJgXn2IXWjQoxo+xWzOPFaqp2Dr+K6
ISW3s/l2bmpHoEhgEveA8PuWjekK/SnK8mErxbU9SEb8DCURduCpLcs2/lA8WNG7
mNBl99uf4N206RCl0orVcGSG3MBWntD2EF5jmiqMF16SZl1IQ7zh5tEkWRlp2W+s
PgylrUCrkFE4YYiOa8LT4sjVI1r7VJjcZbGkOnhIMEZ+jkj8luGg8x2TiJtf0RI2
nqP5+3+4W71T8uVEEGyWo5iU9GWjmLreAnmc+DM0BcLwS3/DxOnnue9iE7wPKjRR
AzPv1PEjkCjpDgfB72tgDY8b0TPvCX+nEUFFO1+Wypyh9AAk48TneX7C6OlZwtfm
K3f2mIDt702aOV4ah7cmSEsMNrcw2GmEIVQOFZQkFPK29llV3xp2Hfj825Qnlfzv
EOb0z0k4whnWOt1doj8B5nGO6dBR7vfnVgHGK7V38VOWWP++nAtEGOLzyFc1epyr
mjDq/bY1Qn3d9Y9IlE1blyZmbyNYmGPRIgU8q0qUUP+x82CyGUCIL+viPVVbtN99
NS68CBObGetp9NNA2Yc1P7kYXBYrMfuhQS9lnPMWWhkv57OgjSB3FMTlfJDuf3/6
5l4s+EiWc/SArlcXQ+cZrfG8s11gVDo39W1K4yeNVCCxEY4KwJJbkiKKOi5PysTr
Gd8O+nQbMotBMO3MZBNp3pPECfQkEYqC6J2NRG1ju9MA6VVMA8oOWC91QTo0/led
v5BVsnV3T2Q7n/6Y2HMYdPWiEdlkkvkq8fJ+K0gvhvnfOjvSQIeGQMt6aBO3Ke7h
Bpksin+FxwbtH6RIvTqIQ/l/i2olY8M7xO8S6kHC8I+GS9MUjv/4QGUeKlWSrI/6
/kjxtJFIIkUyCIvQTRkEXeKZp0nmnJEj36m4+Tj2N4tpmKrSBXfKqv0DHhreexGj
v2S/UFqOxth5haR5r1iEnv1PGKE//aC3o67WTsc7nC1rw53r4zL6j1O4DSptbGXJ
I+I+2Jl58DF5OPq73WKHC+H+wx05PdPqx3+coDMHrWxlBOnFaU4vtXGZK3WsK3i8
ukt7hS/qTpQdBgb/ceBBAyg3AGLZbMU9oJAHuYTNw13UbI1umA8rQ6pGkdZNcAwG
nd7qS/VRNN1iz/o+OEfdj+oZpReBCAEySZwbO4uMhFt+BQlNDvLH3522pQqxn89h
QrCBSvv5QZ2nGNvZXPOdFv/ZJU+94npyPzFLh2Zw2kiO6/c7iby6q6onuisQB7A1
au4/Jr7f1NodeB8P1WYRrkeJaA8j9CMRgfv39swLPCYC/LLcMpx1Hsk51arY9/AW
1RXACElzGlLkTGV3hqRYunOE5vq6CdtHjkE9uvNIUTfvnxrZdbRHwXs09/5FKV/g
7RZPqD6Dc+du+8NAgek6GFEGzXYIv4HK2MM9T1h37ig6U2t0+tZ0rUU1f+QVu+Q5
/T6fhyE2NuyjWgQlzX9RxwFBXZcJYJ+mYTaiTuRFlf7AwXQGXrjtaMo0KqCDtI95
beKM2awhR7x35W69A3tE+j4mWDjXrWRFpQCf6Hljn2hMglanHmWBztSgZKLt1Rco
eYPxiuWOmLavy0zm4BNCC6tguTMfDPtvCRNY373zUModqhMpIfD45zeGtJV+hDuE
a6iH2cniKC7MVQnSW3VBDGcFocgQZxYI7OmrcwPEyMej+0qCCjBep50//WMotc8B
8QSnIRw3Vt9Kzhq+rFewrQdgV6kBYsl89Is2uGQbrW3A/FyeQ2k3iJuozC0WuTgs
rnFhke2iL4jzhfBY6BXcCZTp/QRzNvaXR3dB2XXWBYM7U9ibFfHh+min6lfY81/E
KoVvy5RbNYxGioyi7hw7fFJofQl6n7bmTKxiLX01zdp40FZpb1mGfXDYDCh5rPF9
X3nBINGYSW0350YQrCK1ROa3vAK5cKYqhwE8Gz51oP2palmxGNai+hx3EyOz40Th
myid0ClHukw5je8Ac4RY2sloizd+UNCHtXjgmC3kWDP1vQW/QC4BgdpWx1FbT+kD
We1Z16eqkpd2kfaeL6zOsKRbyFR8dnPSYoTKz5yWswGROriR3FlkEsuplDX1mg0q
OtLWvnXT1UU/1zZe2m4POppNVHSBdr6ikhidvu1K/DgjtZGVQEmaleT8cn5eunw5
ymYvc1NT7n4Pz2GPux5PwoaUBV4lQlCuP/2a+y+1wLV3Mw9TtIy+9cBFRMV5j/gp
oPFYI15jGKzuTd6eN4yDMRjMAQx+nXJCwOK3bG8OGyAMV6kde/diEsUfYg0g2uiS
/tfkz4pznWqZ+zFPDCK66LJM0WjmlbMgnzZDe4lzm5UA6cmFpLBPeaVRX10wmsll
t0yji8vwz318mkE6ONAUyGPSi0I2ACN7xx/fnU4Rs9w5gHJBo2YUbqAeNHsxysbI
NCRlr389TS8G5sYDU40icTCKW+ORbHqIpljmqYSaPWcoPwmqyk6buMympMwPYaWR
JCPCtdiwHgy18832RJh2jWw+OmO9jMjpogUViETsD3Jcfz+XQeP6V9pqtQAlNFy6
pTISmgYFFGshHL1BSbkH6MFkNsYcINQmXgE3J8k8UdD4i2vR5pRALhJQPTsx9OBH
gPlnjLtwtVSQAoJltJqHL+WstaZeTNa8Ma1tpTKlztOdkU52JHNeoKk+gYG3MO6M
szv6sy2t1PTFOw+CPbeVMBIwJLvoP46gIoD3515hb3ooHSWQkTFXGyqOfatRxuId
xpfWCzvYA43XU446vOAMLEnqG+PFOs1C42tU2KcgyNl+IongirYghhJB6OhDNArp
QUD/nkALwRvWey3WC8k9poxWGfkLSqLwxdh2OsN/6mJRYRBvc+KizyQM5w0ZeLBF
DTWgXVELw7HZBdOabcLEZbbhv/nF/4IdVQRAlbPpxv+UT7Jiqlv3TPuN58IdJduZ
RaMkQS4Rj4k+4H5YQsDWYXFmk/n/Q2hxRapyi/jYAmerXZQphWC+SvO4yHG67uzh
NLUgEMN2p4J1oz8x5yIhobQs1ul1VU0zN8I1o5yM0PuI0K4ibMKTC+E79BOMLsoY
RQa4Za/U57u7pN1S0jdZwXIiry1nsLK4EpI8G/8dTqxC8YhnKeG0n8V55EkFaVfd
fCyML6gUbMruOq8etM8jHCOrh8lXJWmh1RXAmJswYlB2/oP0qA6HlYcRImZrsxAr
VNUWK+LtzRBldod8xtxi5orDWzq43dKNH5wnqWYubCYmRz2fA70USydbrUpbXitW
iFvVJCiS5eKP6qWGCdkYqjWESm/X/22zzz/6GxtsRe2YOhuBYlIjaBNhGHD/ldk8
o6m/lMjhM0JIsH6Hb73iX15ylchaTBiSL0PE4hcCdXmA4aVae4XoTU+mkDF96PmU
k21HJ+Cg8FsKN+W6bn5SzHh6XGieIE894uEfd6ayGe9WhGn8tBjHJADW+0USK1+q
Xnz01rtKM6uEDYpXQdBpxJzhUhpn9EzgH/kwwHbxCWMiuOjRI/Zc0Z5x8KPsJUQx
UC+hm8Gds7KAC1DEsiWQy8wPnAdlN1NqPCeqHVS+faUS2Ig1KmjCUhvMomOwL/vA
Vs2/y5z7Y4/FbuoxJ7CHp2Q7rtnyCmIFnCNJrD8Y6EKXa+hYk/XvUJInRcI7bUyM
iRqBF+mDPGWef1A9UbSnaCJFZ/9JWyZU/OlFoesloW1Q8wYdpmQLWSC8O5P1IprD
C4xFiV77qCG64eWAmItoLdn2665XGZW4gj6R0Rmx3Tx4BKcg1LHYGTEC51o50Aqf
axOUYEaTHA8TQCQl9U/pMLn7+gvcOP7X/nxbspDynzeFLWk8G5pllTX4T3RVh/F4
jcuIV+M5E1VJ3r1u2pbnH+GxiS0AO4xJgAQNfMJ2N8L6j1UVfLvU6b0VL7M+xY4z
QvPaBtUUJpM9R3RHigHAoltSuqCeG3QwaUYNKOc/U992RMRW3s74mhJ8A99F8MOC
+4BnzhxUxGi8e7bi+S8c63J3dT1E9pQxO6IVOGyilLKvS3fIjHDr0ZTz8ILqW5Pj
9IXaAFne7wEcfymZUnPg73ZBadpvK3DHTeaUmSj4pW0VCQd7r7n07n/+C7c0bZl2
XARJN9MYF559P1SpkWLMpeBtSJb258w8azphuhWkKYLR4bjXmB96iMOmVRWd1Cs/
9nESCNRcq+/QhgKI2QBhQ/y26Yjt2Y725nOs015Yd2ScTRnZxxAb9ceZck0d/3Dn
YJ8KFEwPOcl/NsbYGurcu1iMAvZBJQw7bOiYJpZIEH1gsX1qZ5xyOGAs5bo4uEIz
wsVvh9PTL7YBBeDIMooJbyIlmxkzz5KTSD0ipJAhYvdlbNXnbuYO1WZFsauOGf1J
8N1ksBpfm1AA0hdU7cM/7SpXlvQIJuXCJClzqHTxGTvi+DIbe+smouHIGoWbaSlz
zWxaW6nWYBStTPMKiwLNuvmj4NnWFXti5BAAXZrzFWdIgO5ByQ9bzqhQXD0KqGj2
xqsFi8pfBprVPcSleYpxHIACVydgo5iJ3Qn0ArgGsgHhR0nzfQE69x6r8CClFmc2
MBWYkaBIkuPF6HDiVIO+sK9Z/3cwZkRdSxHVpK0gGMJxBRfu4EumkdDLygrrm9Q4
v6BmaHUd+RaEuuQJ31q5FqRadvku9vBDj45kODrqmElb9c+hIFStYua0kLc0B0xP
9qePz7epKZ7EVf1PYl/ZWXhm2WGUCgU8x/Al9tnMP4LP35YnDNJhqxrlTpTiMyLU
qTUvCKWun9ZZrPspPvG81cNN67Zjm41RRf6wQVYPiJdhcDGKLrhD8bu9eC7m8Q/y
exUlHw7eE+R3UVdXjfJbBEYZKmwzfu2AzG2e8tI9eJURnQ5/61B1QOnXgI6xwCBg
mEQ3Xqxvq9YoBqlWs7P3U8Mrop8kGm6FP+4NWa/hVjPP9qqVD0Ue1v6Rnd0n9M33
2DOQSyJ8+sgnWR8gf/HfEiNhU1bYlrYnCdX4NlgSA3oi8yWE6/Bou1eVcAlWWqJ/
gw05sznGJ2ZYETcEBne9FutNsooH4SNqU61bSsdQbkcO4A7OStF+///zI0LyfEzm
KytJ5v2Wxfke1x6JtMMah3v5oKC6/+P80nWchxWsT3ErWo6QpkZ8BB/+v5x8U327
fMZWUqPTS6/LxMm86MQPh1JsdHZwChKAaEtFyTkXMR0=
`pragma protect end_protected
