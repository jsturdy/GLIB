// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Klyeck4mAcTcP7qRFMMMcZ3J/eM+CL3calam7ZCTOAl4CFCKXgduVig/lmhTVGsH
vezBq5MQJN69bugWuJ+g9R97LrMtgZ7N8eDAA1adD2+9VFhX2lvkab5ZTsOqGXt0
aUOGm4AdJfh1s/dv+ZB6ygzRpE25c9NZNp/9Tkcuzdw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3488)
3Bz6Dpz69Gzuh69iMd/HWzotdghEj3bjHVvTHKW6blpc9QyWYWr/bclLLQd/KKZZ
gGu8d5YtpQXYa8LdUkGS0FxLhak27s0jZhchDYlPYwCEzxmYJh3wwTHFhsmI3klH
dIY1+z34/JP+KefcH4gwnR7TanQFPjpD7m21kvM6qRdEQPoXTpyX4qh1pSrxsSWl
rn9WqK6CROyECoFj6W8i3UZ6J1m9Kk+1LOLjsGWdXJUmznSyawKbmGeRd/tzLk/Y
gO1HCU6IPn9q7lV//bqyfimMTxQxh3yF3AovUCVtGJj1R4JyEYOYhLEOjLXM3llM
rlArYWOo98aH6osvsQ8nEUzdA6GZ3UGpzDc8rGdLE3shDt9Mte0cAVMvV8GrxJMq
1UdeeEkLrW3GmM94fzyvQym4IAUCjnWuIZLUG2Bos/JHXs03pZYRoI4m2JcHH16L
we1MHh6Zt1rx6Ftf5lm3GYay8ic7utwX1m1CptMkJwe75rjDW2wcVRrku4a1wlcC
PnLNQkrLmEQeXMmU3UaqVnLZAXMXn4CsQWCBtVx3nQB8HxXGxsEeEHa8CwwTZ83H
tn7r+Mo65JPaz0d/CtfB5XzLY3YhHoRbskQRM+9rvZNij1ZBk9LyKky/nUfsaOHU
A37mvHauugSjPzzhP2DgGeuNwP9WILSsGF0kO8uIKpyewwAdyIYid+nHfRarbtT0
A6lLSit25wWp5vG3I0zKTY4YWEfseDNpPnHW1AvwLiTH1mlzOfVwEksQ9eFG4HHv
uFV4dvg60vNkE4cXV9MZ+yGjEGZblJoEozzSl2NjkuSlJkJzTQwPSHx1/rMUlJnw
osfZ5Xf+lluM9oO7nQnqERKeOBvtyfWRzKWEeZDjsxm1EVuB45jyggSoqO0UgRtF
HlsWL8Q6sGa0m9CWBNCeXz6DULBw//JPdlb/PDZVnECFRaZ/kaRP+gI51n+9L7Gh
aQdyxUJg43RFG2pttr831ETmEMYvPEo5ZWEXVyYdy7ir/tZLvrQ6lY6mMj+esxvg
q0xgw40fMZeSOsaXz67HWiaz7VIzOMr979I2a9lHGDaj3frlL+Gba6zHTSAGrjRv
ydwt69sqBEvVcnuli3hrtbgD791c3cT860SZGThXBxJwz7YkiADL3rGbUkcTEPyA
KGE3qIGLahcZ+oXpbe+qCisd0EdVWN2PNjLP9EhvBTinyYvKnDu/BnBegzL8IO97
4j3QTp8TKaG9EbgHsuNGp2G45KEikVSt655+atg8y6tAcfgav9mDeyMbzBhEhFc4
H+NoDWl+1dACtIER5NxOZ/gVQVinseuROL3TKvu3lj2/c0GIpSlD/9JPk0QUwvhb
XBdhsgrVO6GxlhfQQR1p0hu74rahwOqVwzgpLVtyawtiQls1VIut3XTiyuoaSGek
InGqLzD3AlQmxk/Ju1R3PiLvbB/p11zy+GPURvf6Q8cqS/0iqsOj/XjETEWaapxC
gA5G3g8hoxBu0lCqn+1UBjdak8IdFNiHBBxgkASEoXS1hdv8flhro1cpAsCVhNjN
sZwIAHnOvD4XAQAJwd0LM7L8/7LKnQPKIF0+XF+lY58uAbSL/7FYuhZQf0pGN9eI
ptk5Vvq4XkoTPcnp5tqkKkm4gdDScf6U/mqFd2gLkI+SfOTlUEjpysqqvqbNwtNw
jQc48YNdRWKu3ej8A7bSS9nsCtXCJTSSWyQP1Ujww57DYepew+M1SeeK6q1SlYZH
idkY9Ztem17Aj/A89AwoCmVvqOcxYPn6KMp7v8aTAp+EM2tPNqxU5MGqQdub4nad
7q+/xzDT9mAp53ehMhOy0HqBTP9VhaOLimYLXvJvatd/TdboqCOaq3SOhNOo2PiV
qWjPiM2HrU/mnkt4MIWgpgP85Rt+2T/9t3vifBBBys9WOMOkXw8ESkoTNtEX5P7P
cqI+skDerfLFYb5aLEqI4RR042YTh+ykRvXxCmMSGp8RrObD1HgfQvBbxlbznOcn
MenKiX88kHjDLjMjSW72wBj6ZEWj+qlILlfhWTYS3EvoK+cE5/yTYFsrqbFDiho2
IjB0l1nNtvDRRUY72Wjti+j+kBpBRO5Q6yheWE9EvjCG88xTrDDNqCw3nVpxx24D
h7Up3aHn5uIoznetHiBlkgO7qsQzi47XFAOQPdpP2/1cH53+V3Yy4xhtkNA30Oe5
oUPG/EOFAqponbEhzcSbHCKMhznfXu0SvNYmWvR4WKCo87tzfSZ47+FYwre0ODNI
gdPlvtsOMU9KLLTe3dmO+Z8dPIUObxDZTNGQtJqC/AefO0j+wp/DlDRyirD4HweH
MqG4kyr0N0tBgjGuL0zYHkAxivL3XXIAN8Am8QOLWZPSkPYH5giLsvK5A6aOFaUI
QcCqEV2dUDiiC7HRzagFiDxZASs5Pcuh6XOuH2VJJe8LF8U9DtBshDjKJ2wlD015
CYQ+CQswanbg/L/yZFccV3nzLN4K3JUse55JKQ774cu3GIKIXyGL8XImAJr/Jl5y
ZYd1A1/ZPiYJkcLbwqMUCJX/YrpwGIbowHSCrUEHBo/l4lfeeGobQL20yLTqFXyT
+bwk3dwUqCiEETcc67d4UlRn52XDVEkYV8B9ompMEaRRzU21GdhsoQdYzOayqX8S
UuWp0h1oEcHjZLIAV3eaYsrSS4Q9/ASfodLZRhN0bXcTqtpT1rNRU4mJ7hzJZssk
pyoB0iYgRDZ2AzYJVk7vVivlD1TaoV7WLcQ/BXEX/cM4WWUks8uYew73ryzZJGiS
Hz58cbEwhMNWaUz+3IHfA2a3yeGktuHx3iKV4yvSiMVGeEjG08vZA6fN3a9EsxbU
DWiL5CHtp8LotaNeIkykeicLZ6XFzfHx9pqh5V42REHqB9Bm4VkWVc9xRUypJ16R
A9h82XnegoTmzlJ5eNjMbsrcoA82vt0MC1yMJ76XJ4C9UGWgdFk9XauIjjTQvN47
GqkF9U4DLIGcr1lItyq2stSoqX9QJc4jhmEgYvg8Lt6neuSiO3z30uCJrviuXVOk
IbRPVxJcRtYEN04zXE4iSNlNYbwMfC2mOzryj7KhxzVPONoN57ihdD1Tq7VHjshT
EfP3hA3kr30ypz0ML4nple5QX9odQZWu/I5qCiUpkeW0cPNm1vrLvLpn/FZ0KSqx
TtR59WLxgSvOB6WcBdHtsVbzfSBHjXof6Z9xh43uWotQC9A3YouL6Fx5WXr8UMbc
MsaWD33cVbWJ64MTn/7QVFw27+1YyEyO9Ui/XmT1wMMfUTL7Vkh1kRfSfM558O76
q0S0gFzxCxupU5JaX1QdYOavkzWE6axvauKqFJZcK3p+VDlpaZQP7WxC3nkqKC/K
ir+wSOvleRrbFlNhiOe/b9l1fopMtPKhER8uN111r5jaonzxJZbjg+OgjJawsHOw
5OOBbmFLbPXxwcREAeG7fitVFUjqtb24mdyd2y9vL5/Rj5M80BS0DIKnWX1dSuWO
OrsDrAHBb1as7/0TcDMuWoiDB2K3a9AmIYXv/F1tx9VQV5jkDW096rfXyfZEBfv5
ZVS2ISgfftIlt/7UCSbFyktvF2RLzdXBtAx808Pt1kdQnJKI50uo2zTGWaq03IGL
78rEcx4Q1nZxzQ0enaIcCDKcx8DxxnqnPqf1V0Mk+KsQu/CpzS1tSUOfZ/zlmbAI
jG1su7ceE80j2hFsKH1/VivWcNAgC8LRDMaW9l5ex4gfsmtYrVqJJfx2yPaFU8Uw
DmRmXzGxu4PV7eWf3nEZX6ukbElNRy3P9ovAYe5Q0C5U3cLZm3AqC25gLaCwaAJE
1TN5RFunfSGhKVOcm9qYd+T9jekhVz3A3mo88eptNCjLbwHs1tbKXW5ViRPWzqL/
waj0gOZQBwgb6ZmrR5F6MOI/Ug5h5Uk/PAUEylu4zHuv0XcWzuQZdvgP9+9sHGK1
bJjLb6iTToMNZdz4jw6ZGnJWlzY/JmoCiR7HlIaE4yx7CacSzjA6q7t6lfHNl4I3
jbyoSzg6tfuOQSJ5YGXcv9KWaqFweSvLEeIKBc7pF3q/hvkpCnIW/xErQlWx3lxL
HYylNPWFAkBtBVD5ltDaq1CsV+I1pZPpzZSeFKUYpHPtgtTZONNmLAFcG03KKDEF
ugoBOvLCdD3MD5L0md1AD08wFqzWmjSjEutSYl6XJgLahFwCQbAL3SzJJdA/4tK2
Dx+2u7aR3jPF4NJL/IHfkEQhZ/Fgcpw10Y4nUj//vZpQpMTcg5TL6UWV08rZoOM0
REN5pXphMMrVOhr4ZSMN45awcVHVjXbj2JrnW/fu9vpqsmkN/nsM3f29/pw1Lusd
N1eXEH9v5KDlWDQRR20nx1w/CfibuvG7akQT6Hk9wIatYBK3qK8MKWZJZZTJxQhj
ISEedRdicOB3Xh+3T1knJOOTFMTQ1Y6WekPH3mbFTq6IOhkvnoLyJxEJMw3nLNnt
c0fZFsP/5cVBCWGQhMHxWBGmEf8QLSBtVCBzyzVB9j5SnNK6JqqEWbOfrmoJJjyp
Z0nxVAL5AzVXs0Ce0BFBAeR5cMdVZJOdVxSbUJMozyle2bKQZ7IYRWuWDEE3M1g1
/CjlDUUyEoPaWyJAGZx0b5AZ6lskbLACZwVBXCBANqHCczRY7rNiVLR7+RaYjCiV
9pmK3kdg+3tzTzL1Ya/xnZQKRn6+7YyYu640xYrnoCo=
`pragma protect end_protected
