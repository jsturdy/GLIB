// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nfbwivLoFJPdNooIbsBfNz2z5kbz1dDo6IldTuO4YiK3xPlAJRBENAG90c2AJuJt
6nunF3L9GxkjTpyM/fmcyRSVqRGYjcCQKSdcBNSnSkfSoRQpAz0mPPr0TMoQeFKo
dvJUYHs9Yr/TIfdpcgEwksRrKEs5NP8Jih0DfhtAQrA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17712)
IBhA+XnZ9+7aZ7hg0xO2sf22oQauY8HJU50O9/Afoqy6Oxa4zO4noVz56C6Djma7
qgcUhXZ9vFmNeWxMI2XpLg5yczkuk4GgyRo3wDo1YKPmBeNbmtXttL+5tW0d13+j
zsPsub3vO7Cw4oFX4zhBaCigeUamwN8LCRLmrtdGzfBf78smYaTECSaZHpgj7LzK
OH1ayWIx8uy2imh3tMK34WpMmHvjZ0jR1Gq2C8c4JwqhLS9RBNrquTs9IDT3OziS
6DtKnQA0UaeoVMYV1IwPwoKHejEreoFvFDjO8PilVd54Iv//Y/Fxk83azpz3fukP
DK2tx56FLotSS1F0nviMYzxN2x5sbqrx+NEvbkPdI18+3xdNTwj1d/LIhxLJYDq5
lbtNnULJF4oZMw3c0valB30DtAFuiBufqJiJipz94gQPxXymX33tMbFPKxDK0JjG
QBGNEVP7qKGxLYCoY3d69ZG172wK/ZHbmJRcWLJm3h1O15B/glQDHTgrDZQNAev5
gbJOnfUXVtA8eWjQnfILDCRncKiL+oeGBEOvRFfAS9KlvAb/srVK3IY3ABjr0I5W
/H/OdCRTr7rG11ISwqqIcbNj/bE7seFs1GIcAwFg7wMCFFsYXZFCPGCUa3xPTbv7
wpuDsebTAQ0a4QS1dionmgLZ792bdGSyMmycxi7EnCRrrMEBsuuSsYSSp1K51xc7
bhL4VjdRz6wltsvQ+OgwtyF5Ha2KDcjZ9KQFQ7jsp0SsmoR0K5rsfZRkJjzFh5/I
9b/G3I7Afoqndv8wK37pEJDm0jr0EWKO2VXnOnLnOdhHCMxbE8Ho/Pyv2w9ZDr/I
32oI2ccibXNitFwbonf6kYJqmLBtDi+PsRk07W9Kzu6T3HSPzRQZbjGeJLcRFmTk
dHYlGu/plWehqA29aX3w+Vci6frgf5MNupofj4vRMTM+ru/psL1aweYRIaNH7mtK
DnogIbRd1EgpUJMOA+9jmT0eweydFFO8C+1XkBz33bU2HBcPf6BUqOSrpcgpTht4
DXDPqc26H7cmDF8edTRykEGTxse5mjMjiyEUhhYuZLS6Dgd1oEPiOCghJfOJypiH
U2rd+wgNfoXEGWXDBbM4Wh/T+bmVr0I1/weVbuK5nPfCWc6pCeJoap7lgAkXXXZT
pb/nCFw3iRZ4BSyKh3x1Sb7F4ul4sttGv0+PyE1aRkcXKvg9DboS7jvT8NX8SgkU
Tb4X/kKVxnqi+pNR7lbe7hUiDY8cQbZc1d+EM4Bco9SexvZrKrgfpih1+yE3W1Sg
2/o/GPyGrWiyh16w7UrN6vBCI2QynvdNn6cx9Hnkl7YjsAKOvezcwvuwgbrIQj6F
UC0pUcjoy8+txGVwPD3AmyMrmWSvAECv5byeNwEfQiMpF1hyLxnHoxvBRBCm86y5
LTKfwRIYvuAIcFn97FFwN9jCFPgbBYT8w8+SzbTDusNU02Y835z7yTsmEwVAkx81
agz+XPKD4R//s9deVqiBwS22365haZ21gnu4tfdsg48q6V5Yb6k0l3+qw+J/QguU
/vOy8+usKlm6Fny4qzN6r3UlrSmWzwfHGDdb9PDLzLjlWpjfsgXfjAGXEMgMQQtB
dqIYFVtZkev+pEndKCQRva5Lss+MShxl1W62wDm8xigRVvBvN7eNBs+CAq1qttYW
rZOAjc55KxSC1CekdVAU/oYI9SnRh/oXVWKdU3Hp013isq4s0Ja2S1iXHf2358Wr
G+CQV24Koy7K1Uv8SKGf2bPekUn+WzUXFEbw5CA5QUyPHdR5M1Cu5TuzqyAZS/jQ
DFNvtWeAlASoBJmKlTTr6P4ju2/RcLvuqaRejgM+Ba6LGuIlZ/tQjXkiKqsPdQm9
NmpIHXjjqydQMlybb9iNeQN5sVD9Pdo9b5UyZKznpEHrkvsuU6Nc8t2ZIHeWPbwD
+UfQBv8uroIOFBV4/QkD8IZS/DTQAQkivI2YAxnjMjTBWLC+N1vIaaTGYAh9YuiS
p42QckbfCbTUAY+dwQEEW0l/ooj/pnyyanOo3iB3Aj7lNT9MXPRjmrQdFf67pwVu
m2DyMSP/ql4G+4TSJMbNB1SXGgJo1OlCFy67ZVVviZs5sTfl3ciW7VH4lcO7jeu3
mBTSHpZTF/gbaXpITA2wTl7JIdYyfK0AJjpkelP655sdGKGIZPqr9Gdme/ZeYZKl
tocY8oOY9kLfcYS5bj+eNFx8wkFKW2j47jpBb5PoOJkAVCwlURzNXlxyE3s+crSi
6XomYL8AHcKSb783TcOPuMitjHBvVQ2VQdD0lonYFPOSXzjiwQRTja/pYnu7KfwU
iW/UD1Go3462u+hP3+0NKB+yocjjz/BBleo00lV9Zx1iJoEIYaalYyHFRESqvKp7
1/YIWAKBjGYDre3yW3cW+TEW0LvZho7Y9mwORIkjIUHZ/t2Vj0fm4f6VPxtqbRBg
WHY9FW7voxXDj6Gw04IbbSqGJTYYhtm2VvngrrSye4wxuw/24tTYnZpzgAG3wmqJ
pzkgptXl/2jwjptPJscDAfaYBfrPP/FevvLnkVhEnC97QTyAXxalmJWByxcj6rz4
Dd9nUksJJ7fm+ZN0qLQEbhGO9V3IPenVApX8b1djsoX1L2s6MmBRH1Mxgn3jxkrf
Zv4VYCTvNziq5heexrM8K8lSbjitFbXciywu7/vOjxapUUJnqDkgfKWg1dKZdNFS
aGOW5T3Io4QTUFg0/zeBAsCSQOw+tndcP+0LPukSqrb/dAyEaxBPe1Ew/nV0Z89q
61oQM3YNO0oNSWRirCQfqqEqrquXqXMy8eP9NYtM9nKL4JKw84yLeRVeimerR/uI
FhEyOF9/whTwp3jSj82iC2hn3M88u3cSTZETNUgw37MWZ6se4r9/pIsM7h7JPEow
houI3GFGWtZMoOmxaZludVJfZhoBDE911s82qLINwAxGoZwkcd9CP8iGnyOAWiqe
NxCOXHOr4PcZlWBM55psvybL7/wbscNXGo8LsKryPfvVyYYrtR/FtnBSSLnBqiPQ
uRNzQF4eyW1KTcfxj3jDnY6GZIj0oTJRUA5dHKy9rQdS3+6UmhItvCUBojnOO2qG
54N24BDaAx0hWZpmVonth76TuPwhb6SQ4Fc0JMjnJrQcAP0GyXuON1bVI7vh/3kS
wkOu/B5EIsvJ7qeeSykO8Hry486jfFqtk9B1gL07jQcivf59P7X+By9ulFkg7BtR
Ck/tiFGAuXbhWjoSz3IOD2wQrobF/uEK0eO5eIjyce7xpvjBIzZHau7PJd2Xjts9
PS/Htb5cMcPziW9rc1FhP2NmltwmkG1i5mo2esk5souvrpQOlftW5xny+rtsVzOp
qTmL0Vuk4I/roBESxF/u+m/xAIKRwWu3LhO1gjQCauIXFxfrQSqdmPToNx7dxfp0
XIiQzFCkLfbYhjDYnm8eOxgQ/Je7kgIG1DaOO6vEZU1BqygJHOCD6m7NEpOU6g6j
8nA9rCIfiRSw02OoUZ0EGEWLq2qF1EZ5c6O0qO1dR7wUww5uEKvwQ5GhPB2RGW1F
YicvJUWg30jN6osQL6NNz1/mYeX8exPs3ibVHtszakOke2o7MFd3iJNeN6a13Brv
glgTBaWNCInd+fcCqDaguxbtwOqX3cSzJw5fmczeoAZm+0fVAz1XaxlR7CC0iXHa
2Qj/qinsEHXiPhz/83o114ao2iYOCK/oO2LBAG/gSVNdqTIxRKCSqTvI0VnhAEON
GFZUtQ6LWB/LkWOQkX4/wScUK54smqRRi8cOwkWBRfpKBMRfUhd2wCnvR67ia9QC
RoWzyQgBF2xWuxSktR51rwhnPrU2TRPRHs6L4/6p7IiP3cWq7TGCHDH0oVaq0/hN
CbhP95pkSBLnyb+C6IUw1g+OpGGjc9OgNpdZSGG1wOoZFtqthCoaE5GJ3Md9l3Sp
UZcmNKMdzbclnyffnXabMUibqOzqYWYjWIgo17WkCmuvgQFOfC1GIqfQuIL1E7tY
87YpyutmLysNv1O8dpJHa410WPlEgjYMBCHyfI07qiHLfnXxNkigpOKYqew6pRf+
fA8z+dBfZdGOb8ULgz+8iyamsUkROyt874En29VF6ajqIKp9h7tHODnqoQv9C5nY
XJKCDlX+o0zzoAi/RD/eeNgj7da3pU/mqizifJbWktbC5bcX3P1kPDge4M2fKPps
AT6B+V3xQJImz46vMxRAtEJgfU0PlxKuKMJPv/1iJnx2Z8gwVM9OxvqhQ6Azfy0H
q7mfp2UPKyTu84sz8HUdANUpnBFe7GJQAwUuThV6KyBSGfjq/RNQ0o9VartHgBRY
2QdqTCl/bR0zm/3jV0W7tJH0W0ofrOnfL48sKhcXZ5G0QdxvbM6eKfOPGJOzeDxH
pQcUoKyLL2pCdXQ/aPkMVfh3kGwpDRE+ZLdkii7RB3/YuvA+ETn7DUjxgDntPq2d
0JS9GgMbhHqKvuRo8pQvS+fQ23o05Rm2kvjRDsFtv9gelFiiIPkCwLiHmLYZcqDx
nQPaYRj9yi/P195xDhsAeAPi0mnFtNS67Sfn8U54+Q2Bw7rLN0CfJ+yZL1bpaMPS
LyJWs1v8oWzJBwuyp9k10K5L59r+sjaxbO69z9FhDmy7KA9AtqTnvuhIIhHKQGc0
/K95a8OFCs2bFIAikC/m+/BGi90+4NM2koNPIorFDJMfH3/hX73lcZfM8Yzu5DPt
TpeEEwkezIGUId1xWWkeZIB27zs/6dJ/1n1LaThyhbTPwkXlVtm4/47Jmrw3g6vO
ipJ/wHF6fZCjqoCzACIXMvpIa6xVnQhAsWdoZSIt7+ehLnGoqCtcPhyK5iC+vBu1
Wl7CvSGraUf7KOv8YoTZU/WuLtAiV0wlWugGXxsnKw0WZZYTJx9ldCGbcNRmo68+
uEGFwmF9WpC7WJIkjqVlS16zB9Gh5liL3kjdmIUSp2/vq/R2Z8cgSrSBPzLB9OXF
fcqruOZNDpJ/BPeAgmkd319Z2S4QZ3gdnq5FRsVjGI++BxyyEH6xiASPvmLodkBU
Dxx3YS/V0SGE8q0x42G8gxcrF+WiT2g4UoRd6jiW2CPsnKw9E5YPEjJEGkmoLw7W
8Xbou3QOCQ9QeRzi8tn4rIhg588Wbj5xyrNRy+DRMw4dnLlNwiooa0QQZQdVuPWC
3NqYm14BR73NDcjf3v8L/QMiK1fxkS0gl3/DJUTr3CjK2Tq0E+F6G0KrPbMEZPq1
pNVwr+yeDnUMR0G38TWjLTjyW5yEyDVA6OExQ7A9pCfVu17qu8S+ddQ4Wpx81eZ8
uQFMhS7J4wlSNXz+95nhOyCsisW6fObe79LDQ3ZQCq2ZF5OAR09DOof4rxoPVIxR
Q8UyXcbNtHWSPyp8CE0mwF8KCA7sqsUiZaUh5DdJMW5uVSElBaN+N1PhXB3TQaiu
CS53aD+4Ki2PTTsrjZBaeeYsPnK7caikOrKp1+uqX/N8D8Ik1Zup0jRw7gyxGDOP
tOGImUu+pvNzmINJ8viaWKAe2g2H2uffBKMvIxlEGq58xEsd2GMxTQm4SLayOcWa
RtkJBUKSNJEtVTy6jXz3IBUligWK5Y9yFJUO45AbgkiM940ZmAlC3a8vFgi33XsO
KuJhb/iCm9GToYW/rPbPj2J5qMGJjtkcS0F8SsVFZqteEAamdHicdIw0LQGKI9wT
t+iaH4I9mwLbiHJhC+WFTz4baFSfwfSWcc586T/boCmUssAXJ42SZXINVQhvPVMd
FDDscAyT55E8gJtk2tmmOVNPH3zqYRUBehSN4rUYK9nvVqJmQqY86ZO8OI2+aV6F
l7Q6ReAKziSGApm5mRgIn+S6Cc4ll3Re2q0MUjCdQGxGkp/28dN6RQ/e+GckX7NQ
H6agQCl+R1p7rJ2EC2h0SX6o/xzzKKK+6Nvz/bpXRhDJi4D/Ahy7uKw70/ikBUmX
193/6WLFw9WcH0CJU/mBKQfE16Q9elvxadF0j2KTe6g+8OXgSQAgGyCzTwyLX9Km
5gKlqeuG7/BN2HcSY+8smeC93Uk0VStXAJEVn8wThEL7ZGOD05c2Yb8K8EMNUu0t
n1vuUosjM/1nU4uz2UvoVpLviWN7YwXtR7pZwXiLJFVag5cHrj+clIjBVRcMl0Jd
OT5uu3EEtQaAYiSF3gBZUxgPKJtMDoqzTQR2hdlkjK35BLei3tkkAE3+vqqYpGh4
FI/ViRguPRYb4XZ+qwD3h1xRmsaUegUiMZeTqDgvqDyI/w/1GXVDQRZgMcjXsiTE
JvyW9vZSVH9jNPIStq3wh02jKYSduwdYNZZgWIsvbQpZ8j8TnBix5vn+Xc0kCqLz
Ull80dncJTVF+Cqck6RtmrlbCOP3WYgcl8LqbV4DWCMuMjQkYDSVfhrdKAlzY2p+
UqdkLYlhuEEE+vnn/roVGN2akCPE6H6hBFXYR5f0+Mf6kztUGB4Kbv20HjEygjec
/MwPDaflhCEJU4UGkleTOhTcJHs7Xfj2oHX6o0AY8huG/b4BJYaPXmbii7xV2hnH
Mj+CIe30NTSbar6qCFMOgrn0MbCOvG7vnT6l9sLoWvWedrekNR/ZNsIHnkSz0t7P
FNBQgO81XIQWZx0FS1LUOin2v+FrHpYE5QCLAVXQ6++UlXiQo1xJru7TJlRF0hl3
Qds/1un5ufMqM3shT9uemSTkInADNNfsjfhO2qvH/lDzx2i/2d2c/KofcqFQfcqs
GfeOiHGaZdV9vmiu+IIy/OGHFUyVyzeWhtKzEXoD1hnI1Rmzqr3IsXDq6jkjrhGu
arE08agAdFg2tTdT4crp2st9+dbevK+jWNSTXDHkzXOX2PBXPALezm4oeQCtMocd
TKu3TK/y0U+V+cbaKYsLMSFn57EFZjvBJSdyg6Xq41UieaAnz14d79EOnAaUAmyy
2tdD22cZEJFB+Gv3JfHUphmBblDJE7Lff0QzMrRWg3G5oFdBobUoZYzS2ItO2Frb
6WUJ0UYSZ5FxE9PwVD8Vvw6ax0PimGjg1eD3luECsIMM/u+/2dA8kwdscDdbw/qy
COKEXy19qoWPCtY2eQBjsRTfD533GVYgW3liaPyVso4qFJgQPqsvKee3Dhkhld6D
fZMizrdoUXD8SnnVr7V5l2aU7qmNcL7tIszXQsnPuzvMcadumPno6GAdJtIfMrlU
zErarHjGW3ZijHsZu8H5WEpjPKiiG0PpdvX8j8stjWbBXYB3zqMHd22J0dQ8lnPh
39rTH4Nnj57T8nBqKfJE4eE3Wqpzy9UtajNpKKza4/AB4zaY1ZPuMxXLgugqd8q6
YcBqlwsfRI+D3d1/qBOuMiEOj8VHYHpp4aKjo3pvn+f4ivmoHCt2an7kL8lU75Oo
jc8xTQ6xBtgsHBQiVg8cXp9Sfdg1ibt0bYmy6/UmEZJeMsRmdKc8Ilqodg9xzE/0
EiNt46MCYm77iX1ndUCDs1zqGEZ2cDD6IsXHy0Z1O7zvu0Zjl08p2jRODUx53jQw
/RLILByZtffRLUBBlnQxqqsXqeTE+JsJkuI7U1hh2vc2HY+6ErldqCrNt/HzTNqp
DxYFeXEXzsCZB+QK/a36t2JsF7e/Fkv/HJ2WPl3PiD5oUdMX1Ag3Pi/+DJ7W9h/V
+JXbAuZhL7iaM+jqMCbWaNj1ThN6WDjnUazcG6U+Wb9iIq4nyf/ElKPEv1F4ImAh
vk87qoQ3+m87iTsE+BxbVaOJu/CYw9nJYlChN+//LUBWA+f07c+C9ARnWFgVOQu8
LnS1V4sYeP+g1ob5SmQ+kWA8Fa2K+v6TJukb4Zyzbf1Jhr3v0ucj4zr3jTtgbE0H
k0goeWEAFiIDxPXeUaVefyrLhSsAzgb7jPDAKmEV4zkxHxfe1rxns4CW9S78CwOp
krtLL0RyoDdFN9DbChi0oIvsFz8pMjpUy36gRPIn6cxH4CwF0D3Vop6bORdT45Zo
eJaAiZ5VqRfv3nrjW4z278//T36bjYt0OG+lYG6ycMo/g7mElVt1bPonS5GZ0DWe
b9Yr8m5j3oDspG7Rgjv1QSiTmu78ae5B3xwieFV0bP0skbPwJDQPNcnW/6VKOcmr
DoOns+es/22gCeaIvougBKy3gQVN2oOfsTYNQi4nwVWl3ma339eSOAM4+B5c7xcT
aGqiCHO4S0J+CQMtyc2Dcuuq2PwLwpwcp2scuiPwTndf1sLu3XKwSrHIdOd/RRjq
LoZI/UEiISoFyLznmxaOCNuRR7T2kAxl3VDy+mYYNd7tCkFcbOHYnaVtlgCaIBwW
YDLpR9weF8sMClccRQSTmbxT1Zoifo7UX85fZOsvWyiQetfmnqJmoUVCgV0C/7iA
1pBZxRtc7zXjCI1ORFZuIw3rxsXE1DXsQ9wQNAwtW50mg2HpUO6byW6Gbma1GiOn
2/6RHYe4c3IWuLic6g5h9XlqJf03INc62EM99ZVFUykxNI8m0BPa1ywx8fxtgB6o
elpJKxRvYUHXfMOieSZgF78FPxyHLXr+/7T+vfDUbfz9cAfgO1gcJF9CLNP0MLcl
YdBmTyPSxikSWLRyzVOv5xYV3wzwfgf0HsVsgcEmjl5O9VD9nUPdLf/jJMAtsP8g
26OJnVYh5yGHgxz5eiGZyfW7XziXwEol8eENDLeP0BG4zdk+0Jjc3SvBVsMqEeox
C09KWH/Ca93PHh+bY/nkg3/inTy+NV+4Cx/y7zn2m0aOWCuqhR6MpY1dX9bosFcw
wxlYnNaUMf3Xl/+ZpKBgThVy6+RDyRY9LmkmpMbI2k4CdFpDUCuaKILkLJvpHNrU
eWtC5ArqQK74cFDmHibfONsSd3Wmdycws+6ibf2czFncWxdDgwoNP4DGiv22Xl1k
IhcRo03t9bYAol1gsoajHGjd3kdJK5huu8HYyer2cgACu3+0y6aHeg2PmhNQ2dI5
lYGCJNQBRym1MiLlRO9cyjs9wDvPKaYGqX1j7BXAH6tGUaRYko++xmHQbVPzVniS
gdh1YfcReG5Jg/yV8KS8r9c0H1iAp3vSF9yLKx7SeXsegiSYIdPnChLrdvJyxXf6
nqklSmdTavefhA4dewFt+EeH/Pfk3fK3ZEUfNzkCYbzXuTDbNvOpfCHw+ujfT+0c
kJO1rcZ8Jpq3saVPDwubofVPfb6vIYUtOMMYAG9lTvpZ6bEDadGbtGhHkHHxHO8m
hwRrNq4644VLCD0akgB1pg6N5bilfuGKV90wk27r+tZx9t5O2c0fENs5LAGH/rEC
G7wnpMewr/QB8kxDhG9a4eIskMBWF1AbzIzK9wAiJEDDUyXWMjsxn7Od3ACEN+I1
PGZOSp/IGa0RmpkiIT4ZToamGhFmawmkXQzC8A9EQWGcbX6qZkFWpIZEIMxS8KrJ
r2OxPaol34qa8a3MVGvPukjpekbfAnB852iQp+oBozRTYAyxZwBbCZU3R53cYiVw
IhxM1vCFQRD1spp2beMXcs45c4rVgqYscVJNMpUCaK5S2WZlDXLz65q/1YtBi/GL
RX+byMs3jlfB5EhJbN8ebBfJT6qdI3zrhtKL5F3u3Z1RVK2NXP59szvSB5yO6nuB
+m51ew5m49JmzNaUPAN+62e0sedrUEkC/pn5pjebG4iLv+Q8semr2hTZkymV6AWL
Ml5reMMTt4D6/SWgSnewx4+q53gL7PihnMWKU3oHJ3d3dIMA8xRYbj4ltvFcuKQQ
xnoHMOAqwikG8ZyrKgmdRrdzxpi7cm1n7x1iqPYS82aASj7ZL1a9WW0h/K6iwA17
rrkOZvsnsHNyvpS8bXBtCw3wVPtXZwYQhDvMaaoSjxG5yYxeMCDZNewKqNwcYSA/
m2ZYr4s9YiGwN8Xkd/iewa6PjD57fd7kzjtl3Z7lcOEQgxzDqq7cQ3TZrGs4LiBP
9xVP/aUOB6lphZE7L3Ro8i64wiFA4D1AZxRJth1as80bagoIvjknxdQSq7en0JTo
PkpFfk7K9jbSbAK7L2Y6yEQrf77dJ0WgzTq2xrsu+c3AWIfk0f5wKhfFBkDnNVuE
q0tc4qUXuymlB6L4BJBJdt7sK1pqzASzDd4/HVbeP0+d3uWzaLlnwW6IyIGCoTeF
cdMJtHMnzj+e3BbUU3GzI590RIZJOFEcrOSapGItq7N3bY6pyqcsgNKLM3o4dZ33
N7Yvrt+30oSTqqP0dNBrn3nRAsvxLrPHTqO1zgHSE4Vg/rPBbG1BSol+zHK2WFvy
53r+g3uHzXnwkzzVHNysGAlK5fgIwlzTIQHlLZiIB9DABN+ZM99KL51xLGB5lWE8
ofyPo+QPa3Q+7EzDHl34DU7dLauCqCo1/5q2uC93hIaPObenEHgGq34A94HyOv2M
RrEzt3i0c6OHTIe1Dk1lTt8TMHoTcHPeQ6f5q9Mnm1Gp7MAag7ZzqNsSwzfKo9rP
9XNW0JX+Xvnele6cr1g7LlvaBB992MV7XLZvZIGY4vv2Nn6IJAXERPjs35JOrPeb
IoLlY+S9BZglLTLSQcrsy7UhBVloyQTQtAlp1Wao5gW/LMB/w2qG08zNbohYSq9m
Y02pzkk/T7CGyrVgJmIRQBKvOQrrwj5Kb6y0uASYkJIBq6UnC8ZixfMz37jisVv8
StuF9M9iXxCudU+M9W8rT4C53AvD/CeG0PmFQf6Znul+dumbRNV75ssnKiBdbZKl
Cd9qaF/Xrkgq8t+I1LDSVtd/7LQveHjcJNEi7MqLARVjh+gSnartD+RWC0mVazHg
mycEWKrkMmtO+Ul4ddha+eRHxBdZMNxJ1Y2NGrL8n/H5IVYsJ1ewucOr7WtdP96o
rKrJ64u/eRP7e38dAP8WesrAX5rZs88CzQYQcp+9Fjht1ej7jZ/dtlTKyBFqnNwL
AqhIuDvB+PvWGyePzFdYuoHd2imDxVFPXeUTZMwKZWsSWcA0eE/QJri0bHREc9Pf
+7eDORHSffuqoFqA70u6/n3eyByvS9Nqj6sh5/J8FOaoQXJBnAkGhVbE8xnQSz80
sBD5Ve5c6xK8LU6um4CoWHsLz726HQ1CLVosZgggQVAZGoBU9lPwHW0o7XujAaOr
mm1pQMBzO4x8pL6UAOm6D/jYnyVEuHR0XOpRUHsWjyGdlfRTORDS7PXQ10glhjI0
PXQOOyzqFssX/T0B9EUI0+sMz/cnDOkElEIPOkbCN6pG6SDVMuU+A3Nksu6PqHwb
rpSOCQ0yS6ttgTEC3kvnRxqqoJsc0qsSi7KXXiHAIFkvffmLwb4Pk/nniqh5n7MC
ZMhnOSovrJYxwGvzzW8b2EzfyKKp6LmesdLzEXElXa3AsEbqPaUCqflgbMDKRyR2
u6E9UWYZUnVBeLeU22F0rjKYHIGYS4N3lotJCDwPcAWCSUsCb7ZBDDhOQOzl+N0K
s2rm17U9qqc25ByYuImkPdyW7QnM0XnFASmn+KjqXwjH/iAmi4XQE+d9Tc6fqruc
gJDqIv3Jqcvn8XEhOit4rblSstbzKYJ1pRMuiCM3XwakMUaslgJM/hOD4S5PcvwU
t/UrOW/9ErWBovaVvXd49kwbf4udOTkgsttDmnhm5PZ8jzMuK31U5kFcMGs/uLz4
AI6ZYoIK+sbkhIjGvv4THj83paTU75f9dDx9kI/dC4rSYzA9D/D0LkxUqWPW4Xi0
MiQHURNrXWDUa0kboiQLqXFkXoD+kHiF3l3P620uayXj1KiWV1RzrFYAbHuexxOt
c4zZK74ehMfejYmicIyltnObM0C5HdD+VHPNsbLuLaWRnfjbTFVuowOkQithVkUj
VoJWS1hWM51EA53P8p+JQAy/ij9Xhroc3pSDLucqICq0EPwlJdSTMsxEvKyuynyT
UMePfRttoz/Atj++VS13oz4X2U4Ma6ixvb9JZJz7ChEW2BIs8pdbIP0K4Xwv9QhF
sHF/r2IqZc5FZ5UEps3xvFf7KK1ihmu5hJ107KifySfWkG/YkydkFC7IDjNEjpY2
90/0/deorS8GtSJbGMUzIz907Q2lUEoMnNF52rbR2oFdOJa/ZxHCCpr67n0pkz8A
TVQbx6Nr5D+8acfNmn7DVJgpt+Q1Dsub0e4JqPHZ4La/AgSnpoDGGVPGcIqZM/yt
nDpZKyIaVtoeHCtMCECZhN4vESTP1+x4N5XnFb26QSbhmJWgptkJ+IFbo/eC2kGB
Q5GZtAAT/QpoSymU6I2GWOvPRo6qd/gQhknh4LbZ+bjMgtQjuMH2X5owLXbC7yqY
yh/OwTwPZdf6Wjj/GDHsSpaVVY2MX27xE6TDd73vrzLCJVr2SRvfHUnEk9qYxTPp
DwY6i1mkjMoGM/7NoQYHRL0kPN1Sq79GcEbpjpLQ6M2MjTDAhfV63E1QYse4MXgm
J4edw/YrBj2h9nGQULdrHgVNeGtgZimL5Rb1NGcGXmO3npXCyuQaeWbbPH9yY8Qm
a2Ka3MzoqT1t77QM8Fmu4B75Vps+wu17h2q3ktBu/ELWSyfHSLxIAEgTpVOOyrL1
fjsuBSsXL+o1zMnkOLFFQpy1cqo8857hj9OrC2EG6+OOf/tLo2VmTTm/d5cvo11D
nIy+4jBJ7wyonzc9Ivl0ACfq8lz00WWYqV7lS2d1dfPkBobZoelCPBQdxqVWlrym
04G8OaAC/dmhP7Fd0fa5G70rCry396DRVrev9y7uGbC86I7J+bMNwsC4wYQ2n87c
CNpFdZgWi8muWGoWZTjPpfDNL5cZ0qamG5vDHzdznJudvnSUotbLTZ9lPUEdmWd4
QoOpRFVqUdjazZCeLMJBLKcEkAqZXPGAi15h6t0lWUwGAivQyh4LMV4gGXU+kgvl
78cVI5hyXbqXbshGObzlPi0QsVp1Jh6PeabOF0Dps/pprrabP80AS4ZZ6UK8Hiat
QHEvfcE/4NG9WhG8qCn4oJ7mDiNTLwkIAEG7S1lpPTUN5lszj4nnr+xmGXm6gXXN
3p+EzFa+2tYNTnC+abPzDGsQryQrnQssbXLOD3senb8ZEOnb16JWBN3xFV1EnbA9
/MAMHxk3yDonCfL2irwF7H9GVKDGLo2xBBbH7V1SbcCPRCqVXr9JH0Jzt3PN5MmW
84SqOndBqqowQXtSX1dgDSJhtnTec6WYI3CmxMAeu2Mvs72bfcn8fMLu5V1frWYt
XUFnOI12g8DF6tCklhlF+ruFH72bVf77Vcb/FskgcJozMMA131KUb9TPheo6FRH8
FJNnohrETWTaoKRtnpP/UKKyDvVF173TluZYgDb/M5F4VtIbCGcs2Wi7HoNSpKks
k7TeYt0Ttcm5TLsNYEfnzqpevxzFiaoh2V9nh4+HT4nlqHMVnGtY+BJoCTHI+MwY
00M7drx2eXI8cpmu1SHtTJu4hKrKYzjRaDljM8Ko5eoPQJLUO+Yf+OPRsXjyYsJA
37BwFtdT1kKbpW0x8YwbnD2v5FtFz6AMf0e2yB1WtFom4OyjKl71BJCKZxfb7SFM
ujA9r6Hi9qKCaVsenuaQr6/r+HHGnmu9A1XPXvBlehj4D8FaGScvfL9rSsqNht0Z
XtgF+IOPC7oIXx2fIoqHxF3Mpzyg9LqYJVeTynn+D9fI3NENvwOMIXPfksB2hhiw
ecznWQklC9WjOGY/uWuJ8//NsDxgQI4yBjK+kTyMahTfnfOboL0u7+qRZ8fBsPem
jxUoPuAiEKQKQ8Q9BWeBwzT8TPvnACektTHkAlhVYiTRod1koS4bH81khZAYCN4P
Nw6hxkemJg2lr9fgvLWUpZ7NIibXxljJJ+Mh/5VS73GvTxVaDarcx0FhQB2chxh/
j/uBxGE3qsINpG/0FqxZWWwKvPfZJse7yYYGa/G1AkpqCDqI2bxAsZucU2G4v7wR
DzZtGVQr+tB56+ZSjZWfOjUqi+B4Z7pksiWBOELc5zRjiFJnlMc47zVJninD+xOt
8lU9V3ySgI0OXdkM4K3mrMZbPeactCYgWtzYM1jm3VinIXpRzyG5W0NQOOmblts7
ne5KM28hv+BsGuYam7NipGSRer1lnLn8EY805lBXd0HziwDn3CZxlsslUf4sxqQC
zsdSZ1Pg5y4a2aRgBAR86IhhsiSqtFYcXDso5qv5dQqSThb8M0mJIELGFJpk3ABo
UYrfcZe8zV/cm18aqChPhtHlE0E7xbYUPetfdvhCR1DnPuALWSwPCtrTK8b1Kttv
alD3X96SNv3aZt3stqNEC4i2eMoiatxaIcGd9F46Sb8majo827jNMQTF6HFvh3Ys
2xkTnVLbbBSM4Np17yQfRHvCUChu8uJl41SMdJEdD5xAnhuL33uQgWcgMm34rf/t
G9Bmys99Hd/n5bMrRQzNoTAPNXdNn+68XuKSVHPoEZ52gqWFBmkf2S8RnBli7O9t
jl00ikA0yv0CWMAqfI1+YjEb5ck5QchDyRdUuFVL//ZrOS8qmV0UXm5hnKnWc+q5
6taftUFUGy7s4cnaX8Zu2swVDHDDIi7qbYRv7C18Xb9Oqj9kAe0oKqn3b0UzM7gp
isDHGUQ5VsvCYuh39jfPis3+PX6VKd9kE8Iem82lNxkYd3fBowLVeiZRA4bMlgue
ytlDfpv10NOVE06icXKwA/Y6DbmqH6m/PfmWIGeX9P8dkQKRmtRwbRekWOuk0jk1
aQNQOg4YQTLRoqXqpxSWK0T7ELh2qOx6hy/txlwfTnZkT+gVewGvhrRfTBatUc5S
QTeTYYh7lVn9+wYV0wbJXJLOCigf5N3OwA9hJ7abltQapG8VzjK9efJl3+0QW/e9
4gQ7/mKbQ5grJ4RqjQdWVwKHBWhUEJ/EbKV8jnL7AQYG+C3XCj0Jx7/SFg0CGMa9
lmB+5O8eqrEL//bVlqBaHUvlmN20YCFSTtafe+hkJFxxcqEInbRDrBOH3vJItiLb
qOBDAeSQG1natDoeBa5QWy3B8bd1Gd+8tKW26df8V00w9psNoFQWyjLsgP0nPPT8
+ow8VrGd47xA7+1YBt+UNzhLIzm/FaGeJo8LR61CT78NNHCO4/HECkINS6k0SNXU
9yqIEr1QrgQi9TpZn5hvx4y/I8LeYCDmpP9nqoIz6GuuuHZBHWj7HQoifTtoNfGV
GzZP1UIdlN//lK2qE3/JeBcpu9qhXnmdkOr8H1JIlmh3QbXfvmXKBzR8Dv6Ubjgx
iBF1JOCElUS1MI+6bsPP+AaBXnLEfIcUiGbsulmCJ/hGnEYuESRKrPeDMxFr/uTp
/dtqoux9aAsJSqZRgimFw/qJb8UeY5BkiDt35HjA7Hye+yBrrLLwE+DWi3tIYRvb
kmb3EnNUczIBNn8Bbbe0tOb3Gd0gryrUD486VaUklXxp5GNfqoKp1TTvdEMtPU5G
0JdIEtnaHNE4aMMaJdnGQ3JQmAhAdO2umjrtY6iWelVy+YiAH4VtFU2Re90CyPM/
FH/RqX5rzwuXSbhSKWBZkJPnaktlQJv0YJgteVFIggieTPZrrV7vKvlOv+rie3kX
GItODRsLmZBjpZ/Wc+xx7EMaAjC6tawCyLHuMrMRXaJpeToaRMcgSuG7OuNoTDGg
kVe5W0MU0dVSAAl8qNzU1A1duGARYZj8t8MBj0pITUK2CfrRIVh+/ZwI5jYHW5VO
J6oI0bSe4AFnMuGO4jXcB6zuEui9RAyE2O2+LlIlvVMvzyK/UDPEFCX1LjTydF6y
szUA5LNaFHTB0xL6e66maPOesbmbeHPz2tewJq0LbYG3H8S507yYYvYyJkIhjtcF
kBwdeHaPPjQYjcd6xuA6mFYMq9M/DQ992hmuSq3xDBeFq6QvnkcNq5KV0lsOmy+q
HM9wjKpLGLMqC0etIKnIlxzkOtkrTMNb3pzzfetxFlJ2q1uA3usTIpSKlLS1LUFN
rqb4ClBKDTNaWSgd3gpKir9F8iikKDoSvjHcC5eepPpHEBPq3/uEWnwMin5rTJpL
lUsNEUSW29kjIRHeaX4xR/cf+xmG32z545p2gXFEWM831CAxWrsnr9tkzh8M+4Ov
XsNGzBwGa6+NwP6F6yJ6k7Ze4JDueB/n5KBVdvZ1rSHAjodMNAF2fkUYaiOZTUEE
HpU7W7diReQ1IXYk9ER80DAvAz41WcArfoO4b0k/IhO7fZWLh3iM115LPvCK3xi2
6UToKxiZt7+fG+Laptxs1XjxT9tDa1uER5IwEswOTmQ2RqDf326cjgvimycv4hg+
4ZsafHqEaYwIpFFyuCNhkS3hh6l/LRtfcuReL9I7gVm734QPC5aetEnR03NYey5n
l9l/d5CUDdK0RU0E8Gd6l/zNvHeTTUzX7FNKipAJ5bhDViGy8SOHgpZKJh2mYh0B
P3pe9hsy9U/45aOLlP0APAdGIfn6qo1WANVTMZ+exGJPEgyQpexx8BnVxhJsoR0e
0AQ86Kx1UQ/sDYGW7nYD3UwPTtd90X2vBjMSRsjZORWGSPVMduzMtdUWIHJ10zxj
BRPYuJmMoemOE/h/bEjzrLyJZYcdbEZWEcwocEjYAtV7mZSmIJkMw+ogikAdngFh
dAbtnVAjeYVjgvSSlGqGd8X9cZU5eLaSPdxDrx3fhx29ejU8SSCA5VBwXxZ2zEht
yKjp/dOBhMnUlab2HFpTEiCNtBqHhwZ6t1dqNqvhuQ+k5fQAKiN7AC50W1R+P2Qr
eSf+vTb/s/UTCWwqaMZL6sUZnwoTNrb+/jayQcID4ANtiLmVrOl+jG4pRn4TWBQe
vsyKRNVHCLAERhNAmYzm+PTphElKJOcbgf0nEK2uYrtZ43YiP/mFJj/quo6Q5zQp
HHKTcxUdZEqvWNMKiGcTbbcsU5Vx8zczLrw7doWDPgXvb8GhuDMb/pCM+SxtG9Xl
ep+FRO2oJMIH2Zb8Bl2YxWtyZrlfAw+hrrUSx00OR98SdSDsU6PaBIK9dYOh2QKK
rl7hLC8TI/Zz5IWApUIhXNucrb9uV41Ap4iOPNji1lcXtCaPu+diLsEZTi/g4Oeo
R5XD84GEE3eznLTwV7A/50Kdjt26kH7BMu9NiAFbBgDXJIc/k+BuOS9U49/jXET3
Gfa3YNqtWCkOLA1TFhH3jDrcKtJCJWWnWrVBf6Byjm8kU8W2nlvES6PrSC3AOzii
Au8LkMxNC1f5XlYEqRPFGVI2PeQuEq6iTB7Bujdi1xZq7dLYmoAEQPuNOsWUCgDx
aDsINJl2ndpDM/G4mSjgD1WfKcXFq6ITdzSOnM1A0/qrFfHdYky6SYLakmFIz7+8
0Fh7vkAQzxqrjffqYpTuO/gOW+46BtnfqGHg1ylqdaZzyTZf89BfAmUyX9fk1H5A
fwmgTHZbBF7WRX81w7WolgieFgfBDLcXkjERaTjSTCTQXeTHNMU4iEMfyhUV50sH
ior+Xt6tlNOofSCPjhcbjn4ft3ahBNJtcUYyFYzpMzJ1v6AbHdYF0YJOOulLINGE
cu+uZWN4nJ6AUTKjeKSM0FTj7V3NLi+CaVopy1gwbcmh50dZgECx/hzON4Wk4Mfu
jld7MUCQT3uqvUysbCFM18GzEYEvHZsGoLDaoVhnzUiFfrcCf28vcVdu0/+z7+Wf
zPjvIpvTjkHTAAS/iiu7G3CmpWVDRSMo42/XM6GhgXKNjZCuXeuyqplajjJIDY2E
Ow2kZlA0ij5t2Ws+2FyM/Y70Z7lMRO9Qvf6pRbDxhN48gtijGwKjtaqlYIIUiKJt
In5lT02slD/lYyux5byPjthJOMXrryPGFNqr9S0/nwuYecAbVURoJBldhUj7qCyP
xyGsQbaPk/vhaRv+hcz6iY939rWLC/Yr8/F29RZYJU9/oxJhqDZnkH/xczVq/+YD
+V60cr36YFhkvJI3Qdtf1l6v9mRalTp1suKk4m3S5OcD1yaO8VqaIyGB4Qcx+fkZ
/TktlIsrMt8d8XPbrWHLKj8ff6cgI2zayQqyPFueYFHFMhBGMvdFoMGsYNuygPzi
yvK7fHQ4oE6G5P8ip64y40bzKIIk31RHspVCg3jgcuPob2e3u06J7vNJ0MZaCqZJ
4GqHg8PjgSV4Be4SoGPaVVu4w91jo7Y0ezfeEQjEiLmo5XZmPBg7FqDysyDHOIX7
i5RtX5wlp7OsZQu2Zox+lH7TxAa1QkLZ0b5V2YC3RTJAme9YD2RyMeFYqyLjSCLq
P9B6mz9xqRUyLaLdd/Ea5GfbShrU+ZRA3VKCpHNgFJJPa858BJerQ9O8aoHmkq/b
C9JuVw/Z6D6iSPPDuF6ZSC1ArPhwuLqR7nWW5WHGePc685xf1WadDUVPleiNxz8X
p4DEqr9Kuavfdqdc71uGkRp7lGa9t3oPRVnUdKcz8H9v5Td3oyHGSn32XO4FCurQ
LBilZeLko8KJ4QXPfmnmR6GFuecVvWInKpCctcSkKBA0a/anj/UNNFvDA0ndw4sv
SIlF3nBhpF79cPX/U7sNhRj/PxLxW1gpUk7Tu/x+ibFIQs0kgn+AM4fdo/6yxO02
T+85Fpk0eMe6EcPSDJpIvF5W9sD85R+vOwW3np8cZcR9Oi1S5fblBuGVGWbBddWv
9lK+fhc5XocTVuAonNleaRB1tkkwLqNsYlaWjUxtd5LZEv+wcY1qNK+4EM6M6jnu
C0oHinuYa0pUj6XOTGPGp0Y/YlR9/7t8hdUNQ35nxhFgPBn5Z4pj7NjBB25zAhaJ
yXqTMUaFdUW07CZzRGyd9o/C+tBxTgXJULz2OWKY0CtHGnSAvJfR9/zbcW07ZpRH
5jsJpCJDztDejTIihDUilB5zFKvumF2YDwOQf9igXgZ1BkoquPw13jDolQyWRsG2
GKkKFRfTJ46+lB6U1MF06YRqKbJ1HipO9wf3mXhjhWbl26UduOXWlcv+C9mcRtUj
cALIEzSh8n7GhUk+qOVKHgF20Nw19jEwhZXWedNOEppDp+c3M8U9RfvrHevHGuSo
g6l8GSDrvD+kWYPYO4z95TIOEPmpI1vVph/V6wnA5YShmvsv8O3YlJytJaoyohwT
Qh9wcvENgamPdED0a+epxI4zitcbPzYYptoI9BniQUmB64FsHgJ0Z1MGOSqpEJH9
kuRYoOx51bdZSVR54J/XIne5p7YJkLJR4EgNBDh7QJCI6ntzFo+uGjURF/eWJmdw
D0LaI/uS3OQ/6FjM/kcYKrzh0421w8pK2yyA3sQlFn044tFFLeIak/fjfVbfkt5Y
k1aA+sfvkubOwlv6aQtFuUg7f3F2ZncgJhoqYqAHer7tbHpjUwQ5xJo8IhpX9W7x
IyiiRDWDN2Xt2dK1tbxex8pm7n4zPANDw2tJRnk8cZWz+xrUarxjJcqct133XCz2
TjH+ETa1M/MMVNejdiJgblvhwBH3sQxvB3782ZaTLVyYxSfJCAATtoWKFOj/zpQJ
hh/LkHiI85Ye9CSr0FyKzY/Bw1W9QF9rhjpyoK/6zYsapfaGiWM9+CXgjjn0qPid
njnVsNjkRYCOnKh7ccm2j8VzDhB9S2pwLP1OAIEJnumt9m+WQiQU4t4KOO6yXPy4
vKvlgYGGCEuADktaH4LaJVbKt34DeMV3ldFEtMpSKmXhZjgTs2f6bi6fYrlfhOKU
cjODGDh8ow913IgLGzLe3wVgCQmZXIq6fLoKLCfFU4Mnk0ORJSikcOevnv0oTUhy
0vDEQUxv8bV0VpWYFjWFkekyDe1woDEEnC+bmneWClNEHyfdgo6mmFTm1vWtMr41
tCddMXIE9AI+deTNyEVx3gbuUQZ10YWBnAhaZK9V8Q0xgyGQPX8lg1zZQ2CFeg6B
KlokFq2sO0re8OHhlHz+uwKSAc7x6lNezJDh6C/RDP1E2pWQRUorKFCNlgvAGsF2
XTd8WaV2BZGqvD1iJgaerGF/QJTWtSYaemHvcAxcU5AhELeXOTWv4pLeBI2jACiV
K3lz6SWTHNnEfy0B9g3M7//YM7suTaBzdxrw227nfaSdoL98HWB2HiPo/k/v6wpP
0YoJQl33pxt34yZ6Oiw7KggVBwRyd0+vj8txWRg2LbRnzMdWzn+5Qo5lTq+Ya/Rz
h+Q4xGGVz4ajBBfn9KpjfK+cpSXYrVcGKrBRKntzbRTkyvo73ZIpEhRlQDCF6gC+
PMum8gHBx6XZGpTZhuDCc1/MkEBOP+5YO0smG42Nm8O2Yc9Y+kTGzTxUKTtVZwOJ
aIBCV2aajhcaSz2agWEIkMz0ptprcwlNinCendcqeZh+fPVyLwJf6OBkh6GXqPu4
9DVe7jhiI4Wl8NqzSZjPOs6nXigLHhSwOnr31EpZK3C8imc8IJ2BYGR041H18m0+
HZmeq+LJiaWTjTxKFFgNZNv4jQ7JhXAXCPw7tLOxqLnkt3LFS0FU+9czeVaedyY2
RpfgdLhUfiqYZ865xcmN0jluYbt6fL9RTbSAlSp3I0NWwHDPCu6fBe8muSABn2ZQ
J4E5v/LYTPZKyNtTHe0SrTAzPmy9iljX6LybY4bDchHUt0jG3uSB385oVMWst5eb
b9xHPLg+W+YOO/CBMoWTcW3gWZabpOz1SfOkbmnBJr/sMngBc4mczoh3OiruVrE4
34ak11Gq8LO4UCFyTCl1fQzf0QIds/sVHDiFBDLK+ZeXtlsvvnnsWnC6XWMt1yEC
kwmYNVlaqPGF2qZEIyjRzktl4OJq4yrY9bd+8KSs8xbSqrj+TBX64a17uTbBRwCq
lFzqIfKZYIKCio81zTVqp4OssK/8+TR7TR/VyqXFFqmHn1Pmy6nHIE3Sr2+qpPTy
pH9aapdCFxcWPFBmoE9quEf0xHlIf874t+Kebfru2hTVCiBRbhmhEY6C7hf4ttrT
e+QPfmn76pJ+zC22i6UdAQ1w4ZPfYjJ65gwRcZTfz4uQCHEwDLZiGJ17MHQA+s84
B3KwZVKF5yQoSWTRQGXGUhKz6bfCbrMFVakKUme4ySmVFcDnz91oWCPqaO4T0hvE
NQ7qyoGpADR4Ibj7NtmTyFtFxQkZnRo7ThGAtVCiTU1GeMjZswqfhJHIbBbwUd5b
Mnh2CS0yP87wJWIN8+AuiyrpjTFT1M++1gc00VcuvAePb1devwV4Ki3KCTG+jAR8
TTsdBks+O4UufK2kVN1Dlp8yC20h9TZW66IEWvmT8fke7ge04Z0Ot4UA8xA9J6DJ
/svhwdEGdBFxY5v/hWQlrM8r62QewJ8C7MeYQA4uuPTyk14y4srunktGBeOufDtY
4jVyaCx8nv8F/+wcWJRyS24W3Szvjb0/GGafVb/m+k/1zbbvQdvxmxgQTxsLwBtx
z5NsMxsHUgcIob1XCAjznsjlduYimazxEdg6z1Nf1szU5eJdJv+hQhMm/Gwx8XT4
u0nC9FeC4hwsESmgpzQgPy86MPjy8MKPe8tSqw4wnA6BuHlB39SjfgkWJnWHPGlV
Awhce5xsM4qSqbWvfg9IAda/7qWAH8R6UkM0HELcRzMHYQjnT6b8/rT0u+ZCjb2d
2AMRxtKnwwHYOSKiyInGDN9ohHgUCZzQYGYXHQdMA82EvDe5Rf5bvZDYmq7tmf6x
QfN/0pIfrAJaSpDPgUbFyvrCm+hBMXlZ98VNwJuvW30FiAeeu2EgeUXttvZWck0Q
ia6hYgzCSONsXG9V5PzK6gmGYITITd17X+3IMdfwnQslA43SzzkXoG5QIt4O0885
56XmYGnHP0H1Q1cEQnaggagOm3M4dj82OEPPMjWD3BjFH6mDpG57X48umFKNtBSi
n8b0TapjXphLGG3UG1fFXjik/hB05o+thCJGYhTC0mViaY028HuZFFsu7rOStAnP
yaEDR4OWL6kk7AiukShEACVokAylUQYjTHxq5n9pt4L9cI5zmu6vF5fw1EFGy48s
3+iUeJLbL2hspU0qKqhOonEPgQJ17w3Ffi9FGp3qSa+KFz8ZlJ+Q7xe7lloFjPU4
Skv4EQ0AAU+UBoMHM1rqCibaKh6sHEEk18oJjOe4fuK6PwOZqYHh4Ss2HsKm5UNv
dUcAUn7Zsn03KzYzQ38dKzWHDhwvWuoeYACpMthd3Qut6Bddzaj01/ii83mbZahH
k9eI+s94O4RNEXmmpgsLq93BHGyEhRnGjCa0I9zpYz+6g+3PospjzI476IKUj8zk
RcoZjYLYry92pTEcSEuYZjrjaZskjgWB/kqDDglaebk3dAQGahls9ahfWg/v0J06
ixikDkBvdyThLU8txBSc/OGiS4wNQ8rqt1col0GiIyCXEe3vZ/SBCwIGB8fG8y9b
zh/GjIkw4BXQWlXoWti6weTwWiYHesxxC/CPZmtEIjMVQq7Wq2RFdDeUrl2V3GI7
zEsJrzX95bSPIgMRImmHAESeBTdSJ7O9wRHmC2V+Kyfg6Xj/l9HuBkmoyrZMz+2R
UNOToXddhoYXmE5agQiqCjSd5UqtGOx7PkoLRTmdyMQT66YA8WUzT2mOHvaxnhnv
w7ev7f7vNorHNJS/YUA31J4ogpayqpG6Czq85vhS5k3Rcm74Hhvz6FVj6v/lgiiW
wQCfeJP57ARk3/ykoMxPWrhUQTYUeWoi6zqwkEiX+08v3zipNkJPwdmc1WqMqohY
iNgQSH1MS72eY1gZNWmOSwIUIMARSz6HcG+poDK4idb7Z1RM7oO5hpkxCaQRSt/H
JNV/NhdmBiZj9xf761NiiLabGxokNteuSP3OSvc1XpivCAKYBiD+NfvAZoDWEbFK
IJPc7J3wiKKeSMctPT9wyLrHCuVmD6FJP4OkJ+F1YcLVtYlNZPHTpiKJOCKAChWR
yAGs4yIyR4/kzpx6g9JN1lrFAH4kbogQSIuozt7lV8m9MxCRxHS63rjoExt+7b3x
ebVWwPe6u2+9IWLL7DIKENYdfnqsuD0T6d3Q2yGV9a6ssl7iKDrLdQ7YwzsDN2f+
E9MjU3Q6zJ4tnYNFSSwmIgtHvcbzYoepOntXM5IYVDtvq9QdxqNNBrovEWNKj/2q
XVAj4wEzEoml4bAhecy6qnVBFvgs6nDQEK3xRBYTvifMjBrnufnxYVCIm8RmTR3R
z8LSLFvOuD0XCSK1Y0K2Kb+BEBwzeIECD43dqLZDJ3a1w9bdXsz3g/0SPrN9VEiA
2aC9GCbO2RwvFbSyO2ynPh/YizgPFY7tNjA47E0FUeA2MaE5NYhszrGBm5iSwz3R
rkAXuH+trA5bJf918lUldbctjl5UqIip5IGFO393cjvX2Vd2ymc06KoOrfUJbUSS
qDZUvMUQeokLdWo2f3B6az2F1v1i0Pr0UlplxwtvEhux1UzuCD6BMrYaD0EcD0yw
xSKKLcL0YM10YBayfKCZCTGmR6EH1qujx5IzfIBOVKjgrZBlGxZrnLALauhe8nWD
c37dO2FUSgwJ6PuUofuvXzYRPFXx/NMJ3avaIO+jt7pDj6NTe7J3Temq06vGh/uZ
+wDjxKle/IdBgS8BgJ9hCdwOg5AprrIS3GtfdWv/6wLu8hv52Q76m8WG2ZNOvAWu
N7Ernl+Q4ynfClT3Quq6xNLcq3c4jPVN388B/jGl3AJjWTWumGAgZCrxK2fIibo3
9IW3+WClbyBO69/qvI/HlSATNsYRqPmNCAQKGhzrbZYmH5wERxFyW5YgVGWvw4JK
Z2mtHYOEfi5Mqm6N0GQpI5eZ4BP+C5e0dj8inQ/pc7DWBQrfMu/Q452oaIaLkrWC
hPHYos10A4NTXAun/CRNzCBOHLDtkE0jXx1XLclIbLQXE3gN/29T7Mz1pCGPqaVk
0wrdgjwoeh536boCWbFehrV1LbTzbsye9W4WIoSVa/XTTRbtlZwYK2j/RhS79vUt
1v3lyDNobX61KNTpfS/HjUIByfsOqL6+txP5XghlMsv4f8ju6G5+PIC2+mKvXjnz
3f8z7XlIb/IBTQuXgRpbl2fnxCKXgbSaHpphLOlxTYJTmGOp991CU2Ls6x7o/doN
`pragma protect end_protected
