// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:09 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ab9WRRDH5H4oO7Kh3r2PMGc6zwDyNDQW89wIXAeBU0bcZOiQx1MXwfnWjLT33jFf
nhVEDUWo8Yj8HIfFI8RAoZWX2uFhg243We/0olVpzLCVAKxMnF5SErF6r8wOocA5
cXO0MWwgRBG4Wfn12aOVQ3NqhUVca8I9mOQqSOW7sWA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8896)
eE+dYbXk7orXQDCDDuiVk1J9J5M647EW83VXcEkBF49QUkATF0DJduqUCXgnxfh1
5/fcDGQoTIKC6+YspOeBUVegZOhX+VMUfMhkKOypF3qcaKUjSzHiWbSesiFIRO9c
qCzYGX6HtRv8o16AjK+eVtj25lBcapkEj1cO20fzcZpJmTEEcagTXqzWRYtuOlxW
MwhNor7O1JjB2GLY3uBs/DOGsxjOAJ0B6wX/+bjeBfgYfpy5IjtiK6IaA/IZPAL1
27RsQ0M9RWN4yqa03A34cY442wT6XQI5rMaHGeR67GWfYUzkreu4DnHKJ3Ok8EOs
pDx/KnAy/hIaF2Ny9y+GIFMLgVRV2Qb0UUMNP/JGJ8dOe61MfePp0qJALXOJltIC
Os7mF/fC3WnD8s2mq2RNbg2fJ66g84qm4F6SqHa4aIPsPIIn4HxqFosv+1assS+j
RUFM8HUPR6sEPAtMfHiXcxhCpHCfXY5fMMwdk6pI9XBle6ykUG79Si1HCMLR/ZE/
67AunmjEnHFaMNgkN3FJMDo0DKMOqXKNLrKut55VWd9iuU/146RwjbCvFt3mnXN3
rfWBAXSeGH1h7avKAZ3g4I3GWNeJvMPMqtZpBk835di3Y4vkt6TeRcWnX/cakgsB
1Z7F7l27wAQknbnLQRX8RfJDIgPCP0VnfvyReXT8xiCw+K2ffJL2NdL8FYeuGkt6
Y3AEKQss90/aqBEqS0hhoMdHb8uOSi2lAIc/2EjV9+YlMfLjeC3J7Khh1zXAOh2D
j9ZzTXXIG0P1RNrkNFHVNo9m7mOcaFqvG13OGfcyEMxVdM39M7ChQBXfhTtfe2tf
SpdeG5/l66xKIONsI0f+7f7ih836waCArTCv6cwgAwqnqVWTpngQaSY85hwm025E
PYKrxLPJ9kwaZEJ6AqwWYpO5sFCEXkqAvv786qr97l0kKWPcIrwFQhid5qKa2Clp
kw+0Uh+9PA7852neDvQeTZVl6+hgt8QZgHqY1ibAyQxd7ySeK8zB4cFek6vCp3fw
m1rYMU/lHsp+5CSY+42ZUtBNxT2POeMOpro7AlrH9B+TJ232runCGmTFY2GmHrg4
G03haDI1cUbF3h5Q0Z+HYilyjHvyza2wsCFtG7uBj7peZnlLbYkgDzulINiFmWKW
Wx8X3TCPtHgvgdVVvZRUbTM0f70V1R5Nv6IzlQl5CIPSc9KfwBL8vEEEb6mGinVs
I6u7qgWoQx3dteBuIhDyaSW7ueHXELt/RPPPGPS2ODzq1jLtwv2JCxDLvKiVCNMO
AMYo8F2Zb+lVHTUAhBQF3GHEhE1sHFYUxpXp5U2cOXJQdroqApWvq1G+LS3DTClQ
+riF8xg5oqEs4kBbXBa+RSOv+069oa3EvQp3gJ3GxG8a/utkjp5xtYtmCoE5dNd0
64UEPNrwg0W6UharYwpIfHOKlomkLm+pdu1k8BjQk41gFC/+Eh2zHPo9wq6BSK0a
zxHO3I/N+Fyjf60YdXMvrJ2pDgj2oXZLBToL4p4P6d0SUhdSh3aX1yC22ja8ZXd7
sN9sCXdE8zr6GTvZXoc4Lh6fRuQlMrXg0lbd4E04Jl26P277+YZi3cBkLuYQMWm5
Fm/SKA3y1MOk79if0mWIFtJq9cv3RH74ZbiE3uK5vBs/9HbOkN0xf6NVmagx72yn
w+aDluAc0iD3/BicILJGCZS/j82NSOfHHFprct4EHCnv8s4MU3cz8ee32UF/3A7V
wruBwnTWMnEACSFTJgubNpTZhOyvge/gIVuvWWQO6In3VX5weK/hwys28tXhGah4
hMknec/k+91/CCOPpgz7kanUvpw4pEv8UWcgoYp8D0dwZi1tltgsErP2sV/8zNmM
1WkrayF1OWrfHMFIvMZyZ0MWRs2Xu42kRlXb3/zXPeWFzowPWG+ETcStukUuRC84
K+VaW8dbjwrRIzGcvksYRbJosHgoEy4PWlaDq9b1LH84ZPea7u/dVmd/Z5fyPWGp
YiPItIUObfMwz0XgPgSzOUFzitXxqTXyamHQ/i3ZCX7UY33W4mDznjiJuD3YJIuh
US+apea+PZ2GG9O56z1jb9FMY5LdMr40G18dZMb9rvtAsfILf0SvwH/sA0CBATFM
njJAzOoTSeexwIUk2AJgAeATHrT30fCeR0Fb1A0F4TSBf86eeDPTY5tBf/y4sUOV
X4neTUOB3RdI6JUaoLQ0/UiNLEuC/ljvd7HvOfeZZyElQEZ4+GvPxI9DKjvYR1E/
Q0ozHe4aTYrF7pzyvKZj8Q2O+SczFh34pdK+0kyejEiiYlfzMKsTDIIbzum1eDvP
D4UL5Pw5QunP1RSTJELdmX7AwLPQjbgIccDc71TeurxMe968z7j4QdFAuB2S7q/+
yKv1pjpIY9VJeVTDa3gFFCBeAOcJWIrh4IHnKPqpy4w1sffAmjiBmrTYKOcwnAqZ
+lmOcWHikfIXmmgeTZQRIZYpX7yBxtAqDctyBObsnMDSFZMtqgizRk+82nXBkuSG
VzPrcQGd+QpB4JULiZ1NC7LdlJ7b5iYoKcbKcjKNk6sIlBi4rPk6fn+F88/DnvJ0
+MFp6F+XAl3qv8e2wPfXKFoj+dCT5Fm+N+onAUBN8QKU2MDn1RNO6Q4UfRyHBkFY
fKWIsqf6IA3gHPYYXmRdgRg8uVPEw15oFnU0yQ6yicQ1Z3nF4fnHG4CE1RonWukO
OBqHr/HjTwQEnNZB47F28+ib9GI+ixbEpAPbiqFHigiCTdpluRk/YKC1+S6xdQGD
ULt84NECtsny3ki6VUSGTtDQm9IbK8vMngRMC+dNHi5YYjIBZLgrPHLaVwWW0IB+
bXT2UdYdr8Uq41edW793VtYMsg3zKDhaNKT/gwUHH/iT2HDM+i37TJdXABx27yqh
6nj8b9BJdT2P3+Y9dDAUd8KjuSeuQZUnJj/um0H0uYtirpkFqfKRxLRe0IUk3sOO
4F48gL3QrPrguJ+bLPnKseheWz4E1doJtoTvbch7bqI4RQi/lxivTVGPhhwz8ywq
FaQiyzWXeTrWdLbP/2CzS7qWob2B3ZQT4Zzp+EaThgZiXb0jRdQUqB5EAW7Wne7y
zKKgbFCRDLx26BhAGR3kTMHSxD3br6eex2k5bI72/DueNYgyKcDx0DaJLmGVb4qx
bxSXfTY2RtzB0CRPoLVXTNJUoIGNbLkMoPe/dGIoDg6UIu4ehRPBgrVLrUjwlDGj
abafw74F7rQwaVc1Jr1mK1BJgLn/UjuE1QV7bQrDsRxxw5avD9S5XCVTOKrmfQv6
fnj5IuuiUWdcDC3CMFAJgMuZl+rIg1A3HmtyShshxMwKnhLSYYevF1YCuOEjqNXW
WAnhbYprpUsJgSwlIJ0WDz3ZArzhbkgRseAQphOe3TaDovHur2puLdfUNF9ToVYm
nU4Vqpojv2YrX4WDw+MZnJv+91wWSfu6ANiJmZ+V8smEoCenNSd1AZTuQW893YSM
8o1I44A9Rlrix6qSl/9hewZuuc7dzwLVTCAar/kFacC73cu4GIIju7em6FLfS4Al
0T/yQglmIwjpeKFyzka6kUqsGcAPTVC8toniJqhLZsBvRHCbz/5zCXAaCAOo9bqU
5uLwSTMn+hCGkrQtXessZnK+dfu7tLbPg1qyUVerrldIuoTBhGTTYZnQTnkmyFm1
YGsrpWDD21C/foUhItvaljN3ClX7p1c1kFXh1RhI0dATgJqERcByxAv53MhJvxSY
qS4VKp06jhNoNpKzGQsuqbdKScSNXwxhOymAyA4w99mial532dub8EgLMvp2qA3L
qZ5rsG2uDwy3Pz3rlQuHrvF7JGmgt+LoS4FlSTRrun48R3lzZKwkTcPh1IV0jAZ/
t/uZ7vYZnHHIhC9Ovp7gpgNpH08XALpNVBSmuY6x0xXRg3UilLJ+X1WBb1XUX++U
17xJIQWiF0XUJ2uD0m3kgovpph8LY+ZHobcl8EnQC9QYA/jQKnwVT+FH51lg0A7S
wxGhPACf+s2qBrnz/igUaH6DCJ/5itepP578orkO7WFiy1rCsxqUuzwV5LolbxnB
exabKg7qtjtDeAJIZZ5Hgu/hUdHVj5Boy+A5BRVSa/eMxKCtz6WnX2jdY1J2paCX
VZLu3wx86/J+NVMsBoWR1qAqDj4ikCkYHVLwLuxRowlmr+fFZVBUs5n17lIuArBw
W4sj0sQJp2zw24HwYPSkk3whtzRzNnZdkQP144MF3UW3SyUfNoCQPea2JX9QtPCn
zhp3cyDr+l9IeMkWx3yalyYq83N3UOcZyfbXxOi5kLw4g2bA7QTiYee0W+3sxb7g
dXzBN9HLOEk+y2BiVcLh9W/47RtdGvKtXUQY0y3yPAC6TEpoLEBmqqtRbNi9fgll
PdxlBM8RNS5mOKMH/5IXXJiZg2wPf+Ta4KH2ijURESDKUeyjbIvs+9ROLjLoJlnX
0sl6UGeUR1DhRA0wlFlm9UsWegDo+Wb5ZDxT5CIchpq14BsKjUQ1D09l9WSjZ0rS
+HVldZGAUPtfmZQtUxPiiKqpg+y+L8/cYu7/iiJipUgTUAHQ7od5q13pCsMQor9p
FCJOU5VurWeR2o3LryNiTwhwwjCYY+J5G+cKz6RA8uMaZWJ77YZj0AHsT7+kghA3
7VQCtRGTtVgnKvcVTaZ3mx4cyAwV7gqypa2paakR1WKtp5e1sum4UwXajSQph6C6
+oclxrZbucTSU7q4zJNDcCFtvv8DDeYOqgIfTXf6dxbalbf9d/6hNNJdO3p+pLRp
BYo1gOFZebOAswnJjjeOKQWj2ZAKQzwFPUhhnEr5lpFnRlQXGqx/5Sqmi88fXRC5
u1bmRox0JnLToI8nE0Wkuv2K8rqmTs6zfXxdnX7eVjQDEqcTW58WWIFGSe8WxTwp
qda4UIUrf1ZM0nPckYx15M/z4BMAGveNNyjAI/ONI0o9ikbQlZp6cPzYYO+AOwJW
fCaqJL/2RChH9bFUMCRxWITn1VbNsH32xnkNiI8sawqPG4XPH/WTJxsMZZ0v7BF7
JRaF7+bZXuYZpGvn+Scd3/OkzJ52eif+xNgaoZcH3p++a9PiiyRs7DlcrPVe8txZ
PYEcBJu2Xuin1KD0PwsGbvHZQg93d0soKAqgtQ+Fylz3kNZnrqo8DgiQ8Y05vLZw
iN37YnUDZP8M9Axn5An3g3M8LqaZkeU71Kar9FlqxXXHoGwICJ6bapHNdPJBM8pN
pFR1rU+W9nYX5sz5etcgTeT6cqchdNT/kzsAgtBJGvvq6d7K8Gqzw9dPO/P07n5a
7204n6PFjDouYKJuctVkHzjLeZuCKTwTD+WRbO8aZmiaMlFM6MfTWLyIZ5abtpku
y5f0gOFqaB7jCWxRj3ok1RK7yjx8p9yfK0KF3PKRh0AGdf9DHLNuJlItbhDOK0MQ
kyr9AImYz82bxhv9j1Tr1Ag9Iw/OJv1Nvv5dsY1Uhkq/u1zDmZk+ASqkROY6dBUK
kxUnoGrNssIztEcglblokh+wsccP/tP52ac0gToUG+3pOHz8biy1s5Tne6yqBcUi
HEyUF76V7VPuHt3wyUJCcK6fZAvuwUumCv2Al8VWsYI0Irf7MTjyzo3L2g2Z76Hi
THDYTz+1NbOmkz5zL7YEp0uuDYkzNygaHiAIxcFgJMK/xYJyJN7YtG1rAGcrJI9V
Idx61VULqIRO5UVWmHTVognEiOVeMSn+59K2LmvSo6GpCI0wCx9GoFT4vj/3RgIU
0m6mHBtf6aahV9anOTGcLRSDZp7JWrglhzIcfUYXohdbLBQar7zyxi8DIIPSCGMi
AxVNvdTsOLmqlxJSKJxgSO5ijQBy3wI0KoHzXa9Y7OZ9LLdna3Qee4KW/FYr5T3T
AxtwMjDoZZ4tFEzr759HrKdOwlG7+ym8gmtM9rhZfXsb53RsWGXGTJZr1tpxEASr
DQ8GriiWD4X9XeO01xZwULFuFGqsKGhxpLBvvj4nqWv9jEyfADVgQLKw304nko8r
GmK9hANVzanaj0/XYvYyb6kShr2Q7grE5Om3MyHfbDWN0/ezd19enwZlVWTINKy9
c0IGK/WSdJ9hi5VC7WjbEdP28WoyVo2GPEySFhJVkuyfDkvRqsuXAH7pwhQj8YGl
U+8uvGNR9cyTfzoNdOjoFEp1Jk4SFjKXcPSl7EyM1XvVYjbid2gEfuF7+YdDCG+6
lWFvkSyGaVsDrEKST853Ms3pCzMFgyemUFTKnfJk966WIwug+jnYPMQD5X2uoPry
7+uy+ZRGzbz37O92L1C98//WoP2Irch6J6BLACeHDH7h5fkUlvKer+4tSQP9I7Tu
6/aQgaJouwiiS07xamR1/5/LxpTO5MKgBXQXS+XehJ1p81NmC2VenZJB4LmyMxRd
LpE2DkqQ99l/IzvEtRBL9sr97+4ZgITl0ucoLNIR6SXUTd/DITg4j6THK1ACJq2i
570eiCgiaiRA5UJ3Hig9Dc7iW7AK5XFI4K8qHu0t42EAXiJGQIwVwMdEo3IjK8DX
uiatzW7MMovtHMKwJGhTT6RNUtUQ1nftNBoVzVbJl0874rULN5TOvp5b47R/hRuv
2TFBoVTDb83zEM5RIHsakpKoThSSO3fzZ0cYKcI0MjKIraSuHiCz/AFQJ5aW3XeO
JXoGMabusWw//0EVaTmWzCrxwc7OfwQoWqoXfZZmVrXDgpyPE+W6f7s77n7thuUs
AS8753NG91XHw3DCkkoSlLRk/LEskbTrbGiXaxUrXWgQkW9wh7ETZN/wkP7fd1ii
kNb80CENlcRgmL8cjDotYamGKXXleuZ/+DtMrxanJ0fp0zB2zhvKiqGoXjYORnPy
B0HrFP3kzwgV0T73ixLuzh4Yh8VwfvYqDs5LrALSJw5b2O9ZC/QDygxUFhN+qeGB
YT9lPM+6lgJXzJz3H91hGst+PjRqXKPZinEBZglCoGzRsjU42Kpg8cFf7iTR7J5y
LKM32SdHWtHE8YRU2xrTa5yVs7xDKPVFb/5NHkbgTeLl8ntPeJ7/XnbRnPvPTWQ7
aDhNj3Ei2Rl74jS4EtCCQ19W5aAlTRB2ZZtQTl64+mVCe1x9SYiZaR7Vn9ZUQ4tn
gCls2mlf2CV5TysABTVpaM+AXsMmJUkszghpF5amKVfv1qJ3DHXQRL5nMcum+kPL
baHGAzdcajwB4Z0fl7JhU2a+P66WToRmEzXsyhCpt1Bpb74zToNfopwwH7mbVVdQ
Edpt73CoOjWySlWlHqdclixE0OqLdervbKksky3SJfbeBnlrTJtxWVYx3ZmWhnID
bHN33LHzv4qlyEZYC/c94EzkJEU1b7h7UZ2DvNOQCzL8zPYU8R/OHezRtXiMDOQ+
SJluV+aZ+ij0YiJ75SQG+igxJFwaUORHoB/ZBrhkiNJv61XuilJJuaYdnSP8u/lq
93tnRy70kEy0jGo6SQdAi64jv7bbpoPQr12opBidHso5Sq0AWhT26M8+iRaSfrPP
7PfUdwvsu/epM7fXZAD6dZO9F6whJWSNpYpqLYCcScExwUHL+SqryUdNtAmusoUG
AVpj3GqEIhIiqYpUEQSYo0A+GqoCR046hQyaRlhFilDP4AL4c4FCAoGHEVZHM9Od
7bRqeSUtDmhIGrIl+o0aVYTjUUYrcEDoOAFhs/KSYexFsgpV0FWdNbwixoR1mJWE
n8Eqm+QupkeRxmsWmGR43cis4iAX7PlrZAPkRKy6VahH7H7/djOxsFIK7k+79IiP
aiTWB0s3ms1jm62h/174q7shh8RH2vguS3gP7OeUbDDt5Hw8/+UDCqDmtgnkngc+
YZurtn2GZBMrZ9yqLwnauP3biHlBuTShdTxNdAYgsGnS3Ywv3QSSHJFXQnBKBsCV
7D0i91KGxNOdIWyFNLL8dWS3jityFxxJpaL26vkznaomgAwTR/MhkrUCa9GR9AHw
EqQAWZbsmH6H13Oq0Nb/prtB7KSx2X0GneDNSK4N5y3chTtgakinQ9fxThoIA0b0
k2aKjMTLnuJQ0XZNXjKsYX/V5RNl908fDpkAdf3sh6ILDEdYyZ48NghcPMnI1IGx
WSXRHTbojl28C/TYFGrPhTcSHgk4HFoykgVrp8JjtQj0cxWBQ7JZtiMk8Zc/czs8
wRJ1PkB2/Z1iwHESOzHHytbYFbHlbujU/oZxXyX40NvnfLPw38hgPwqFaAQJfvOe
4fSNCzAHZiznBh/OnlQHQigyXG8qt1/0GosLf0+L8vwPQHJHX5fNu2Zblfwc8ngd
6R8PGqMZTXgyFAxQLfKT1sZa2gvpChMq8kYYMkhpEovWooWPV24WJuC6d+6G1Y4C
rwOKOJg+WyuQrA763LmKKsI3eOokvX2Cq/AbLPztsseOon9sR9MEvzeyADUldC8m
gw8TJwkxmZvU9krAHk6YQXnLkDYtniSAxo/AZfvT2vmW9veijOBxBLdsIWNjENYV
/TWSr2EzYDnCc9XEmGnkk/+EWkglkFsQl5r1QkSxieS0qZxD78c23uin4R+B1cnk
qBq24ybi+zAmTwH2Xs1+KHTSbvNFbVIXAxt/4wldk3PJh3XPU1HD2dddRuTxxI0f
tMiHssaWmt/orZKT4aYIrgwUGWTbyGrZ+1L2Jr6Y92wjt7gbhaYkfYihlrrvArJW
ETRGDOJG9OgIREKkRnhQgXm8YxtoyO4UnU/fJ3K0S3pFZfYZraeV/LxV4OCWbRB6
P8/9zH+p0ZhsL541+vtzDXTWnjx6Iry/a9J/EaMzdaDWvtwCZJNs+T/TRHNT6WTW
C1wenNPa+SB+p7E/5vfG979gaUUGbkW9+N0XHitPEXvntwOJ1I8JNB1iG55HjuBb
5VuBZkL5M7GiRgBQmIqvjDd/sqif6KTmM8ARoLpkkvBkASZE6ch3DzPeDIru3Vrz
IKrCcwJnVMl+V25+dHGt+Ynmfsn/B0WcmGFhjYY9kAUE7dP5kJSpjvxUBsnNw2Jq
kIgnH+Rv53JCnpfcmChQ8u3qHiirc8CksbemopEy6ZcHOiI8wWQFckkBspUKfUzj
tpaUZn31EQPLcWT6KcZRw6Q033XCjNRlAd4Ksbk6sphsu3X7Pmj0HQ3nJC0fp4i/
BB7Nu2vddhXUHu2VTbmxPXBW8VgxwTpCrxGzt1256S/tu6VorsNWAGegcfhcD3Sz
UuucsEdK4ypjPwLM50xZQEcLsotURONCUAO15B+opRNbIaS/7F0nLHmRnr8ExFSA
nkvROnMj1Zs0DOnYJ80OTAG0rFg3ibN1SIxI2XS/+XgR259iFTlqdB0Hjs3GBLE0
yMEy0tW28dZtE6xvQN7YipAd8OhCW0v337nLlGVBmmz6ZFxHahkLTDP2jBEf+16t
JP7A6h44h+BZyjreqLMh6KKnYw/M0jWfpRzoWil/UYukmpAPfWpP4v8S/a/34sAe
BTzTUR+CNdE8Cu/kyDzIY8Rjh2uC4D+GtWKjFqAkwSG4rB7k6vub3PdQm9sX6ULf
MXFuAsBnauDcH69Bsktw3/54ECHdGvPQoJIXZiiVV1Av1jyRW1p7loKEDuLogMxI
5IDR9L/xY07lQYhu+6LXEHuDtvi30sLqs5yeK9onThy/22C83e5ggDhdydJCeoWa
QTzSHvuA3QOydLNZDEv5fUFBMuVzlFma0mt2kZn6wvKtL2x835JJY0V47cBHxTl8
E/CQqGpfi0V5W+PMJfLhN9RfVfNXBtODMDf6jR/Df9iAX5QI9JkFQM5V5kuPsE1N
xZybLvCqsVyV9goNqr4sLB4Y1rQ89VEVGegMMj9zeDMDCgXcNF5pmpkWWmHR+gGO
dTofrLXbmnz+3gZMLBW+w0k947tT/lXZwX/1zkzTsAz+kEDR4P+8vn0UVaxCfLYd
Ph3nNvz6u8Lu3u/tI2n28r4uvZswjIdQEFHZGyBK9uOILJP6wA5jpLz9qqWzelff
xP48v4rCeqR7Ul/r9ThZF/piUKGfo7L4PW/H+uRMyE3POsWUxdfbUAWC2hVLUoOU
MUaT0UhKrorpNWxkxbmDaXrV7xUIwLx7ymAq74IW38rVZj0rca6uKUHTWtHLWgt4
GIm8M944/Fh89p+/dV/8UZ2lGkhWqTC02nXzBx7j5HNFt5zvPhtfwt9wM6aDxgYo
RA2Lt1YLh94sqNQ4FD6kOxWyXYN5xCd1ejkh9lYgsZv40uDimDzOxljMnutBYpMf
sO5wKaC+gMg35RHV6/8Cotsv+WdsG10lOKpsqpdXkpd7AOsLsWd6lN0ktNSAZdLa
yujbrQq3EibLEbaiWc3itlzTkSe75pIALlSY9c19L2nWKPfdjo/cdHHqKpMaUmIS
eA6fFQb186Q6Zv1yAzyzMjwfj92BHOy3lCAnZaESvTQyuzNcUvXBjTSoQYoOC0KT
93xfBbb6RoeKTjU62OChfbxN81vI1fnlAXPHlsomtkXAMhuBqYfwe9UEn8IkJWyc
EoJcWml16dVbwObcJkxtgpV+vrCgY8IYLxf1KWYXaZJ1243nHBhER/uQy33jShWL
n2D4U/UyhNYhpsnm6Yv55AiUf0SgT2P3dohlYG3JrzNxqMcNqjb/DtVh2lPhtlWO
m/+rtKYEUkU8mHBPPnGOcIGkJHiDWIL+/vSQRymsf329jHFnhALwBDQB5Rxwnv6X
Q+IkdHUQmChvs2fgk/QonJrFN+204NiQXYUiIjdS+GfS7weL5PwcNGvcj7rTmtme
ovYFbvKbIeeSl5vdOqKJ0QjBc9y79TdeGHeqT/N8G/HCwUlL+NhVemNT0dNrguzW
ErfbVT818sLNG+rkybQBP8yJltVhW+MfwBre/Nc3SATFhCfqga8oONeAvyZd2yRJ
SJNF2qegIZhLHTU0BhzXZrtexc6Iw2HDBt1Bn4ZqMXM5CrIrdQ1wo9ic8ooBWpKX
kn3J7aj6GkznreBvbahbXxUkhLFvQXQk5PgFcnZVSuFK81YxDPMm7E4og05nmlAP
7fYCumL96kz6WrEPntqxXUQ7RM6wtTrUwXtIGXfMATt+WFwhXRJps05v+xsf/sSF
wYxlvt5fbPxM4Y0g3ny0k5L22zhnVc4fUzcYwBCEJat2U7m8dr1zJdKUX/TEvYnl
zH3zY5UaI8hpm6EqyDmcVt+QCUpPtmYBLr3W7X0FSBIRbT45rypucsHYSGgTCBPW
UFRYxxgteOP1jeaX8wjxIq/8gELLI3mxpk1gAdue4rFvezMBfsTqFi2te+2k7yKY
qeG4iKqH+4oF1Q4nVlvDZn1H+dORY+CWEjuht/UbGvRKm1DSApsHA2DBnj4DK3/+
zRe8xnO0VNpXU32X2aMeNlyef0w+Hu5oRcHk51ZAo9sk3XBvxchrYCn2/ZPVydOS
6mK6+snXAFg9d1sQM243Z8jaMhRacPUtF+srz4pzVicz5qo9rcFWcs5xz4dSqnCs
kGls1bG5jhINdyS5ZcgOhNQQxpqgb/ob/N+fS1ZXAF3/0quYy3cwjakWuR1pIxqY
s8sSooP9RHIQ6+CS6elKE6TvifiSb73GiD6NkAO5WpZEmHQknrgzpeKz5qG5gJqv
sL3icXf/7RSm6QmH/YzpU+oFFnNZDwaOqIxX5sNf/uXpcchdPwX6LndwAhXb+OVD
aizzTj9sqQ2wAJLUNcE0KyuFSmWoKJnWq62De4LQFgvEpqtCZqUQzkQxGaanSEcP
8/zgauNsbvHfcuK/nTX6h30t7E4iEEZrY1vuhvvHlabQO8CUvEFDPKoSpMdZ+gvV
hIxtDAcXao7WDeIi5HjNKk4PIkry8G0rkfKkkKwrIO87AX4k629PkSJIZC9bqUHf
VKJD8wR4FE8r8IZCjTcJTa5YpyRzpHfzRpwDiMWyYx1ALP1c3J2jJv19qvGUjol2
8g3xdRB5ePivoJNaBHOyE4v3E1BHaIPzl0pElNg+i1HzOrukVENFsCRowD6zxI09
WdNKdrH8el2b7TOfsB8Cog==
`pragma protect end_protected
