// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mOLa6DlmzUdzTBBZ2hzu939TuU5FbLM6EaVIJBV9atW4U2tRdTCNttF0NnV8C9CN
94HuvsgCWYdU8PzVqknikb9SDsAhVvxCdGe0XdFYotpFxu+Egyy6JC4fY/PC/RRy
1fNwegbeHWyJfIQd2KVBzBSWbrvjkFU4j7a995RTLLI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6048)
KQFnW4zOH2mg7txz4KHIUCiJ3knqHS3qswAunI4eslP1kMqSsdDVDEGTnYCpSN+q
ffDxQYFYLoWtmWwR/SG1UoFkoZ/To/SEOsJIVRsqvNhq1rqSpT9qVkH84Mwb+WTw
bbuauR0poIBp7FHqWRxk/XPrG0sB/qj37G2UcIn48/KOBCHWfY+pLDwuCI2+pnvP
btjYf/jYF0hM5UcKAvsVJcF6DfG9kLbmQx69nSXhNOqatoPpccNfzI4jFOHrDOV5
bMZ3DEXAhnmu6NLpRG/zIFVGscPPASJghANDZQQxnNUC1bPoi7SRjj0eDyw3bTEr
mc7d6Mg2GDzv5+RUefDcywNNW/UugEUzIPu+v07P7N9uBt1KxACQ6oeJ/kE7/h6W
C1ofXZMO7WGx42MektbHM5ToKcxiFNSVp0nr0Fyc2+ctBLUGT8v82lZw+b879K/7
FAkNOguozvK94xzWiYy849E2NLTLYNV6wV/2LnmPRYIeQsJ8EHDxnVhJqjSaKEM/
P7WqHY4TkbFJTXsnb/Bwri2COHBev5c3RKK7hZ+KhZF9FW/DQNUdjF4SPCqGSDYZ
ifaqSTflZnC/HKFh1wtAN5pAh99RMZwzRdS+3VT24ug72D39GarpUEI9FlHVqBUe
8fguYewgOTV2DGcFfsRibeHGX8aYljeelFagztb0FDl7ZMTAUG4jBN/Jj2EWfxe3
GHgiotzDqXofVlmZyuTOhntiiwl2TO1A0ctf9/0S6Ppv9RS/ZghL192DlMl2bTzP
QMHkfWx++wWc216arskyTD2JVoebDnlOvgSQopVVKoIRAO157iIUhnw7fZVxSTdn
D2svhUCRAsYOR7cWnfSny/zZekkTYI9qdreEwwKZ05wKp9WkaAJrSdT1S9GpTQgC
/Elg5Kk7/IvZJ7JeE8aPTYL/X1s6GDu4IwpQOkzTfmIEh10F3BkQTcHhMtLkbw90
HFpv2Bw7dheMwkyvsMmaPxC7uCOTXTLRQJmB8918rAi65ZQc1o83JDiN+5XAYvQs
SqzXjrTuMYnHS4ZFLfCOlma/8q8Z/QiEWkQiT+6ICGSwL/GGclPD8lK9EtQOSRnd
UBefKujj6OSDX+ySeLrC4tURvPI9E21+tmBKu7hh/bthJiD7hjE2y12Ir8xcxBPd
D7eIR1afLBwcaEXSExw1ILJsaIjMJmgi1GS6dMLjl8G6Dx/gtT8nzvjPhqGk+KSS
pwqceC/XWR1MuC1xggrjlKHiTUC30RNjCFtlh+HpvFzuQyQGaZF86kEOO+MRWE+m
CqHKWtrrJrQt1cZFsd3gPfXCRtpE/VoinmNtfSnXJhEAVNqpGQLzg7UnwageUArD
H27GwRNOYiYMcfF/AwDjveWgsyVX+dh9cKWDIYFy3fnWvb9lvddqa7l577IrEbc/
3XH0fIj8SRXKm1wm9h5JNni6zMGQ2r60H1Uxp0Fx52NYdfgcgGdSguMVDTzyn0Yn
eGqStwBStuIzFB0m7maE6xwuAenYnJi/vVHr3QlYzS16eAiOvtedN9zcL9JR6MrB
xMPVTxN1+Wm5Xg2Twh30J237IcCDQKGANYgJmLGqGYMKDN2jEly3Y9jsT41IxQJ3
dqTBJK1oK7BkwVXY3M/MCfmmuqUqcf27wQ2n79oGq3fUPgQ7G9jKdkeh/gqlDoM8
kZ6mgVwtbYLa5/gew7SGD6CJUHuoVwXKvZHHm4HVhhXpowYkGRUxcvZe+cTolmO4
1EDRb2wqQnj55qDyMbaAcyYrWdWAd99tMGd5+PshzVi14Bj2KilkJdUmODR9vIyC
7LJ1sRTy5J+vg1U7S4Hic9rExLCycUXU0Of5S89AQ8pWJidgA5UWhe8BlTPLKCun
Cg4OQsfUzdukf8NBAthHex6J7xb/SHQ4OJqlM1Jn22Dxf/tIrDhqNOimC3Gf3jDu
QmpLtLgrA69VYEIhmMmtFKyi7nHTZV0mu7f6dOxfTUfL8qQzpSPtttYO4h8epYcZ
F40IcqSQod6UQNVTf0dBdndFclPzgiY99dq/IzMU5I/7EhL+pclw5pkF/6P+dXjt
t4KxghoBbkEVLCYREkaSvH5ui7qTQMG+8Y5jS9oukBihVPmMsSlrl58EystIoctu
5Vr45c0iE5a1H7E4SZ02O3AGtbx92cC7yjOg1ayb9iLVkwtAIjelrjCdUOi/anUC
Gwj6RXWDsoak0lKbpiLlznD8xnWaVzR44dNDtBI6G73jybaASwnwTCAErW9AUktf
M+wxstFsPdsmyjEAFcC45ojnay8FJ8tQUZFUZPCaGP2d1/6MX2A2tOJHgIdZDaHC
7z3aXrLtrqYJNSI1OCYNgjrIIGdSrCyODXQ918Ull9kkn3sskaqCaoFJLkLUZod+
64dwC0IgUeF/zE4FFAtyT3eXaI493z2vKsOYUbHgqKG6U0EwVg539NpY87makcfl
st0GR7wwuM2n2+Y97JlraSf69/2tVlJKxkimvYV1SG4k+CG4Hehq4tbHrC2WrZf8
Xb4zJN79gyn4BYzY5qQgXmRILQfrInQc0jkB0Td4rgr/BJJ6Z6asJTC6n7c8Ji1e
fOMZnIx2xPJrUSt8dANM2J8QfhDJwkzt+b950HEgc4nJ7xyJcEMmHkYyaHxpCm8S
9GPL6CzG6jz/kt3zOcDVt7eIrMatnlRBCfUQ44SdR44lfOWtAdZBmMo0SGmNmlo4
bEFKESDXJf10+DM3PpoiWP34iypWPlYGWIom6F2j92wGqvNhoA4MJKYh1JoIAVtW
Ztb8usWBhtPqYj6x0Eyk6tHDtBHDNe4c4Ke+FOpFhevvzsLKDK10aROvAXE6ntrl
rH4arjV8Q8FkxukK1w+5hU6Rxlr7DmDFWL4N5UaGhymDWTCOhx/yQ/GBEz44v9Mw
e8VU0/Qn8Ipnp8S361v3EkiFvExBn6NGawHM1zeW2eUmkbeBf3aEMmIM09nbelWh
YBnafJrOoR68Ha2Zdg7BaN93isjJDGIvcWR0iazMGJTBOfyEI8eyJB3j+AS23Sfj
sZTm1gylJRbO7eo3DDpzoqy4QwZsEhR5Se8EVl7HG6gLfiWMdQcI58PSsNiaS2Py
ESFYpuTXFduEkWuBNd/Qz65ZoXUFXcQ5q5iI9XbSvpCNt/mVrCx3nicDnBm7w3jJ
wbaCYCgsJ2FVD/XnBMLHP4n5JnI6wpQ0euDt3TBtjjaHHuTmCyT9BspqHxsAzuRf
GFT55ONwN344JonWKSv5e6Yrcd3+Ry1cZY5OGoY5DSAJ+pCWxigRVFD5d1CA39MI
5u2dQAxspYHG2DphqPevOYi+9Oj8Goj0tYJlCutVaba+JsVQI1axJqYo30RFHInt
rUhAWfhaos9oVnqOMWuVfVEPGQy0ykvp/bmr3Xl9J3QrFPJmQfl9maVBZiG3Jo5y
vVT3LyS+sJvz5pgE3pr8P8SwIomwprEraM5zTGWacCs8makuscrVUa2IHhPQNN+Z
QK6JPyPoK9wQq2C76SFI43FdnKaeHaWamM8VBdGaGx3zvJyUUZe++WCHYPhISqHd
KmDysJ8Z4hqe855A06xOqgWT5foPJvh+HUfVN/zFYDi4RYiMFx3hgw/mMiPI/gMI
HbjJbK3/2Jg2PlEZQqUPzvgyZ/oTrVOjfj1aCbofiE1BrEOzijql6NZtXy1VIvUg
DQu8p2/1Rh2/AdXLCoMQnQUJEDu/GTHqznRJsp76X6TtCdHdlxN00SSSgzhvyG1+
IdU8JCFALEbDnKa5BoDtUJy582mjCEtxgLVrl3+FtOmRYKzwHDpJiQG7FxcGVNAP
XA3qxNVt9kQ6wtBPRdonIA0PhxTwGNPBx7qXOmoWT1wLOjpe5z5hotqKlpzFXll9
7Y617PUkCcD60eSGSiHcdxsTPZl+C76akEzp06T7LobAzX84ORcPdKO8YflM+Bxl
QRdDX0jtWv6P6AzyrR/JUOBxjTlCVk/JyvWBB4qLrhPoowO75WAXYndiTLNfThf0
rF+A4gdMYX7dHSrnDgzaYO/FLaNCNFQf/+50FzpM5L2VjhinnzrksKH5WBReMjIK
iLXZ6Jp752eY/Ahv5ULu2gzWC+v2a51t3xW1mmrpDs+CFH/J6fwA7sWIZvIFoM2A
D6NT5j0e90Yd1nm2udBSTc04sKzdHoX9PivbhIQ0VTZ33FSvaL1B+HNElQxGo2zc
d4RrS71RguSHBV8BonkunVsBVM4wYdQGKMd5ulLaeKxdjj1RqDEVwrzsVVkFVsyR
8cx4CJstdWHIr2YIMbaf/wZjLHk12mU8z1ZjJ1GOD31zOAP39ZuDRpJSaqM6h2mQ
dEPVMtArKlNzuSzx6YAjK/FH1P4VjEgkxS8lTmIbj29iZzooN1fwHnWztYkuZey5
ZX1fDCpfi090liBMlw4NdKQ8vBT2xfGEqSvRmHzI4dL/OXbJgkLnqVopzsL3uzqc
Ma3JPuCxXVOTx4Z1Dx8bTRoMnmCAOsoGibIZkGzpIJ4fJOvDgZGl13faXsTzrLE1
m8//WRzjXEwTHVq0rM1mEnp6DhS6+OGYKF8bgb+UzeYJRhg0/zN8X5qxm9Llho7i
x19oTdhACkeu1Q6rq2jPUv5NISEJQXwtSMtVIDdfsl6lm1e9gQsZA1AIxtcZtNQC
WjnXHZj6+vAncil044UJPtb08MJEgaCpnsyaNmyNpTyJPRMdftVTnfsxprSBUfUS
rDghlTIvE0TsnMfVgG+hdbLswbBREwuuKNduiVijthMjBbKp6LGqgo4N/FgPXfE7
shZLkVnv7OQHxKpTtlrRm0Ddf9KDBmdbI1LNiW27yIcs8jatZeGzQXk3jLq7/ZMG
gldKMjhGJSEP2nh16dNMAtC95u4MFJm5gB5xh/iSNMflTCP/8prz2ikeWtfBzCVy
Q8M2LVm91yLgMucL5W7mmq8WgVH49y0pC4aN7eUqkJ/TJwgsJtwZFcG6WIE5hYrQ
IXaO/Wb0QmtAzRQFLHfGbuVuy0Qyv0c8fZFW+EFZTHkpJzNm/PYY4jpdMw5oEtzw
usVfGGdiNH0Ej4B2HA0TppHzexLQQBYHBxARMSgic7JSLs1RiEgK5+npkSWG8xpe
6Tnst3ckJI6SaTFsGKWsbIjvzm/2NiHa6JhFWlxSqHw+1X058Dp4leL807PUvSCA
OVSv1qsgBhP3p2UZQpHq9nZwshLTEEnxxqq//wZDbdlIfKbZgQf04pnIcy6GdVgI
HlhADstC4iu6DZhlLpecl1CmBjLcjiyytSGOnLPyJmr8TYUPR1RHIwIPyVdm0oDf
oyfJD+sA3kyleUF4qp627nrbh2JTNzco6Ev6ONrML5PpvQJyUEpf1ULBLU10LUAZ
zluAtpfrjdjACoWYSd4qVdX6tvRwtsbl8L5z3FjoaDuA0a6dZxT6LOoVxHxohXjz
8wNnRA7D0SwPxqUU++ZXRCmKG4TUCaA0Ed/FL+Iy5uJXahhG2sTXrnfenoVOBdDb
wgmqWzSJ5DlmxQ4XUWVQpSrGGGI8UaaVCHM1wzUbTie2G5Ru+njKJQULowsAPCqZ
h0vm/ov8joQgp4orHLkZftizSbUORGGIlM6QvHlBiVGUZaYOj88bVb6pMDXKdVCE
ZbalLc54XJfDU9pEoVQW1V8WLGy+7Oc5lell3up/BhUe9FsE8g8m3GOkF0sdIIQ9
FJMyIemZin/kJ1A3oK2z0d2xVGtD4ceJ3LibLHwLqX2yYjX4oEWYKzjE3KNg5DA0
IHk9h4cYeFqlf1CaB1w1zruFmXbUTZvqoRNDWTf+nnrPZKCfegaCbJq3XyAURAG2
dkyHM4nJCpXvESAnRb74rNs1Fquma37xTfEkGE6BAl038wsNwMAxBptDIOHzVfyB
FzU0kHyUwXWpJ0r+qiDn0i5++T+PIoN6hnwLhYks2e5N9KKKhsjdQvTNBDV0OaLf
tz3I8+9k34aVsOilJBYr6GyZgPsgDEZGZvtlmcOkZ9P/inwhK2JBkAJTelahes17
HkYQIJ98Ze3suYdl3EVQ2JLcNchQPHEE/VDR4IZam0aK2qT3xj8UQ13wVrZFwiww
nvY2CQxX50QZ++/YBF9TiGjOadXVWpxjuUjSOKdVC3IKI3FewjZMbfeZvjPV/qRA
4id0RwhQ00GTAlpu8VNS6XZusCmIHlEzsiM0KpSH2AkOAVe9XQ/5L5r4U220ZKbe
dXLVFwb57nu/QRPjdqN/6ww2EhAf8oNYg6zRElYJh+7i1vzq1LYJOpSOhcNmaTD6
CQBgByo+dSnMd0kj2lzlWxdqGnNtxr3iY85wUZu7o5ihwBe2eulraxnjP5v0QuMV
+omAMbnxV1RcknxFVjFvqQSdLS4CtBrjI7REilwIR22Lw3CaDkewrd4ns017aTCc
XpSi2A3/am4q21BYD6wMl7cMEErI42Yv/S8DSkogPF38UZGl7eGmFBHlOeOuuhhW
8UbmPY2/zxGr4uEPyqMgbF7AXO14wly5zZ/A42jtB58Az0+ou5F0P0UCZCksUCUF
R6XeKZLf+c2fkiBTlhwwzgznS6FRxiR9fKTUiJT0/DhwsZ2oOJCtedcCavrUfG9w
X9tSkhcnQaINuRfTxdwuQVaoAj8gFhYKxdG7wWN+pUhXzm4l3uTXMu1belzt2QOl
ERrGx4mJzt0KeeRyIIRW3Mmusr5WpVKXtE5gjzfMvvREvwQCsZuuHOVNKABE83IJ
zXgnlfV7Fzd6TNJgd3mPsiYFnyFt6nlSpvwAEI3f/OZhRuBdXrDewn4iqUAM2g5Q
aii6YDc42JKycazR7Gw2CHKWRzXZ16ES6gaRl06JqcIT6qaQphsB3AeiCxqUGAHk
QkRu4H6kjiT6ZoHkiOKTnLN3zi/4tmHFqtTevp/AnQTXWkHrk2L/MZuPQGmWL1oh
qkrS2+0DPHwcWtxiFZB3n17ZdWP1IEspkL3XAILqRjd+gEQA9poVcezRd1NYnQAa
GSWOdgbGGYvZ3gfAnhc9BW33ya/ayAurebgtJQzEDurENpcmmqVuB0/MTfDQDJuZ
TEH2goz1WVD5uulr9imkV8d+sPrfrbqkqhqQwIaqksfF+5rOtIkZZtWfznhtRJMV
t4u9mVBMeei8Nj1IORT/if/lDrUy9ja10jvfk2tOXAmOUBB47ZhG30vzZJ64LqJ9
iF2zpIwVRIFkIO8tg/l2bHIS9V54yZgX29+H0ahbBqrpb1HP4800IXGjjfdc4U/F
5OgNzWBsldyYrXINI03/Ev5ZTGKtOrG+iwjK7eSv9vIbCQMLGrs/c6V/727jL4dw
P3JnE90HiS6MnJ2PhwohFR1uZd4q96PMaivnNxVY1dEwZqzYRNsyyIu1/slPJ/3v
wQNMIu2spYF9yvIYrStN0NZ4n03oOc/c63PJ05apwjOnOOPECpG9OKxTv8uz1pNz
2yJhtrWNy3qbu2GKFHNtlOZmePcgDhDSikiZ4zEOLN0BGHWwMy+iKTVHhyc9sQdV
X+MPAwx4rEfGnNLX9bjDFrag275Y5oq39OlePqz5TiFlKveEQNDnqZHKU4NhhUs7
F69JBVqHaKtO/hsSrssJoVqkeBjVIJU884R+QjSgUMkj9xntbmET51PFEpS1R6QF
CstPmqoYQeMbQQ09rqUR4SvGKHbhHN7fh1WzlkHM3MeKoiPjat6utgQQsVJLd6nN
0LNgDroP+/V1Cz+lK0oKxdSeytvPeKScaGqAP94i0V9qjX76gQYLGyPayyoYNxTM
uBnO3O3+YLsmn1RxY6PGiJGfR3wEr7Trn3ADiy64z140f66yyFIagNi+xaNGl74M
SxglpOctUCO9NVC3iLR5en9nFcBrbaEHOMtFshxo6oomvGDYR+goSVpFyKC9xGQD
lKKnPS5zqPwCoOKM6lDFFUlUZ6OYRL9sU5Mc7jzrkNHlcTqve6CNBseES5xFcLw/
8kB879bqXQNE9mfBrf3m+QW9bvzIKT4fCr5SkVT4GrFayTe2S+Sx1oAQV78iXFz1
BTBD03CyHo+fny3ZI7R3r/f7zc5D+L9Ivqqtj1IDuSRdzncBfjYAEAf8BxLywXUw
3AVrDhE+J2rdw6mmZllYAn1kb32vcLFRyxree8y/APNScjf8r4tfLkIIRb4TK9Ty
`pragma protect end_protected
