// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jq8Kl2348Idn8m/7kamOlSocAePqLqRFVvjy4MF37cUe6hi341BO5Rohzll9A22n
hNC256QrDiqfnORHehLPHht+SUEEHJUYxAzTlnr9xBbByhUNGUvT3+tL6Ac7vIt5
WPzsC6ld1evbQdXBf6cZJQQdRrVXjR5hZc6UKrlIN7M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3584)
8yt2scAv2vPIRuAaJsl1DYWRUkFRzLFXrxpmcVIhJvR587iilGTs5iinQ2eQME3G
ldwOHz/87DAMesxpXVDXVClFCM0KaQ9rG7KNSuM+WKNYMmvxBpo8vRFK/Va9zbvk
wp0sF/xYTcRhlOx/s5yq8aqbYZaAzscGq7ilDUjGw2GiNHwrc7pXqqnAcXLypn25
2MoNyKnDT0PgEzqYjkMmcE4ijbilsZleHDYT8U5bortIpCz0zBOtx5ITVJfeVk/6
o0enlnz3Tdow1ZlH5oRn9Czwr6TaQTysEWEKkJ62MNSWldCOwDfJh6ZDrZSQuzMD
I7zTlkbtf4uLUQPQOj/ujtvW70xU7m/+Em3uenPwOQ5kYPXdXD8ie9zjkB9aea6b
XX4fhCxcSGC+RwiCUiRmQb7Ja0oXD42pzyASgtZ33Y3PQxYZvt77ThgZfOYO96em
5MkqJ4VImCeFGgh0zI2aXFUFL9T1usFQfrd9bV6wD6Vc4DNiyPYL7GO7NZcNBFGx
NJ9CLQnB8fS9CHRhy+MO25WcoyqWMaKUiyYwcHTkgLx6sTEQRVvWcBOrxsRcCFQv
9Ro9Y9bpi6ITIF9BYz8hDMke8gx2J+ykuB1WzyNIgTzSLPqdggqKYvePV6wzIIO5
WXQrHVQ1WWuWwqFHIcrX2vbpNtdm7EJzt8bhpl+I7UanisGS9SY6KB9b4dq6ZMYb
m8yhQyU9F6VF9mdPpWqeU1RCRd31J5zoHrc3SFIEIh9oahiQA5AYwBw1H1mD2fm/
5Glgv9cGZ8hDphSfDSj6tGM4hNzfeuT+lHoSG+2vFTIQT+JcXWMneczMlk6HpipQ
2dk0Vz/AH6aZNPAuFYDG7bggUVVO3dhuCVz5n7wFFSPUAcDJKIJFO3JUgoNFLaPz
QVP2eBSbekgM8l/bR+5OhAD+QT6Y1+KhXwUYHd0xfJ8C7ANIWo+NZ33UcKgdHf4q
JKm9Kl5z+UdlJEWw9CqidSvQpCa9JusJ4Jpsq3p8LBcUEkTqJ06IEeGqfc2D9f88
wH1WFQhJXaT6fI0Rg6xdH9itBA+r03GQRI1JGEvz40ybjiE/HnDGqMtz6uswqXxt
KYYplrrri+ckrZbt5sAz+gLilkq8JpdugAuUzHhltK5Wo3TTHhAa06D53yNalWyQ
cDNf2Ed/P6sBho/fPKBAoZbTRdxAu5ZYcOJ3uu/H4Y80yS54OIV0HCOfMI2h4bso
MwIYivzZSKTtFxNwW0D9u3UV4tWxoPbDisA9sZCrPrP4DAEgvFPNMXILPMmOhcdW
Z+0vG4sdLkhPIwLIRQamoaennJm5D8DcS9WazXkIlc+U7wuo39Q5vCKy97ZAZ8Rg
cLvT0Szsixe2wPYGWlgLXmcMYltvpC482VTT/foTkrJYM4tLqF6N3wFjWk2oQOeA
Wm4RQM0uwnmT2IPex9cFUDpNXS3ot6HzzQWVw7THBhdS2x+iQN8UHYB3h8ySr/wR
/obEtE78Qfq1Nao9ZVc7YVU0J1wzabzETxFhXhz6nPjZUC81SPDHU9slA0qfLv/b
n6daUk3h0kTmt5JP5FEqMYjYYqn+sUK+TrGufpfS7dhvu/u/wBmzEMm5806Ub1i6
hmdjxMQFZvkho8HEjEFJ1bsB2mOrQzeJs85dhUWZvbAiVhGRJdLeghBBXvEJfiKa
T7gXPpqMs2oWjDz2owYvBjySQL+9mU9hXsGI/irTyLbJAHN+ss6di5wYhvbA3I+v
sFTEXTTMLbXk0M59EYE2cLNwi9nqhxCQksV4R4O/vTj0SlKG5KZPuoc032gvZD4M
euiNJL8qwvMHZYkmPUNcq/bfw7ybSTq1S9j22UT9T9Ly8rMB0JLWe7XSRyaknNFj
Ik5SFtJt/NZc4eZB0dQ2BibzBWOfawSdGc5aGRKjiMm+LXbjEIZQLt6+Mmko/otX
nbwFVMt88u6kW4o/lvv+QlirZ2vFx7qol3CiOBLZLY+HvEmOEAMDdH4osNRCCwBV
CmPJnoroEEEir5kROXUbaD+XGzkNPut1Gjg/MGCm9+CJkI0+ebutjXGMo4VyOf1l
McjjRe0NR86++BvhRtSy7NVI4+Jy7mQj5E6VnT04WJfVu5uieY9czwWkGpQAjoGh
JSa7APdhumxniWV+jhK3joBqBF7Un2sAdvOLD8owjG4jlNO4eJZNe+UtPtOqVbwo
VeMZNjQH3ydEOPwwHsIaW8v1YYzapWUldlN649gejHhxwEwVzE/Xqpn2lSp12HAH
0W9+ljY8EmKXzhfnEtCkrVJKJCQEctB+XYiuxgOl1qW4swPTGqeeHI5wjeZt2wKa
Lme93Ug+swjLQ7nKjjmCAZiwcegAqLsYBOPdEb66ZNHG70+ciuUZuCAhRJ8md88B
ka3MsCaU1i+c8vzeCll/OosdoqXceCnkx76v7lYk8UjGkDNNXiXZR4iiLSvzVj+M
BmORZeaRVdbzxywhcQPhc5pHiW8OzW5UvJvad5mpx23ZmBRlJbp/euTmTsIoOf7o
TOnnLql3aH8rtZIHeFYzLhXE9y5KGhJovoCbQx0i08bRezGFTse8rI2OzLY3ZBVO
vOLE+xVAbe7CJ0P9ch9tNQBaIcvbIRR06VShE9Z67lkn5+bGDj1YJ03+GbpchuOM
cml69flgA8sFga6LIV4mwm8pEy27eyOn7eBdjk5smzfgX3lwx1OjDF1AjOcwr8RA
O1AmpIK2+ihfp7eOQq1U24LhqauK3LNIJQcA7MruM86yrLtngE2IiLPG43YkoArO
fqs8HeaOXM5Q1hPntfkmq+rd6cqUNHTwouJPfFCkCSulDP/RjZe35GkWmtPp87kY
vDW6qyElL/7a6t5rhOZrzI1epb4XwB635ab+PjVm51O8S+nSZ53TM5qx4+6oAs8H
6aTago83wYLWvvU9+I5x4idIFO65LQ+I5NSggi1GPnP8F4OpOuzpI8yZF/wf8jfn
RFjk6JMlV3Q6NhADUHDXh3w6pYJRau0lIJGCy9rtRYNueYbuejQY2Y7zLNnj5jIL
88J4Ul2kdtKHvsMF0jJVFHItgIYDYINSJlaBNLiXO/rlknmoPys/fSWmnfyBMhMu
KzA+wjeQjmjZjJveBOtyEiwsKzBAspSrZmtzrVBqWaUWX2Rr1LFNnrMTWHdbRr67
bWuDXX5ZBjfL3CrPp9MYosWHxVcItMYJyL6opah4khoDdtaR1KnmuN2eqKKmO9yw
IpGYxMia4MxmvJDhWjr/1kOS+ETW5VZkkJNldzQ/D3YR4K2FS0CNATyiiUBEZ2O2
HqOA4WpPGGXt2bTqSfq+OfVPkux8ZgbVX9xzGS0wGglrjSnkHBMWS+9Kr/2B736K
P1dhVvUuEskADpZgTgUwV0bm//Hh86sk494vM9mSNR8m7yMyOMtr4oerI7LBi9MQ
tNvEtjasvtrCjgLxUSqeB3QdZyklJwZsdMCrHTJ2dqMw4BgvWxIH3eznHLR0fJQT
TmOoHFi1aWtRKp7zl1Y4v6rGCGYgbjJ6xb+R1mpo/LjhrysFq3ctpo9/TsTb17A+
AiwloQT7QA5Yq833ENC0GrXkatrtlmllTiG3+U9OHc0updXu6/OIw0y2OzpMUcqo
x6aIVc/JFhYJlF+t5Uj9TNYv684k3xu30Ums+cjnOSLmVOF7sAcv82vrPwLEXLic
RezDTpI5JihtQHFbrhOrGmpit/8DGoC7UaBQJMAxPNZcPFCR6/TRJZFEIU2BcsgL
hWHCCY7mzZEhQFXgr2R1frR7nrNvzKHYT1eWHpqMC+qq4F4gVqNpowyPpMYplLvr
K5IJOafarjTsuG6JU2Av66QKSGIiHX9ohboYqCHWzXKrA7YrLLUP/yYp+knGivRA
9ektVMbcRVdGn2KjfEZ3QrKUybOeTgd6cQR3Qq6li0fuabOA4u74N/4Sta9iPpXm
23IlqGO4idnKlwmTB+TP2yI52NOUUSh7usu9bVxTDtFt9f3GhMJPvEGl2b+Rdz0W
24Ag/dtO8yzVx3CayLVf43rNwk7WT0DnTYbbIW4A06ZMaj1qYCE7Or93BM2BysoE
DWUlw7SIGo6IiPzi8JKaOSM8dpeMsEfCn8X5mzberK8UBjAVvqTOAwOvf7E3rpSW
zbz8/xuUmKJo52G6XTjoJRDiC8O6pUKoJTuVB10OaCgahZ52vZtyC6jcyY7cL9oV
GhY17mqCkTubalxdM/mPyTFGfbIwI9DVGrau9LNdPcKY28IUE6R8CRrcDgUtJzbF
HJzc3AN7h8zYPYiZxsFCjjybDMMIZVnBdbogSiQxTDNcbxMWSKTaVDoQaL0n2yU9
OQgZjP1fw2Y7AVTl8U02NLFXO5jz3zpRb6zS9DTyYc/JJ0TNGHfO4mj6zECyM4On
KRvo+nxKKbFQ24Crt1ScHMe+t1QnY0o066W3XnsCZJVDSCeqhD+N4IKA0CRX75mQ
wf1PDd4KGwZD0IPGu6QNNIwb3/uH0e8wi1aaBCaLYZmnKlUOoxysQN4hNXnXfgrz
O/I5N/VO5FIRQGOBXE4Nj4I5Hs4EQvlMEkFJqOPfsDryb7C5IPkeO8ldla6xv4rS
lLkfeaxEz1f+yovKjd2JdmU1Yd4cmtgzHr3Y75l2+BR13Eu50HJiNoEzRWGcihfY
0oIPzmGY5XKtm2hymeYvCOELRXt/vpyJZsnTU6Ee6BcYHCrDXQKzF3pTu7TZCSdG
g+rQNEqf96Tokuvq8f73lWwkzMx7wn4Ez25bb56CCMhbkRRr5/nvK6iSs3KPO2hc
kglFmyIO8PK2xwFOq8U2jpYkaqYgnFsTKRvo6THnD/s=
`pragma protect end_protected
