// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mSif1dRdwl9HU3oAJxwfuPf3wI3m4LwVnXyDlcD9lYsuXbBmtI3dqdd+XBByIPNy
fQVrv68i8ZXodt9Q7PhOflpK5NPtYBcorURP3+43IHZ00dfd0lfDwOjyaz/fo0uy
sbOZAt8tX1vA2iZ92s7eeIzqFV14MmeJTUZ682PAJQQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 135456)
c1ZaP/a+mETpzJ7dihEWWfSI+EObD+oK/2SCjgLkAPGvInRGrBtMPNJG+8liISkZ
WTViQuUPLe4mKnZrPHlntY3at921shheqPZKip/gqiq5KnKA5zZBGEcXC51d3/Ds
FmgWlKCdshOOvsBbwwGhA2Ef8YSe8GvUe9SL4dr6W0v8L1u6oYUq/fSTUAXID1le
c0MgkJDrU6ztsrwisz77SBOsI2L+TtAhWAP6cDPHPIMaSsmjGoqg1GB1qfG7r8Oz
MXPIb34YJ/ovhxSB9UuMpegFQUupID59GaHhHtQuWi7FCVbwGpWxfwMAzZ7vfhik
R97aR2GXfM/+NaTJRoO+Ab+2gn0CQU9YOrHScecUKofQ4gVQWGmBFS23rLn7P8Em
ndpquWwgMBdA8+1Zra+jN1+ldrcpMh0YWxxUaljBa/x3DTFVzdwL/7jdfGx37/Jx
4NPRmauYAyMTlXobbAC3QJJolx4h4xTpXTIhgASMZGLLMIn0ei4Hv4dPuIi2Aty6
mU6xYWN4DEGjGUcbYZ4n2WiyyesRu4hDeL3Hq6GDbav4jh/93Wb+GuSqtHyP8NWF
lx/QB9SCvtoqoNbwbB4rY7VjhCB7HyulpcwyI6e3m+h14JacaPh5ZXgEGeQUOzqC
HW7tmjWOPQ1E/JmjvegYUF9isP1HgCXJ6xMLEXkj4bSLCA/IYi8kjzR8v79p6TUQ
YtGnIdaxgEXS3bPspBJXOXwvCLTN2RMY+/+lXjZInKhVus0beVvpRcwsz59YoCP3
dyu7d6/H5WZBb4PZUNIQHOFS+a172pwPYByMnq06Aeomw7Be3BUgXNxPIbMUU9mT
eDjbU1kmelZlGJscZlPeC3v7OUqikAB9bSr8JYgKTFsoCkg6s3hgStGBmafDAT28
4YyrIgszXiDZp9ppGzZ8d7E/F2vRizTCmroy28ZLQRG+6LR7bv/5/EjNed/N2ZyA
7buQ2ucJmpSZU0msH6TKvENftdUvjnww5pe5ZJY/H4nUrk2HfFME+mAVvgaXj2tB
NW5YvsJTRG1ZfF5pIRncElwxgoZUnm0itZXkSzmYNdDKEWiXRAbl6VCWjIWza/Y9
qZ3yxVwjjRUoaDUg7nnVVCxJ8KFI3oHq1XuXoQP0hFu2fLX/r5ieOli5aQptlhD5
+b/1/KxoAYlPlsZSiaS/267p+FWsyUDV2LbB08tw7XRG8M4Ew7NBB7SB9dtCkeWo
Q/EOf0fd650rCiSmY7q/DcTPgIA1PHc+tLrvRcWhkmb8x/3Jc7rOxmh83RryqWxl
LrHeA1EAi7qUr2gtWk+PyCHHb2N8d8iEpuLLAB4RXAGAN2RBKI/oPdkWbHiHwVP9
7OYxDsgA5m/6JrEYpEsTfCMTItxbTbl++7GQre6VN1nqaxKKfXru9keJOeWTtaFn
U9Pikik7cxPMwpsMFCfcw4qieMr4cpgX3EKpbQbbxAeWy4UfEIyErp9W1kuQHjQH
PmxjNXBHrCdG95IuYCjEihwLjzrxhknmbgRbDxYZIUKlPomKZSs7X/OQ6lqa6oV9
6zsR3gJRzTVuRVk82ePEJaAZTyOeznjng0zMEThG6tuMm2zbeavxuicS0+5ID4uZ
SosKIHlKA+TqOrdDBXMDsvVrX3wKTE8sSaUaEZoXDLbHEfCfgy6UhG7WKhHkn68M
R/XwdyAr/dT21492O3fPJIR4D+ohWWX2R+IRsmQiFzRdT54uJddXbsFPMiKqmFAb
B97JFUIW2M1EpoqFLZxlsazMhZA+snKIP2GsF/QMugzyqIFAgsV6FyjVr5zHhBMQ
7+Yh5snI8EGKa3qj762PSupvENE7Xn6tRJ/I5kGom8VYboPzfnRsd2CH7wkHjsKC
A+VPbJRej6OebxiPwCpbOsaGGsLrc/P+Pz/71dcAUGnq6YognKvCjyTwDVtMp8Uf
Mo/xJOlZMpRWLxJrFkRsN+JKVM2yJDeSrn1+DqXt6eyF915t551MZyTylRfE7VMC
qpUZKtqKiRDdXt3stoRhtPGkpli1vD7fcIL+R9ZbhwevnI5dvHOKRyPNXMbeLC9M
SU0scLwozy10rAVDQ5cYmm00JWj5djiAKqp9hOZHbObZx5+iKHVyLeXsgdIC97yU
Aogf4cqaofv4cBTFkqMJrAqdPH5TSK/iUkELIzYa55qFBmMCMqs4WCUhvt2O8Tf4
uH9t23VbDqjIT9+g4LLtTNKi4TSshFbcQPJprCZfbLq4gOGRYFWCifOfGKMjgi0c
6zYguEgo4mRmJXUF9Unsih3MJ/JGj0SefySUp4/S97524g8opYZQmP+TvmQU3C0c
sMHgwieSsqqDn3TGbhRDQOCqUWgx/letZnNeF9uqubM2ExqQ9h6543upKclllANq
xy4IGr3OKeSdbK/g/YbpC+TDjEmEALKNN3PDpQzlCQXM+dBFqGLVE7whxY7otDTi
0vsf9k03aCVazXVEGvQT1pKZXlQMCiahh6ha8+29Aiy3ewFVb1GDCmRktfuGQY6a
0L3bW8kL00nv1C8TS2Jiwy4dudK2yn3AS15UeIFwm4iTCVfWGJjkT5g0YfD6g2KC
z8TSdJ9uT72sXWVnQthVnRpyQbY5hZs+5nJ1NmINRXZa6L31PPows5MCDNXAKHG3
ZdHbFTgCgNXjIJH8Np4MWB3Wt/iEodptsusC2ncGZRpNMJZlE/0k8+NjZeNACcnQ
WjuKrsp93lfz4OHi0NNo5rWU9zkofbbm/jAKkSu0TVyuK7MFSpXjOgpmYNWeHIec
G4yDqmuFMsYPoqhQWYqJVp99M/JnqwQ4bkoXBLMqcMIlyIwaPy+AmSWolqDva5Gc
a7xB3zUZfZ2E95IWexm+DRjkCuEZSyhyXnXRyMcjXIVtToETfKanidqboFmUpYNI
pmsnXbXSDdAX4P7ZDLscOVJz7aD2uD/Kq2OR+19E4Kd6w3WqOthpqbsuncd3TOAz
VoLsCfH4M7I9vpdkONWSR/JSnsEuFo0HoxOna3+kTRjKmJ1Pz1R9Iwdrm3fieAwF
wBZ9LcYJN2ndQNzoFJnek+SlDsuTDTqx4f7W/8vm8Wu0DugGux1DgD8c7cAjyjsv
pXEmv8zjZ33F6KePZZlsY/Ifn+KexEorzWjXkJ6pWwEPc9aIu1nluYPOdepcZp9F
LwZ8fhXhaUaZlwzqcEaGCbHVjMP0sN7vQqb7cCvSm4PgdL/9lczPk+nrz8y1VMNk
bD3MAI7MtzmjtGkj/y5qSng5kALh5vobRvX79xK+VrcRrzj3hyJ93yzq/2zauSBa
C2nrQvCcZ6TdlS32JVLT9EbJU/ei0BBmxiVc9iRK6+0x5+++p3rTvpyAwPu6QJai
JSeuhrgYhOSiwV3ASFRDm/xE7jHCQxlgPVNM2yd5smtFj66xslxMR6GoGd78a7dP
p9o2shJ29Czp0Fti76iR3EyDgGXF2BQQAa36seb21xGNCZJ66rQrB4mpYODOE2wY
qb64e2lQcSg0FW8He6Agx6nZbjp/isr3/M7oQjuKKxf7Wex+41lyycJwrX0NVZRN
3aYcgovd1ncu0JJYm0uboJkp3XNGOfAaEhQ8n62IS+fKw2LPix0dGpazDyGhpM1w
qpd7MkyDNLVX/0dDCcnexgTrWuJ/p+dsLDdDfhg5zZ8+AOMuqyB9guYNjyDrOcoM
nZmepK+u69a1gF7h931F/rJMdGt5bjTQc64K7d4aDUua3kcwTXkxRMN4bD10dwDd
s9jbXMZvc+sGVecz82x4508eVAfuVgKyIvRowkwvkIaNQPmzh9SIkJxs5xEN4vJh
Io5z1YW7RWNcw41agCmr3P1ihZPuheQXa81DD2aVk/rU8pDEH2jZJkKkC1qc3afY
UkV0xu6CvX1J/VZwLQzhLpzPvw/28qlx10bPdxOPkrBlkhEeSGrF7YTUhD6zQhXs
tyt/1khaAoHdzHu1Ba3gTAHaCbZpVtvMfPiiBhfh2fuEv6526Cw3YF31jvdzx0Z1
kx63P41AsvG/s/C9/yhqa/HOXdvcKf9gYoVQ9jBiGXnzas7DwavKEpcIeY0n71fN
Gsx3370c1WVn4a2HmRJfr0+c9++/FefvRZ+uoVjnwxVRnAZmvyo2qXXXakfiirs2
PGb40Eg+WX1MXb9LXGgNMRWtCNBV5+/P3QigUo0FPcXS+oR0HQd+svA61dEDrg+b
aqr9JG57HyzxzTC3GH3NC/DrNGx3xrMyNLRKZ1UEGEVPdRQhMKWMK14EDCGKU5Pd
P5p9q2y1V4Oayth92ijdrXqQU4BC1NK3LGfH3nm3ormusjUHq4WBYRtoQkZU/w30
jH841rpoutA3mmNRRSaka7pxeNr4G1UhU87rC3aviYiluG9g/SF6sci/UuspllRc
EfC+Fr9s5XWjj3noCVSqfwdJtz+SBejGchigM1ulKtGcSjQT/nhU8EfblXIxdpSP
ARZXNYuQhKHGATTGXB96MPxvksFCuqulmrEGH22Gv6PHWIwdTxODPVxw3quiTlSZ
zbJqSam9YB3A9hwq+mvjd5RLHvBoefuvH/aSCE3L/WW7dWbwSBfmqaoWSP5YVGgD
U/avupQXm6CqsGstXIkC+nTwqLxfHVUb4+ju9/sdxjhcC+9oyHBPgXb2SxzeKy/w
LLWXzVH+1wIF2DqPJImJ6wmrW+58jWxIw8bS5uUPxxIK8wfTd0Apscb6gm9yp+rZ
e018/YbV8tBaZRqp1pvlGr/DQA1tj+A3qijRVjAjPQkhsc9ON4Zhx7G5++eqP1gl
g289UmAHWjXFT9Pz3agNZoB6LFqycbLuScOjxymHI/kUn5nfh5tvLh22f+unwdGb
MP7KjDQ2JYaBp7fdp8ywviC+qosJiqCRTBHRzhOENSlsFbk7f+ytxyarcOMkegp4
21jcsBFoSXJ6/y/fL0/a9RmRBv5ctQU2jRLXvBHtVKl7IzegOQqLciEM0Pr47nXc
FMghU5g2S3p2yr3fM1ZrqYaYiFKmT6/GCom4kZHRUZKVcrB2Ir2UTA01vzpBukvM
uzbe2/80tHVgKAFA5M4RJMQuM1/HVMTR48wRsC5+9M2uPVw99Kx5hR0nwVF1fRlS
nZVjPvkExkkmBpRAOYjLHWeodPPLQxnOdWzCxYSkl/t9/ozBCXrVkWaOeCPIKZYj
3Gw5NDIoXmwysmTeUJnIR9EgdUwLYN8fZhaYvHM/uBkB1eWE+5Y0PwOJcxfj3Nfz
43Gi+jecadn2rU3moXdCS7WnZYNKlM5PbcKqSbEqwqx2Kq8I+YZFAAytLmQ/my5d
N5CjNGyp+JKXnAeoodpmO9/pM/QrQbreBGbxVKbXDkfmCirpWoAY/6JRrJJhj6D0
3PxazdmypqV2/t1fXWDN/8yl0IKwartR1zDtDrd9nPvnMnt/iMROQwLcm0KTbo7C
ZumTaM6yOKZBZSowXYqwQ0b2u9051HVgewDGhXoHSvRD5CHBw2JXL6kVj3VdJMmy
1xi0m4vCEVZYIk4v5ksOVaZSynRySzqwRZLSz83HdOLaT7On0nGRsJVrYmTwmdnw
B2zMYUQsO4/32RznR9erRzzQAsaViYDNzIisv5OHjXcag9BflKJn5hVVqVW2ssls
Fl0yI4kXM4B0F5IxE/W6zoWIRyiyZZBDDB41/u1Vn9Nh9YtoHbIeLCcn8EPTzIrB
KHlGersmteGflbdZJNNL+e2J4kb/p0A0usNxUXcLJS9rl+OiknuBRzr2qZESPBXu
ig5f1xzIPAPKv7t4MT+0/joNCQIMsMy0lZqq/o2SPNJZKzvNb6Utv5yhPNvBxXyn
GxrP4/HL+OweBqbnh1pf0bFBGg4B8ADgZzyg9MF8nlsZ/ZG3pddIU4f9rUhLPQv3
1sv2LVlJd77A0K6VVb+6bq/41yC6xFGxFverCQ0+4+QHfkYQ47Da8678cIQCkwUK
6rjt/iHSZgJGcRnYVEarHq/VMeo4oHFxKORGIBzuhwIRP+oLH9gn4i2zvqy4m1io
GVTEMv+HsWXsXLWVuge2+E5eFo+Jpz1Gj1XJ9L9fp4hVFNZhmwtblpN+wqrzfYqp
gYWeo+wh8lYtFNuhbMiwCG0DiRKoGLrCExxHD3dEwG0c+1J/kzxKV6QLH7bfE6JH
BtMNk4PNK0WMbiOlDKKzzy6D4wIa2EGeQfvu7Yj8tJujY1jQ6HwdZRAoIxNXGv2u
TlvE3lzJF8kamnsvngfrPeh6kjmm+t2dpMsxTOHAycZxLAcGtZqUX+SGV5VyxQ44
PSrrjKLfNQIXRuXnHzyUpGcPb6t3lwCNeIVajJCDNx4SurUyT9cPACrt2Kn33z4H
+bEb4CLk5xDHIHxxiEaJ1d4lZ5x+gXomVZd8w3nUv9SLBXcuWetCiW4b5UP8bXz6
iyZxeKDn8Fy7eGUGArEUNCQLr+gYL2+5cpZeVUgx/n0ytoTrwkRrXwhGTL4c01ak
N4p+jERRjK6Xv0eEH7ehxaTDGf41hIJY/CfXP5Z8DdFUNHSbA1fPtBHsT0gJcJ9W
aGq3Me3y1W9Bu8tPqCr6RWGH9DCAPjwkUBM+vtlaXSX7s9zku+dpAT7CVE+vuMWP
LPiD2ua+nfIA7e21EjsFmaWHUPwRqc4AkX6HgS0liCJMJYxTYisPk6Hh25rDO3jR
rbjvsxp2bem0n1im5dbqz9tM+Ojg5Ffu3omstFrMpczxxqEd3cxCPBjLagLmNgVC
kYKJWteIOecx6YUrSFPgS7F1J1tB03duwJxL/zDXlENKDz6f4zDW8220dN4xp6e2
Y+nW7PQnUL6FR+2flf0HqhNgh65710rViGnELIo3fqdEesi4X5Oij0bbyvmVv6fT
bzHAlzFiCwEOVHwCRemXwloEukAz++ZsqpralnkaDfrXw8SmklFgJfzCadwd8oB4
786MexhBZaXyTPNQbp7V+be/u2bpSV+TpDfhEiVkesKslJj3dCYQyfdVdVtrM7Mi
wwNu+J/wOEM/rIPZa63EOjeP+3As+kzpzoKiWniDUP8IS1n0Onchzr+Ms6kMfdzh
6BuugW/GEremo95nYr+8oB+TnS4jaU1z2gZEGoHacnp5FpWCtYky4Dk/T2Mkm0Ah
P/zPhmwUgz+86VIQFKSs+X/r4Oijfk67ouOGecyH8M6/M9XFQ+E8HgdskkinFa3z
zJaT/hEoSITexd+yB/TcnVLBtCa1sgjJXVzaidb/HuaskCZW69RVGHJ3jXjJSVRi
xvAzRJPVZBk4gf3Pci5yItX+VvCP6unaScUUJdyxKfMglmBHJfAl3QqioSeebD8x
6IlnpuIhikSuPDNiNksfu9jcMreEoLFAjDZA1azv6wuA03kXynHRbHTK4YgIXWX3
sq9IhIMCwcqfHYFIt4RuHZ+xv3knDwWx5t3N3E1fqP1f4V9P6HJsYTxCdotycCw7
YvZaBr0v/X/pVUdUKTRkPdxqez8DnSK9qtDfvQQqcFZqWf4/rbR64KtSaAnXfoLZ
50OoXhC+i76hbhKQLtjio7DlWn1577xYc7N8jWVySx0zCRHsSRgMGZ/qrP9gzuqz
eYb0k6vlp4/h+CvWmhQrKCam5BZFb4BRpgq0bfRHkvthwLxOJWOfd/XjspntxD/g
hfg1SbrsV22CgwMNL7JFYUmzk49/Cck2Xkf+oi2hTZZlQGN499Jwcs1mjFbBMXx0
CiVmduf6oFfC5tMXQJAVBU+Z1x5gNlE2A7qAsd+0pdUOELGTSFJaSWcjGdIKDP5w
NzzJmyuw2RlqZAfWrXSs6OkDzmsQ3YC1Is6BRi35DLRZrKsx/sVGci/nGt7Bh+Wt
hJeDaiUm2bOeOiDFCD6WWYBt8NUdgaVnVlVQ1k7IbmnmgsoebAu3tTJfN37HPmzi
w+ErVo8eQY12kUU9FMrEDlG3gwQNS7FPa41+M37TvBlkH3H9Fb24epS/NJKjqso0
lIb8hT9+KNaBQ5Y8BN/pQo3uwn23aoYZgPLeIlWb9AwV6I7o2a3Xhl1TwTWSf6UT
KIYtpf3My1aiS/zkm5QxA7dG+wDEm1YaJPwdRxz3RrhJWj2M+hY13Js9+MTluGiM
W8W/0kH+RbVw2kdePXq2+aB6ldHUX3KY2ctpjfdOIuGfobPwJWGdsKZDBZvGDXUW
rUZnlcfpS0DDxSJiqz4p991fjOApNSp/PVnxLdZKQlR8Shg+5XtkDSVF90uxxQxi
c2tLpyr3vesyethi3T6wFCMZxVyLr+gKb5eCI0W3wJgROOfTFipd+GOXfRR6RKpg
TyAF1Gn/XlUE1oYVp8i+JmVINo7WlbWCTr6fDFknNBPyuVi7i1dQPwOU2St1Ae5c
so6X2c4gBwOTjQh1GKnc2e1vUpOfeRAShKdqAuIsqsZHaMfTWNQ7Vx+aMEXEd4IQ
Mjhpfpz/iSlF+7bNzfQ4y9yZ18Hxy/NmRpdP1Yn5PeUKAlpgGLvhUejHoQwbL/tx
zKVslyiIPziSiyENgkRNP1COTgG4T6Dk8AwbBMejN40YpOhDXEAvQP3HE3njbgqS
g96pNXcP7yVbdid1ZHT7souid/85kEo0ErVQY2fih337Fj3v3ahujiOCFPHP86J+
2SOwTDHBjKyyO5IybypLBSiRX1aHevsQb8aGvCqaDaSVcNeYOSURJSLcGAkOQH+R
WvaQHz9HnRt4rllvcPs8Q2iqZqKKU3B8KBZ+xNB4TTlWIBN/Cgm7vDB40napJ/ce
enndpm8Y1Prp+hfibbJeZjcP/RcA8C6eRsbCFgJd5slWE9kPJ1sr9/wyP7di3gV+
oVKTzGuPzuG21+Bxonz1srFAUOv1epumQ4BXV+AQ6lL2ofhrqcL01z0lEfaYDF5T
MfQbFuUFJ6LzDU9X5OYxsGTKWfYTUL869jGWZS3xSbUfdIWyQwkP6hjsT6kFqWcK
MI1NBGeMX+6e1dv+/Ra8YJ4OJjZUZP23aUKjfaJmqTB0pyi3EnB+c4bDvcjfeiMV
IfAIwRaZDlQl4USgih890s8VaW+BdQQN7w6d3QqstezIyuP0oVjc5z3DFjvms1ju
qGhvRHXs4FplABC8KXdYFYf65DtYcmaJJ9O44VKagyE4rSga7txmZF+GatbSH8bP
ChhDrOBskbQBNK4KiEZMOr917w4KC1o3pPWh+D/cx4votyqRPC/BvxvguovKuJh1
qe0WLKPtlm8ftiXnMaYeV95M61tbhxwr9Ypry/8whNCHkK2BZaGOC1un5wzwQbaZ
VOVu7kB6oCsoiVsn99XUmZFQ+MeEGZM/JftCUAG4dHgXNyjcR0vzuTicknSS8ZjL
O+AXkCYk23YknRIqkEJOKWWDdxGUF0ejiE8Gv1F+05NRMB7sKHEnMtqRwQIQbOqs
w80yhk/ekPfpEzbAWA1aKt7bW1ppl3OC1O9wsGtyim8voUTeYTZskbLLziNxZ7dT
FgXD3WD+MzFBSs7FEQiSV/yqtvqS77NPxclr34MsazGpwQlqPZ4VTc7nT4ePYBYD
vyACclnQE4kkS3dyB0aGw8vtabk9M/V41s4M7fE6E4d4JU3CAoQh7RdwqZsiXbkL
Kz6+DLO0t8dj3Ou8iGj7cKGXqUmmu3W9MKzk7aCV4v98mg7pJiz7QKTMaEcWgNYq
OukG30lyLBkOR32pnNlVdTmGhhr48rPzJNIbuO4Aw2WUkFzLBvHGOKCkO3NW0kwn
ibK+k39MLKtBDmJvDL5Vn+2QlTWZ1iiXQpfXjQ//IincbJAbZ146Xj1fKrU1KsV1
7DQSTP8PKIcNTzXxRTOaKjoj7I7ZmoFPitzJRZAtC/J44k95ZKqvPYL1XbnIoNmA
GD8722DBqq90GKXQxwsGJgXHsmZAH0exrQh45lbJJiMWS8kEgqz5b68Wdjfo/gY/
gM+CyWSNNBiLGi97fpQgabHC2Q+hfCfI7BUhdSSybTgWGWvCUDBW1w+4EfQ8cwZM
vMNX5ebBO77pGRAZbWhn/V0JEz1rMz8VKLvcQWopKQeIaA/hHs2DHsHwQGACSID5
QOAe8siLJ6qt11L57IagJGr4xRaWPiwzHLcIRSMDuB5ibu4mkVzW+v5oqmJJjVpD
ktE1f22/dUD0RIr2XnNJ2cWQm3zRoWCI3pyeWhnjM0sOJn85Vad3mEwzsKGg5XMs
5mE6D4UxzgpbwxaL4kNCdkxSZ11NUJ2PzPFi5eHziHracO5E6DkBr4iIlnkJX1fU
TegCHLTdw0Gb2UpIAi9tuX1wjCHQsgSJF5Sx7s9bfrcOloS0WxGdqrS7GB71Oa1Y
nW+34fHnZSbN/YWiXnhQ/n3IvvmGIs3WtxELFtN9KD5dfGKjgn4dpLp7NAh94PzN
pnIpJPTYkMMHS1Czm951o3wlpMxxUrQCRnGCuwP22Fnfxr0HLFvahDYSLPrpeu82
F7Tz6dyqRI0lV1x5ablbRdopFUnOTcS1+/8dA9Dc5JtGr0TFSmA9jC4ndYhuPLaf
X10/2dLtB/fqIVGtxsWniQ2IV56Kmzr7Baw8XWOF1I+qtGb+Lvg5b3OqfPfWUYdC
q0FGz93KQw4Xu4IlCMAVUlLxwAewMU2v1tPm4FJf0DS73pQDT2jWTRSW98UahQUh
jhsgQQA3mwYjrRb1l5q3tulg80MRVP2GkSsgoDgTOV25ALG5qSOUgSSPHRDaK+h6
5URs4MGqBEixL/qjjg/7KgRUzNLxETUhDAqUrUrnnCH2JkTDkc+QfsZ4I+gxi8Jv
U0+3TbMXNQfuE0Kx3bDWJKvjcnX4eszf5NA9KmSVlc1ZbzfhYEBOzrFcvKklMQJf
xkJVlFdjsGIfSc7e6+FmmN5v/fWpflTstyKlnEttDxR9TwM6uET9VqJXbuZ3GstV
9KyNyIzOpyqXNa+h1rT7gb5N3cauRylQcO3nP95rDlu7Wu2oWrI0fArUQDXHbK4A
8g7wd7zGbSXcbhQu9OoYTThcnegFfviBKBxlKZpnHjwbMvM4rabb4+78Qh0Hte82
npgidrzXEu5JmJceAkEj4yUO1EsZJzHsB2+uKw35b1Jy9GeruZT5UXAsJeS52BaH
GEAEsx7HfKWdTsGSwDLklDBhJdoiV9C3BQrsCjO99g5drGklvw2yklNf9HOthanN
X9cxyxLd0xsgRe5O7PAR/kTgGLK1FfTJqd8STI60IanhtKr0cxZl3lzg2wJhN8fo
3uRYBfyJhHHpBe7Q02LWMKyjUSdC/A6of04ctljJo2dTh7adPC2/adBw7K2jkU3D
Z+UY6Y3dduDU2YpytOJg1lbl9ks3mag6TLhqQorhaKk1uhv/UvfxVw7FFuOgr2Xx
8XwEn4d90PskqniDTiLXBACyfEAQHzPuULy6t9nkVOUMfw3kuKgWQB8tKVs6nvLc
HGRT/IsH93H8C+nVSQsFTtqHSRC1hUGjCf1RBH0Egp5aPlwbEgztXVTkRIApodX2
hBIJv3l+ls5mWvBHP7UI9iCaDws0rlpxGMwxW46wn3Z+2JJkdyD+k0gBB03QG30e
qJ3pILCnrnHn8C3noqssa2nFNDxUDd8uN3lcmrzLksZI+kar6TSIc3KWjvMEmZbS
Xrs2lOCEMr9tG/P91imGTHfvqHEFM8a3z85sm09SKfEhH3wfbBo13lM8KnhK7lxH
NTMF+zkTu1pENXZU5KCBgjRU/wX1/NYwmkGxvxJKrbrxHYKSX7yHwWYiJAhXtyVw
LQLD/Xpw2KPLWO4Wyd8/q5QGsyaly5zw9+6jO9JECEGglb7bEAQNOc93oI6eZ3Zh
hdSRdVgWt6w9xf6SvN8LU2ka6SFXj/d8vMEGPpfCXtw+ATsstpOB6piZLO9Hdyz+
CuX6pmrBuPye/Ac69uCTd0OAtsja6t6fMFe6bqvEvwjBD7QeqAaADzQzm5e2VYhn
qmGIutTTuRU+pbfFtrJ3RpJ1dMsfJKBHONk0fper9Lh2SWxTyJIy0jskdrgdlnVq
AozzBonNDEZJ0rJcYmXu46rr+j3oplAzsP0JNJZmSuKokvWzAU/MOUoZs9/rsGQ6
z9WuqaRie11r7xziJeU9wxNLFj6jkHUKZCmu8pxCDfWNeu9Of06a+SYHXfiDyzE7
3tAiFekNtwttknU7TNtAqoHExIPCZKR4prjAax4f2/+prUytNFhR4yn6zUdpDLx5
zXwToGhMfTkWmgD1dCQ3EdKxumEVS605NljfPeY1+N9+rP36jKXTZEPuyetY7yBH
f+MCV8JSrdZtGdAo0jA+ghv/jEbgLZv1z8/6GRDEr4RIT2E+1IioOuEN/2y+K52H
BOGkQslvbZeAeNNbrTJtBSyjNFbqPtU5ErbHAl7164gi2BEPpo2a1UzhU229dl8H
xp5Tg+if5+DGW72ZDg/N+2hFAwdkl2XZcDE9OU8XGwXYPD9VQO1AQgRdp4QQVgyP
RuSiGiIJok7ptGsCjHNrlN6CH3z+TiA1Df6m2deTnIVJq4D0/mLUpSqCdPooeqGu
vfcu9nrN8ODXzxyCGmCqmh6FK5OnYmkhVfMftS1WdE9hhjFkMQriWNdUJud8ZEK9
tiHUkvorW3/S9gjUl/7q3XP0JfivyJ+m+ic/1xZWNtclavUBu7H07gzJ8zzPpq3n
s6Ax4Zj/ATQqNftzpNvG0DCwQv3kOWKT6VwjK/v37BqnSeKOMtJeKr6yIK+dPfXn
gvuhVJTocn5lZi7E46g0mO8jCfZ5Go95ToB1oT9Ne1eGZLJjIBB31lsmmn4RB3vA
fuTHHHcDwFtEnNqC2T9TX3WM9woRyjFgAzEPmuDFVo25r4YGlB9SYwkVbJ01IeUd
nBWSGgBqQSoi0r+itO+gVwQ68aIxtSsjMJ8U1cmgLZmN63FevuAcVjEBYXRGzY1a
n1GBxvlp+W2GRAfd2a5Z211Pa9r0ZBI5xscrsjxibuLI4OjiqpTmESpo09+IqDtJ
bue6eNfSvmUzF8a8WXzd5qIfe+w5UeObg0FoMOFCxoaII8TUmJ3mPCqPsDzsPpCR
Q67rS+dJxYx0BMzlcvPm0eFY6BVcc+arkFEloq0cM0+24vif1hZyoZ6PFVQ9O2Mi
WmgiWsC0VIrnTM7cTUCAnBUgCdKhFrtBHO27kkWqmgAzEyq+jb1QPvjPWgvIrgpE
oZgigX936GwruGExptMU71Vlt8I1oRx4veujGjgw+e3qUXPnzAEIXkxiHILiGrts
szHNK2bULfZQdO1XGQEfzDKgWdKFedf42jflmysx3U5OFZZdx00SrNPyJZtXoduV
ZUOEMGv/KzIIVsZZPhBvlRoAXWcdIxEfxyYWHvTJWWxVSQUhBttTHCibTY4ZdbmL
RCTK7R5WY/6HKeV1gJSRZ9Wn9hbWV9/cuR2o9HSmTip/bwDLy8YoFsuWeSo+lFTp
ByY4bNX3NoEiCUbChvSJXwHdFj2TWxz6/uceFLJduvWhvVxSebXP7+uqSjQNlRmt
lxOYG2enIWhcJbKegXzPzyQ7qzySqSgKQX0rd9wxRUA0+S0xPjvl+3Ww+d2jNrWl
TGJL1fUae9ILjZC3EM7nMCRazBLP5avWlEFSLlXnXXIN52e4Fkh+w1VkRoxC+FhJ
jGp/uSLGJrwSlVBtfFsLJK2C1OF+Y7yweq8AAGLnVtABJgNVBSPAJp9wTokEKRDL
p5dDq+pgzsi+ZEE14gWos4NqDvreQBJnHIdu8G0NI32RNviPx80cSBMyX0oAkwtb
0Mza1owdhHNP/SA5dN8bU5Iel64/wVx/2G/TTNJXuKb38Y0vAxuFPlCM5P+eC/p5
QXFLs71/hz8JGLkqOg2va5RJN0fA76IZYC+0iMWczLl9NAu8iPPYgx6M+q8WomJd
HgeIytI+5JmGi8SCGawmRuDsv6NdpUABTZHh5k9dx2KzaIeSVTdO+qd+Z/UqiGmJ
PsO3YSPZanyuHbLcECOZClI1o8iroUo6jAkMt7alQyHe8roNYnjfTbzrff9+8tlO
00BWEZu1njU5tPiMNzH/rmi906d4ttBJVknNwgGQwUgc3C5oZd8iSa5A4uRG8j4D
VA+5miFBG/dsHLNGyaVIhCXUefbqIple7/0bD3JGoIoWzwhOdgbhTZ9MR+dWn57w
GKVGmWJdYekyxgkwmhKWqvwAH2vzPWIiCk2PHqZkLHpAyPQRC1Zn4zDW3GKS2CZb
94Rsa6ZHb0xIENCEA+wNu4UUYghNKA38CUG3TYFbkIUrd+3rfABdvEwUBwiXpUo3
3PmQ5cZkNsFHrAcsAkXy5iNWmtY/QIGoDknfEv26jdwy+hXW2hL44Z7EmKtcNwov
4ftScM9xK7rTja4bNR/PiVYa9yPV+8C8KjpgGe5Jn67FtILGyLHJaSWln4nZazay
Za3L7b/mVQPsNnIFBMghbXjNWCFlrAgeGz2rdGR5Z+a7/pE5HweuKgypV3ZP6C9I
YknmqHj1NykfiAZTn9MClZutXjhruKGoaqE+zNAUcfANC5w3X7P6TPKGWZkBFEnD
ha7lgKPjm5TayWwBJ0MJsTlZXLNKtcTDyKI2ENlmIsHA0snddPmXEwAVaXzKIam2
BGkQEeaL+RPt+V5HxmW8SHvD5iW4y1zm/y4jLfQjlV44+sicFkxuRzj6H2fuJKZV
G3Ks2wKXBlVDoI4UYO07pg9wXG4wRjC29bAqjYaDpWYTfbD/6uC3sVLArTz0aZYj
WpZ9bf2Zmnfd19MVQ+Fadt0NfZyTJzBtCcpLi6a9gArPWSK3sEPssJTohJUdEKJa
HEaynwLntSA4CiKTn9NTUmQZSxWkJ5qgDjBBNddOsF6MLCKoM1ZjddjFWPjS+tet
w4JMGYSEuZki2yo1iOvBuMGODzlZEEkHS9tCBJBZgFY65F0t1Cd2IkrT0AMJG2Ro
z18IYBbvYaVt0S9itpDZFLs7b14TbsPjILAuCE6OOSPARjx+tF5+desrQIwsxUF5
O+r/S/yabORp2o1AyvBVxhMDqDIpFzEgejYdngSauoPb1ARJjSXYw0UIRVFOWuqj
9/HyPEvXJcz2hR/zau+8cpCpxC53n+HZ2ty7RBK62NbEHGnuRFbAtd30IGKLZLjk
JFq/mESoui89gCxHslpXg8hwiCSB8SxGWfWIN/Qq0edu0khiH3kF+mFuP2jdIM5X
Gdie9A9PpHPkwYlPJYUzP04bG50jfPDiTQGHdqVX2lsCvzEG+dxRM1MHjRrXN6Np
Hhd6ukk9BS5uBxV467n0VA/MLrIXaG2dwHjTGbgnA+5cDC6QspQn2doBt/qUpNyy
eHd3Gg62+PtUfIeAomyh0gqMwhM4/n/LXITexUTH1c/7/uZMaiUdsDw+VB6GajUx
/hCaPm/NgZMijteF/cIJplNvfanbJU/tmQYX+SYYngHir66D0CdzvLV8COx9VPXH
hGiU3F/1Ttsb5dJ5b81juA+PsHKRtnMfKSmk8aFOyvTrdCrijY9qo5FQx3Y8chKe
yKezvIu8g2++1W9vAO+r6CNA9G7dD4pk+9l/17a2HKCP3uvueXPM95xBWbMop0x6
1SbDaqnLA0Y2BYGux8Lox7kpksIMmhgrQ85m42uFXU7kF/eFRomow+mgplAyjdXw
5Ao2nWfUuWtoZBnPwv9fdowzmL5ncxJtNNuKieN3UnMFHiv/PhYGVQV9T2pV1dgT
oWfV+xyAW8dh0W0Q28YNFBldhrJvP7Qxrk8WvnqqkrI2VB7In9taZYDahmuqNiRs
AtXfvwI/yytPBqJvM/zOOuDzI93og/zpnGNzSMkX5njJwaYmQMTJwU6j9CVen8fP
+ALBKWdJ6hM2m0+RQ4trQ/zu1AlJwlGmhII98eCCPseeDJmu86nJxOHeGChepnWi
3UuG0j0OeKupuZCKDeLz8vqlFs1ygmdQjb8wYoaa3fQwQOGEJQdgKswnbrDPIX/t
Pt2dT1SkJMk8uPcoHbaUqsMuCUMZ6j42VjegiVj8x8bWdXO8WxnFPahZqo94Jgtk
gT3cQg5/YyIgzRieGj34R/jG8EuGQ7tesoWzgT5re/rwo64mpsz74p3amt4XB1zI
JXwyhw8mJRYYh0r6QppWMqj3+C/Tth2aLdaM5UP0aaMkDPJylMmJzw/PSq99S14G
2InNEE95Luvop243uxK9Lid6/zv0XT1nh8WsgwE6006XMTFumhwFWiNdht50R+Aq
sCOAg1QWI/clpdITaYjhUEhT9GLgWJVjOhMYkC3CK0ycuW1DLDa+W+ajA0+0CeYT
KYwPvvZJqZSRhnhPgdRK0Ey6e4xHd2plaPset/C9J1IvgKfJxTd+tSY4mAl1G5TJ
5hT2yxqIw+ZPuJjCNFg64/MrnLh/A97S3KEjH8KeTnJ0DASd0rW/P6lqVrlVBrtW
hrD7IpfWvwZih3y1EKYQguWfR8d8ZGzxE5iq4si/9BIwrs66M/IH1Ixz8RvzLD+5
WfqYZAB6h6z3+sKpgfEZnIlay93yufh2kG2RX8OQkE+adfBhsblDnkrssm7EftjJ
AcnH2uO0tbXPQOgevmdMaJEJxWgefPRNDvDDEhnHZ3aztG72HssZpViRiGlQqsGu
8QvtSyNT/Vao9LzKVJ+4UKRAkF7Gw/BiFkS3S7f1iKbfpCwTVch8RQOr18FKd2br
DOPDspgMRzlZOGqkqXMnFQSs6rm6wV5iDafqBpkyYjZQgv8BLxG5WKzUwwapapLX
yHJgyBw5cVaAp6Vs2A/0ffUq/Gm60pMz/iFGQYg+W2Z11Jetr4AvDqavCCi/wxPf
czELVjP8NHe2FaA9KVtK8TJS8ZL/f+3gRalSiJsKYBbC97pHsiLEzdL10WrEkwWG
BPBd1FjI+KfrAieFjR8gz4xNp0touwp8I0iGvzvvd95gT++LNF4fLE1ScGplpURp
baMrSJnZdkZjBlOzYH0/bmfQnNGNekYHHWSxybYZMMyRjwO1H63PK6V4eygKL5vr
DHxrmSCDbe1fHD5+T1eXy3DiAChQcg3ww+VTTqYYveqKGWgQUS1sDlz9jmdCIQRY
GrJ5+vhae8scFenLtq5crFka6yzhhVpUxRvvxef6yxCxnwQSHie56UQAOg6Fsrnp
kr43QXQUpaoiIqt5++3lgefgKSSr2EdHDDC+XoWoDmswmO+OohhrcpOiik/6ElOz
vMo1uKhT5H6fJ8Ls+kXqklXR2OlLVbV7VjFXFZXJTWxDjBEwh7MvW1ZndCsR8iJf
pakhKslC4tpnV1aHpf58PnqL2lgyQi0MltRE6rF8DQ7FPwTPnqmA6Ybwg3C2dP1c
sI7fOphrIoyimYK3Q/jwVE4sFel/uSdZ2jjAip0n9dwxN7wXLz1ynZcM3EQg0eLr
3qNgeIe+ED9Qa1P+O3y4zK7UezIj8m0nSnayQdIsp+OCGZsUmcHlBdMDQ0/YEDm+
PSgUf8i0TRKbKkH74VhG6M6fHTLCopx6a7DlTZ451466/AWhx87vxtVJGEw4t/6D
6O7NOm0Ul/FHKfTPqagw9GFWwLpPyHWTFHjmAqXRdpf1AljUsPTanBQuIZ7JjfX7
XYf7sUd1U5JezoKkE6NiZHxckzdoS8lNeHad9syhWcBvHff1vEaXdgfAV445Y2Lr
QvUCla9BJiMDND4t52EumaneA5peaNbqNaYD5S63+bQmhVQ6W8UfVmzTfGyGCwA2
VjYhzUQlFqjVVDUL7vd3OjByVC/ntRXff8b+YjdCPiqo1RfseWulHr/yZp6YLk+P
lah3881JyRjHSzyV82Nx3JOp7hwJh3TpgFG2epRfrtPrXt3XK8tbw6bcNVSG+YKU
XF+7PozvscAo3yEEiDkO8V31OMddL2zBuKrWBFW9CHTP+d+fItb1RCfdy54qJsvs
NxnPvoksYiK/xJFlJ9jGIZD5OhNFB95VzEs71VlpGMHiNHJGBao00Bhaz+XlYyUb
5H/jylA55K96NpXkkjTeJ4P6xRY78qLmo5sC65HRO/1hi0mwt81pQiRL7Rqnq6Vl
LZNWBLZU20SctutBIWNxPmyyvRqNJvlHzZ5GZZFy2wWHgRIfse5GDt029IYyU9s6
gGF4lzz0fo7SIEs+BraBrhLsJzEISikAgLjArVfjqPXuvovlnqRfGgCQUVLpIOtp
Qoi59GfmRwMCWiarEjuc7cxg9W7UHF5QpYDFP7S4DX3x+KAOxUjpE2xsCbSr2Jm2
Y8lfhWv8S6JMx7wbS2AH3Hu0xtU4AMwZIhOb9+SGQK70QZvGlaFNGiioeSNgGcjD
fsaluVUYFDd93ZbEvmM1LGE1meFi3Tl5D1dyHAtix/23MfDYlvxzcmK8Q9fBUJDF
5YvvqmXVyVP+ml1YO2BGpjTlapBopZ6s9BWJTnW5S5CRtwMqtmQLwqHkvgWlKbi8
Gxn+n6m6+uncRf+pdrs6Qz0OKNZYsuUlC7ZiZzhsBjBuf4VQ9b28rZoDaI98HPSx
zWTp5IdcDlwmlZB7aCbw1Y9QIRgjhxNgcT3c7tXPPcwIz23MgC0a0580ctf2hKFk
k/D91ZFffxe6MQ0JK3r9t4YQV2XmZP/6IxxntP3+Vr0Hy5LBrifMVZi8CFTDevSy
2pqJEhXoCvYH2c06lNdDgbjaEF/nO+YJFxDyPn6J3qOtR14EYlaGal4yz33L/YRJ
zY1srvF2uStcFryijyIU9Ohf1edgUwyR5oXw9pZzi4zl70xqnIWQk7VJDHoA21Pd
a15SFYk0sp/OWvRLsGI6wjQ9FuS0PEcnvApZdqGO5UOJrLYywaHOVorkfLamC9da
M3lezCzEvH1RLdZDNAEa/IqryRxqkjMAK0VELawVYqU1ndRQOF3WtdjDtG+KQSF8
fl0asM3HaST50H4lQ72RFIx6ItRxL0CqO40NGHeBz++H1dwztckvBnqY5WxqegS7
xEnc438VSYgTs/8848rmxboifj8frOVB4hcegvJxlNWNqY2vxUeu+qgiDiCP6Gcl
aqk67RWYX4Cxlcu2/YoEdodi6Tm7w4rtu92Z1HptQMTZCuX1a8+17UVz892KDoA8
5Yl0hbOze2dkqmbmsmEOJqwl+36IZIa0P7HhFOaCDYzuVVjP6vjh203P+nVojr7O
yPuzB9lSmGqiE+wdUgvDF8glzueVQ6AZTYt71V70gjwtX17h2gf4xQC6kaTwug+N
Ajp7PY0x8LfgS1x2wwDkUNuiyBjrLHVMWx3DQPcXi+nNoq1LfdihMgHgpmWQ7BuT
M1zhLuYapoR+3E2m3Ruzp6CuhTZn9WmETWVQTrrNlh8xen7tQ6b8nCwwQdQ/ZNIW
+1LxCMv0xyzzwxCxfkxbAvbwiADpQ/pfgeCWf3g/AWs0E3s+2qJ1lQLG7Gn1y913
9Lj1zpJM7chTk0rnHDJ+1JGoEw7nMAmmGypRzxartv0GpPWCdh1o6F2su7v7S1pe
vSg+g6uprS3qBBTHkcLzhXiJX3C4/pyXk2L8d4MrVTGM8O/+o+1J5rx0lC/hcPdu
d7bpeCnBlElRZFvZO0R/Jhm3noSgxB9wF38MrFj/TzlDFlAYplDGNH6M/Qp5yqak
onpBQ1ilk8xnzqqzcTgBOYd6F9zkVo1EaGs55r2kNaz3PWl2hYSd5jRvaMrdpJgq
mcUY69i8dSvkhr6VyaWeFtaT7tmNtpRrWws3GwW+EiLM9xugoyjoKKh6pApEQzja
Elduo5GQQDNMCZgB+k4sgi1+79vPCh1DS9KAU0Vyeegu7DQOGebZzluspnBsBilm
YhuSgrF8D1mr5Bl7eITG5qeOvzyEcImg3lXZloz6hABYmYZoGKNKymaMiiRVIdBN
9gQ7rBKtEt2/E8raQfCGG8aQM70n+pAhaYAXKUjXcSspUtOM3VNIFw05oykx9G15
dEen1ZVTofGMpLWlRP5RtdnP7lGj/36dyWDSi7KuKowzQ4T8eNvghrG/MUZA2/bC
+AdcFR3RiNFKhg2D7sMoLo0q0xL0SKDCyPX2TID2c8j980oOAaCUvmEKn7pMiRh3
4MDVaR4uS5e8u2kw4I7AV0Arv+uSWrQ9pI41JfZ+RiYxa55xxXRfw9d9DFCe2qv8
efFZ/EepL5K4a5q9ONpsktHDoy8l6znXKi1NcSg5MJG+rcjzEX2t4xYnF2K14HGC
qjj5URnQyJOSP5tVZ7EHlJBcgvgg9dKJg0iEop3s7fukuY7KxkEq2bIiqQsohXHV
38gVravvMDPJvk7JnVLfqa1oXqmtJAoFRGg3IWjbGmJaZhHwEYvJUtAJafzxmEHv
aDKDKB8Snb5nrtXkqQXj+TJHxg7b993q8d0LcYFWUMaxAhS8ZSSKbXmXanNrD9Ip
MpfbFX+CisFWOPcxj7RZ3byOhn/UQ1SyZDuTPaBFZ7HFdLSdCifC59CF/uqQPsvr
ot83DDEh2vOSapOJQQ2t9tKwto6uynIeKEGG0javta7zcVuAnDTvJm0S+jYZ4CnH
L8sIT0eDcXhlP9YuM25I91iTDNGTx+h86QGAdU2dmejC6TDWrKlap86asY5qESLy
rHcIUM/4zv4awq7tFd4OSn807BS2Iku2T9g6jdkc0zQ2wrOnjyNKGLTAJ1OJUNjn
RQwSXVgOH+SaCkbERqENk+EgHh3Kkp0mjaUHrzc4g92+rSbAFEET/1m0Rjdj2wmx
isNP/x3ymb5iPuHdkBi2HPnFYNkQlejvSOs143Og2/yNwZAhuObDkuFDejMIe7qA
ipLxd+w3YOv2YtZx6vhY1VlcNu1AXL8dd6CAJKrloFaquN815Et37Onwy4wZ9Utd
Gg0HJMvoxNhu39AqEgpx6/IfKEJHyQ0r/GEyZXCjnKdyBuxmUNbq8j3e0VBxugiH
LNL/1N+u1Bv1Q1SHDkQldEcLXZQY92lRNdbvHzLqrG+uIPBi1qqbqPLIfu/BZAgL
hPOTwtgfeNFp7kc9YdVjV7ygX/eWm4eGrwlYm0yKuNugjQ11oOaqvrmQl77XSlIW
MEn+fcpJM9KdiSf6hqPrrZVPdCNusBI3f9CNhK3aPCFtwHsHe2nTENFQqOpxwOSn
pjJZE7Rj6iw/hjfnQuLDONyFL57v+PoOnrkXJ92/MzwWxnGWNvlAeavek2FKO6oA
WOLVUUsNUzx7tIyJH4S1sRrNncyxlELzQF8p002zmSq0TseNPjk65J1t41MjcPit
8niOgCrhtz8VyPmfCxTTDPakEnvWYVfH9sGxBMQ4Am831Hg9inRpP0003CVx4D/T
FgxdgkxwODvT9Ljg03zPszjlyxb8G5ctfE4ILJvajkc6iAHwyniPFiCTWGItM282
ksoAhhuvrPUhbHB9J3rgdzms6q6ATJQgSJAJ6d/8VlLpChzklZbfNDPt580UiiPi
zOUWYPpnn1dIF7PuL6LMAd7ZlMeF7t/4AaJsODxaVbZRitBDm/Eo1qWm9VDyXg6f
l7UYvHs+6j47EFofmV/Kk3N6lmNH7EAR61PPqNC66m1qlRTunxKdz4WyfThK4dY3
5NcL+qR+VCMwL32DKYUQcW7lr5Odr5Zn9M/4w4A/mzWL51o/bacQqf+4PmCG2xqa
TJiyC2dPqtzBfmtujPOURFZPQbt/KaFdpjVm8jCkuE5O2SYDu4Zdu+BK2XiYnI/I
Z1Et1FwuvL7M+PV7fXrm80wozNdHbnp1jsurVF5aV6vDz6SC7bMYubc7AL43axNn
t4MJjXiJWUFNdwXwRpTELOQIt4+fWi+cVZkiP/vqPLv14WBfzJC/zQeWHK1EE4H6
wfKM7Sb53l/dS4GCd8mRXu3fztgIVWONwXHRRnxTf1Xemw6xSrKMdp8Zoi0qU2vs
AK6r47v/rMfL3Plz+M7HzCQ6Xb8KeZQNBFUYwvG6ofahT16RDnPhWFZNorWFDCVJ
9dJ6aYbJos37459firda+6im6bDQLaNguFhd2PB+UXBMhmQjHWi+k2SzN5RdxrL+
QG6p7k01fMOo8EbC8dw2PNspSbNy0G6qLnGd7nRrgiDBgCehsP67iv9MsOWNz8DU
MH9rWPVeMVzrUpDrYwVg64NowohtVhv0eaCPrOhoddmny8GqFFVa//0HUWjmHGrk
7f6CIYg/4M+ocgsFhNIoV1uyiDVwtFlSCvwHufGTHjR6S4RPjmtlhtI0nzJnTge3
cWfw1GmVrTSw5A6F3TynQFbRhLxKAU5gj5wy9o9yzRZ7Ax6cQ7bAswiJV0DxIU9O
USQs7zBF9/hhJQ4TDD3s3lO/0DjH3t+znIHAkChwFbR9wuWzDS4RWc/JrY8Sw3AO
TDif3WxJL6ESZWKUsAIf3Ge8ruXyKD4r8EbcHCnOFEzbQrWtFzX1CTjq9LUu0QTc
vJD/5jij/90hb2B77QO/AFHRYuTuU2TWzw33agrjcIGYmlXUdnDgnVPgcSlTxCgy
+gj34NSwXz5KjmtBEI6s+xhK/UBsPy9Nl1rldaBOc4b4Il1wq2J1GLZRF4qMnOQ4
oX7GjOOiLzM08EmxA67l3q18pkqljoULWQb/7cl21cvk+ZOM3KCE1MY1Va3h3T7L
4GlJrit9m0tqWsjAj5fjR9Dk68h0WkckrH1Yr6jDhC/O+/u14rtQn2UZh97lB5ED
Yh2edClog1PvYJjiXPkZmYXwt4KCgFKWJ46n6zu+VBHIOALuZnz4SzVFykpGsZlS
bfiYIeMgGOW4xnb4EjNRhcMjTZXAQMKhTDFkSold3EbcDYamnfCJC5A86sCK7hck
bNGOUOQqqbJinTJHHh0imw0mOCJccykYoX7O+T2Ku/Ug+Fx7L6jgSOHP1ko21EPR
PWOQWouF0Dz+qOlMEXpsZeAf1PqqYsSlpq6iltwDUsV1jSkXJjw8ouL3B4CHkMDl
G3GG8ID02TrVOuhzygXBK1vNHfV/Qx40skKCvKlNfsO5rbgmm64l5luCl/APmQ+A
OAp6a+795hNIRnrApplTewhsugM+2SR5inDR7UjTI3xMAi/xZTiYaNFuq9y99NYh
NhYFDiMliaBeCxeTLMidGE1JsBXxwTH6ANFa8/cQsYgc3zuTmIBA6lZrx0Vc6OJc
RNQq1SPcep9a/1TWuaFf9rK8mOdToNHp3TX6jyjdpubS+SwsB7N9P8rGMnXHV1Ti
eBzvwEzTY+XuwhaksRUIU5MNLIpseWohhUvVPc3GUkv+dCnKqcytlqCj3rdi543h
/BCmEIcOCJkwasQCiw8d1TNmUoFCKYqCvpD9F9OUlVxdLuPUI7f/NW3tmnN6zpHu
0p4GOSMOZ5JvBrnKUX7Ou29I02rpflFQ1jdfg+y/yxR1TAoKYY/1XdUorgJ3ynP4
3zGUHVCFo6Y92E+VdghNiVc6zzG+FqlzLKwOSOI62qKzmGm5LvjyQ4WPTpKNGwDA
WzJeqYp21VRY/eOKARHmqoVUwBL2LmueqJVAyw9a4hTa/wY3ayksDdsOQZfOPN3p
zux6wBaAGRQiCALf0k/Tn/6LU83LS9Alr7UIOvHDKHaM1By5CQRJigbyVtkWnK2J
14dQ+65Rbfp5RU2qFEzLhxU9YKMSkI7vJZW95FhEBE5U/0uj30p2GjfZ9KKVANqi
HiuFxiDGD9Wz+6t0rt4UqI/TL9mzUkhbx9X89sM7Bok8vPRFU84MD8OSdX4XekwO
TKkaUSeWb4Lon5BQnjjgSclbjRxVCTiT/IlhAjfYXX2soNKH05wY6hV0215yTpjj
QsR8jyxPe3uGGKxgEp4hwI+wMK3Ec69fTGLpaqumR88/thMY1E8d1W54s1mICSKA
x/fJw/T60x+x9oZ0IhB7qJMqVkHiyX3dsvByPoBZ1+7pOpb9cIJ2V1ZuoyJS83fc
boqeVSFozDXb2uD76q6Yv6VCXpMSi5jBL70xZHCKeivD+T/O0FKKBwv8MXRmRaNL
BSdFdtCKaOCRm8GGFFiiAZzPoJBDURfVanqM+e7jCnUDAORrWqAYZuLKlECBno/N
6/zvtMww963gZ/ybxPlBpwfVXDXSSKvOKKrYT7SKA/BVdYhaCe64MGzQ+KZlN16Z
/WWMIKwQ/c88DDkGo8y1AQ85ke6ACCmuGqKT+OkE6Xn5yC8x9eNeecdmUG7VEm86
y0kOXNPqMTBiyLFIf0D/UDAX3vsv6GxjPrGqZm8iTUHFdduLuo7HDNcWXRpRKTEA
LzdU8Z7JtPbnegq9rJdnZo1XVyeMhx3h2w19KA6ajvJLnlyVslD/d0bid1WlIgZ1
ejKfLCycyGipE7UkUra4d1n/WWdJDzi0a+3hr2+OhrgmnBAcNoG9WhHRe695RVGS
rnrQeCW3hqdSYmNVnzXZGlButWJ6OqaATNCw+SQ+M9rcREkPmDi5BjTbheTLV8H6
Sp8gjpsHNg/GOOjB60Sxfjz1OWqvup6twn4bqVkl46ZYAXCnYEmf2797lvKiu22k
k15riF8BYxtaO/L1BsIhAFJvuNEELASjFtIkm2ctQm3//SDnud2cXSBcOmrLjQta
wEYA51tcu4hLsa2WTboTywUFrbo5IS9lHf2E2D+2pOgGeR4U4YF3cZA8uEX63chR
2k151c+xtNJEruRjjqXeS41S2gtooyewxzAM98FOwsP0qisPyTKS8JBlJWBrQgNU
NP9j4OGywWQdfQn+r/uqQlemXS7MT/OV7EQLXAFTFaME2JLzjbNwQl9/jAr1rbwP
mRf/W8JmWEMbES33Y/d4idjxkDHNjPqF/f+OW+YyyLcJ8pKshfr/dTma6r25CUZi
tmWm3oOF/XFElICkGRSdVwNIYPTEXf92Q5a8fbrifmngi7OJtHfOdoF4tcTrWTEA
JjM4pOxpABYDNd7Hg4YuUU+c2y5ghM8rpvuEc/m7uuZdI3d16ESKApQ0FtYBvi5/
8dH1BOzhjo6jLn/Citcp8JK1bHJ1UmCjpjhWcqddZyiXlHxCxpNFRz5Slccjjxx8
reBtS5DI3RthF48+l9A+9X9jNOX6qsOfvL9P1B6XsrUTn0KevGmGX5f2VPaaXgPX
xD3iEPUCzO9bbqfHsisooIGkd3Oig8cLkQjMiaZv444XSGyIHOlMYKmsGYOxUMln
pOXQ+0XwH+6VshxBwpAfetebAadfc3YvBz+qW2kX3MXV8C1H3PCMSNcGVirzzeS9
kdVqQbmP8C47ISd5JzIN9yTxPCea+ovRn/Cx45J+hLFnptDbvTEvIQ4tZn9rx2oN
TSTsXO6udkBc8VUaJ6VFdh3YVbDiWvY4BKyFgwi7ktS2L9ARz2IdB1CWX91F4ABO
iIkSM4HMjboqMUCP+3onk+tZyHhVTrMjsSaYUfnWfkO+3ZlpOBs7wfPs+JI3gPPT
Ur2blZnF6GT+5YxY4rwjN/JlCSINR6FOBMegFLyalykX+9D3OT4B6UQ3BOjgtWj2
9I+UbCxJFuE0d6fReGEupy6Otn5Zlgpo2bBLJl0fcGp3HAcAg7dMUvXxC2AlWs2M
dCa/gy8rtdAOUjCaLibcmpbPe73ODRPPdDSHLdgodPLqrHkbVoIg/9ZnBGKzyvtd
0LcldXzKaoyU1uKpI9eSENTrCUVP7Icrtfu9yd2YivdUKE3ansIIFEesd75TDnAp
bXw7jsaGOI1ddTJd9LDHgcPaJHZ1GcX4YvYdK8POaz+uWLgMn9B6hsk7/6K/yRq1
AdRfHOV+tZgaH6ExxFa1cQ+xgA+lUiueOtt9jzsW1+9n5/uYkQ7Ltnkm0sQsHkQW
4QZStJvRj+ID3k1RqvnEshY6E9AWvx2u8kJ64XB6e9WGLMfCj6iDymzEVRY2NP/Q
4ldaTOPegf2ewgT2NZBNcVQ/NlgvEelUQ66X4rFef4AjzjE2gCNiZqNNQReKiR+l
qxU4y61UYTEtJxHAz4gByeraVZfbF8iAyKtM9mQmvQvjh527k1t2MGrWkQ+0yZkC
z7envZ9GFB6f/fplN3MklReQ59okwnsuoYBk9ecQMtOGZma8+1Oogl716fZu3DVq
cjvGrinopbLGXzc366uIfdT3eMgb0mWb9fG2iIoeX5ZU8XKt6L+POzZn9k5JMkdL
Co+FjSER+k3tjMai14XJJqjG+ZUQ3PXm6VIM0VIpGmdkxWNcyugB7czGqwvtMM3t
naWb6r2leq8Z2MAR09dvzftRtMb8AtiedgAIT42sHmONUd9mVlmqn4qfjH9U2iSw
Mycj4nWjARCty1daM28FZAC6nqKr1lK6urkj5AFVV8KdmqfV9DWleLUUa87566kV
/OfPDdGNQOIB28w4SI7cYyq8JDJhfRDLBOADkcgJUMd7g0ylJvIrjffm0U4JO74G
m+6av1L2DZhclx4AmgrQhtMRkczDDrDsdUjdMI+dFtAQ0vzHgje4bDqZ8Xsa/1Ys
/ik1MHZVfP/fy5Gw+IvasZiWTLwo12pIJxlHb0SJzxtuUZ/7A4g5oIHU9WKGvGhZ
5uHy3ZqXvlWzgaH+dsHEcIDUywYCyIOv31wRX3PkM/eWdZXXk8UPpjYldt1d++WI
3mdHY1APzNypcMw/ZlcNOpJA6KGBrXizNjULfuUtYxYGnz2FidHckRTVwNW5wJDQ
fxqWORL56UJUMmJPvjFnDqI9K/+a7v3uBsDSiZr61FW9KRza7LyM2ds5V2fUglKQ
fUYsoOahSPTYtWLAvcbbCn2sb3+I6kvE0X4cb6fUdm8jvbUzCHdaXGnBF2vlXl0j
ZYe0DuKY6GOQgx8/PyB8N1eKw57CbbsJTqYvrGLw/bAJ2b86T5Wuq9zW1EXSu/qO
4EYIDFhN83xyhpnRvlnrdOyHpqbAphk5PbZOGJ2xVVGTkz1X0/oSHvM4jJoQ/iH+
oD9ZsU8CwA6nA6qJuzYK5K38DdXTjRIM/oOXsi+P8E0C/us6s0eMKmgwxG6Omry3
7tKJFh2Gli89D74tiF2LRkPYEvPOpStd7Xt6qTRpTP2ruNopOKNHGWDdm/nQGPDj
M/BE4k4/0jmhLxOJduM1g05TYiV84pFPZ5szsWIa4YUmfH4S3JmtUws8a8ExLg9c
TJMNvAWIR6d5qBr1ggAPlGdPfum6g15HOO463BJGnh7tsQAk3jSQo7gsEDLV4SAx
2NOa9oCuwMA0KOFa8VeAOjdw/CTOeF2/G6EHp7B8ZqVGage3OEed+gMwF8rtwCo8
jT1KDQi/KEbau7/KnKNP5rL0/daRhgGf4n4BpwPs4cO9Fnt44CvZOyuxpxc04MCY
GlSnACjxYax9IPy7e16mvnY9sX4Ei9eDxen/Q4RVFkEswbPyr7syKTmoCkOHeDwe
C/AIY1EprSegPZbXoYjK0bD8BLKdVBMeVQA+6g/EdGOtjdxmuQ2Kesw3lqHJCdtQ
3hpUMSlFNyRzviE6Wl4j9ecpLYOeBF3RFJwGYdjkMX0Crtoj4alf3nH4+97gEhxW
CXa0SeLaL8/LafIR8lLihTJ6ARETjPsgJKc5NGl7Hdns+TrFgtEmM6xMuiEoi6GO
dGXUQahCYAa5dUlkITUUTIUkD9xpqcimTTEr3/RKm5+MRfaEbE9vjXYHMHwlhRJa
4aXg4eCp2l8dfaTPL3Le68IdxnNGLzW6awg1tcCnB779/+eQax6iQQIykxB0tdCH
QPCx/0dFiXUDilQGPMpqrN6s3IvjocZmf7AYBFR5a0cU0VAMfq1eo8uhaTm0SVaI
Zy4zKfCBHgCg6GmChsqy966hLS2pzpqHpLQQjpTdsGmzzVFRAcmaIQAE83I04+ui
vBohJm9xBpVbG56t4kVCfrbCsmOphMtLM76B5iw6jBi/gaEk/YVwJwov9t0ctPxY
po3gDIYasF+uZJRob1in0jXMCvg9ImP4y3mnBT0G+aLP9PB2kvx2PRAAPyLe+Kfn
PJWVuCr41hGB+tplUmMqzhCbrvgttt6kdDkjzsDT6oIqD0rJ8DAar3em55PMemYj
rCwTHF6q54jEujcR4/7BAjZM6Ynm5EYv2pVlzyBvPKHaRlkstINMIu274J5nGfVH
+HjV1KGQlupVG+PuS+g81o5X9Wz263GshMUqOxpzcuxECrwYUfjkg7hG3r3ezrBB
m8JIX1y2avNPPPt1RS3flUfospIPysiHI0AagYC6idb4Ijb+cJurtJ/sXHK64m9A
Q9RbYQ5p74TXlMsM8bfnW8kMEQK1sfS/rPdjXeT4Oyq0Pl3dUSX/w4FP/bJMZP66
MdeMVOCmDTNW2hMCUzy1aJXMzHEHhTIP7QZSupm3UYRx9+UOkxjsDZqFc7lGBEO2
jp0JtyunJekdHpowjeSKNJTLeruQX3kRY8rdP15BoAUQk+2RE6mSI52Y9RCtYci6
x6cQ39yUB+TOvnG2G07eiuJNnkwdoAfR6GsVxNQz5RyG+22+ZdcCx4AVIH6B1LkB
cP8GnvimOWSDkYNQqhwuobcarALbagGOLL8f4dtc+JZsDNMOdeAgVLQ3ePTrXBy/
6EkoaGW/XdU1gTNjABYYorQSl56+Q+8Us7Zw2UX+wNarIm/wQxKVIaRZNxoPN0Kd
FHsWJsJhO2blD0YHYE74PvbS7UWlXPpIXTqQlhabGlARWa2QQ53Ezf8/8GFlMM5O
PXLr/xYWOxvKhiDXCF/WcJ9MhosAZnwY1z9JhteRMT3lx74mr19JgMmtLjQ6jTt4
B5p9fDgGMM/o5l6xM/zv1Ka1YDzCqtD6IjpNtdefj3J/KWXnNF5Koq5kIpG4Qy7A
jhRfKypyH7fo3krEO11DVD7IM1J1qSnUcHdhuOyCzz9azHfIBNHE2v85J9OOZdar
nky//ozf5SFd/pMI2PZ3t5d+zmlnRKFMqtjV8MWf4/B3GEX/OGLez9X+ASYwUcj2
pTyl7iqGGO/3kecJhqq+5AGHlE+GcIg2p4tygBxC7FIpl7Y3jbEP6COXRZfljRoI
uaY+2pToxjEGMu1nMB5VSDY9m71GHu3BGpsZvGMQF7AyNhc9oYkKDXCqmULtPF1j
p3picqYi8R15J3mlrZfr6mGpCh65WVkW0IdIrLemAvnpRk9A1uaaxEBWGHb/HdBk
f70Xm1g81uy/aDZwMQapEhEQFomu/Sat/QwHaVXGQhZzv9YVnSosRp2Ds7BmOhM5
t1WskHu5bO8RHlEfhLlBJjipiQuo7Uifjh31mPKeSX3w0MWLxfcneAU+SIBh0vuU
nqn9DOIPgVwpN9oELqqoguKFZbMhAmvnff8R+XtG/LEGCipR7QwPDULRtBKPansA
N2Z4iphdDKooUouvz8tHOIE8F2XZ7w6Q1utw83KMU4xZBbmM31nHy1TfwDK+18lC
eNgR3yFcm8mDzoMWNpBYfFmaAlp+TryEM+FBzVl42j5UBVnoszxMpc6ttplTMadh
9KtwJp/ye7aA9SN4DhXiXRh+t6XORKegmVQR5Sx9fz266Ul+VdPQdSFh7tqGveoL
9+9RduQg9xWrh9Pk+CuGrhCmJBrLFrsmv5Z9NclfGVrLe1RFiH2Tlq3l8BhmDRID
W3phF50x7LYraQ4kntELvS17SpasKufZdMBKl7Drx8TxeVj9Ur+9wEK1OUfS1wns
sieLCqVqplR+rplrP8645CwxvkiYoXq0/BJAgfxn3X6bKUVUQchBuupipqJ1t36f
tihFUeU2fXMrPeESAFJ0R3TnEbKEYP1aCIIbcqZBjTdxqWS2SRtlRZwNwbgz8was
ztq0whyz1FpIXnGx6tgNoW2ifOtd+BLRHtUF2O3a4TXZk5qMsO26Qjnxp5F8amLq
XNZpUoWPBA3Il91HTUollmU3bqsJDlQeIqeaESe+k2Rj7LXHT0E+qUfF0q1PqGAc
Kqnbn80GcVet0NJuCHMzR6/ky3tj7Io3vHFto48cHSaisvBA5BXlzO5Q/nXwf2P7
3oTUDDy6OsZD9fzyll3M1V8ltL+sdBKrbAv1fP8e31ff19BY+6DiKh7F93di9DVq
wgWSwaFGXjg0OTBhh7eNJsJ0RmLGhpFaGh5O8ImpFupSWupF0q8tzFrLHnuPyx3B
QfDVCEk24O2yMG0DsIFDDmAI26Aj3JVNvxh9mTZsnHrpcX611qGcUyDSBBd1ciGo
8RuUxYZ+XLv+rwZsyMoV+Ln+ew+bGUoGGbHahYLKswZYRDgDtAUjZ7GTBJZt3ZYv
xVvsRB9Lscw5qCu23vm8eRFq9eX51wGPwdBQi3WudA6oXwzyS+oBsEi6xPGQgucb
x+t/V0x9taV/pGSCbERxyM8rvrVax0+w8T3YDng+5o0Tv/VkfqfP74goAwoijZyf
RekhuZKzyq1XF9yDTmd4e/mmElt09jWJ7l0wkjf7tP/AeZx3itoP+rzp3MeRTrs+
KoPV3CELIZiVTzDXZ5cVLTuZCd20RwZBPMjqN+5ZrVaJH4Fjl30p3JTGOIItwKDR
Ze2hnSkMtSv3BZ05rG7os1/BaEDVJ9c4xHmDRpRUTbf9+y7jM0ssooib20KxXX6O
IH4aRgwvLeydzU/ixN7t9qRfmsBhIMQxPiwX5tEuivzAmIbz/dZHPeZf+9dQaQQN
HDJ9sx0nnOJNHkcb4LNGdsNmi+42syBEK9+oUpmM2Xl+Ul5j0z5h7zKXL9I1JIq2
QThJrOH/kiBB2W6juzYbrgZJA5A20dnWSrj4p4d1BJe7oBlkvjd/NpIoXKEWrvUA
/Q9xy4oyrDGkQq+lhg6jgUe9oDipCiqTmNiaqOVwo+ecOTf4CoFYAhKe9sHg1zdr
IzYLf/z3VMzf9rue3NkeLYLXz5yXpaOEa7GCWwVPTwoG8ZNIG0NZSZmVjC4WHDXz
ngIZu1RDzBEW6sYP3AjiAHN7sVIxln03Hw55Jn7eX5dPfDZFIjwO4GqFzjmcoqqK
kj/IFt8KBper8ts5MUyP0WkvBnu1rWqVQWjADLahCboph31rb+8UZUIuXH3BN3cD
fdYdo/LI8QNGKZ9haJjI088ViP74WMHk8suhAlSNwJ0yK3tN10mRT13hoAOQXk/J
1NIIqaTELYvdToe2UHwLVOM44tCGzsGqq4IHRtL1TwgVLER74WUntF5QdUuFEsre
HUMA67K4zZIKW4fUbDpROkzSHCUKRG/Fgsesr/sDV0EMnML8/2FEsNQ7b0+7hxUg
E4iV5zjzddKsWX+rnMFnWBne0OqMIutoTc88io2+N0385Sdz5Y1LifZG2BDjX0fK
UEsKS75bRPL4gprfm7PAc9hREc/vX8xS5eQ9qBwldgeV/9FdbWT4yGSl9JOlfYAz
9m5HywyKWcWOxphV6YWrtzoXkPzmQyEz6Rf8ZglRtv8UnKV8yMTrtK+5IDuOVBpt
/EyeBJRQ6Ys4TVs1ioOhQhJqP5/uD+q13lQSYFkM3Y91QtlQVZIxuqJfvpn2W2kI
+//iIzn3wbAR7INKgL7MNqjHh/GJFDTPKdpALQWLekO0+rnVtgdWgNhXIOl7Lxj/
zfoqzHkTMAXgD9n3Mhl8+ZkgXBTeJZmf7OGVFpqVOPEuq/rBTSSgeryXSOR2OJfR
v8iy8/IfgjrJZOTm9bMD/EczOMUjmKjwKl/mlCCpBKOg7jNH3MV1jvdD+cHpDD42
JmKNS32Y211VamvCRMJfHO1Ek3VOGdU0h3Zc6494tpnEgZ8Mdru5lL/a8DvUTqQ4
r8lrtvm20uQ4sKozpMYKNHaJCSj5F0blZvj3L2G3zNqAb7ADKxWW20a68Q+EPQ8K
+EIAvwm5PvmDjz7vr6o/CW6o1eGiGaZoA6TP6kGNN1X/m3pWJgP9Eq7nP7xVSiMy
TFd0EmAQCWLjwWIxHx+gmR+/FUl5QGSU7uDUeyuupkjOMtQjQ5648hYOuXDJvwve
cQi00uk+fj2RFYVP8u1oKFCB+SBpRog+BKxZ4I3CecNVqqPnkhLdLheLp6GPInE/
NJGAktJ+2HoAu7Z1ynVJWIjpIkQ0XyE/7U00gvwGd2InUfudRMvH1Tsvf7Im/9hm
8G6MlNqRo9Q54MueB0fIqZBKbXo+vmlXcOhS2kNnRScTn3u0c/0dP1C4DbI5IUkf
5Iy8vdUGxuRE5OGo2qdxUg3QeJel1SMexANjUsQ+mUUofwsdAeLnk0sCoz9YcVMp
lmEPGghE0gQ4b7dnIarTDhw7ynPTJ9scUlluD/p37NBUIlO0Fp3P9uT5w/G4B+10
oiCg8/htvW6ybFeWZebAGqPyhgv924o0ReDz+vzA2sDQPkQiytOqsRByMm9KXiLs
TJYjC2yEQCTOkr2awJ72M3L0i1IwBS/vc4X6ZaKiJngoxxk6YrmKVvNIsa9D2n/Q
MUb8XANB9kzbYr+PYHhXMx5GPXdTKHDWu2rx9WWkAWEQNQs5kG3W7Z5ZENMDpY/0
QYyi6Ho0rVo1ytx5C4voOO9IgwF6oisN+51yuTgwWIJ1YntKNBDa1l2iJLlC1qUs
kOWDZAjtFCA3C4bNg0+J6bPm6Tyl29d60qHC8fv2mnMK8n0H0xFBkmZ8a3pOY92O
T6zJpb03tSp5ytC0ZDfsSzFGM5EJYsJYWOcUk0UADR1mYQvLNjXsrVLdVKwyrGnP
wcGSShaC3XQ5ousSyk4nHz9A1t/ZTQn42sfpwvMwhQWtRpiSuyoKToqCI3FMj8Kz
Oeo+UxnnIoKvkdOJIRMLdsLG5X9NyZPmJoD3etRT8LWGLFFk6YfituavU4ydc0XA
ii2tE8Hamm6mIDZjHfLueRCiOLFASyVgQHFbqjy2srNrAPMGmWRlS2sZ6cHosY7q
IoeiUXVf2W5UAlHFjHI5Vod8WwDKzVqFrtITQHoeVQkqFGqMJKcOvBprxh06uEdR
dR9AbSNV003ED2PXq4F8xdx+PyD1KAxK2sMX94FXxUN3V6k8W+lotRivbPKNBQqf
g/CxMmEeKkArdhPRx7dp+B7DpggRRKVbSMPu+Jkd/lD8Wb6Tsaj6bbrB0L38ZP8U
5jLrePNHpCLy89gQtgmo4JTOXxU1r3H2YzSmx/nqPU96EPqY1eCYbzDkWwgqB+na
wgjm68VGdWiKMnbtfsUtaDa8B/WwF4eY+b6ubvoN6Cj/ZS5RZ93RT85wN3QEF8sn
7OgIA96DBY9mhygB47gUk8s1LOECEdvKHzAn4+4xZuOd04Q6msO1JX38k/gIlZ0I
k/2lPIF1G8+ORSEDysJTi+hK/H9sNOBGxUKCi9sL7uNKzM9ZHE6shkED2VjQK9xn
/0bQ1cRiHA3YQk/CdgijAg3h3PmuvPa24ErQXHappKHfEFVMT12d9grI9V1m48eX
Ix/yiCnmDz1nYgtkU3U05cD8AZlFgd40fxh+J+ayDB4S+nLbZLGBi2TBKjoXcLzz
gLe7dK1fwDFjjc5IcEC8/1hIeigc6lQA7Fn/AQNSeZYZAgBSI+nZDCQOeJvfk0yY
GGKZQYqyopLn0uhvVtlIWzL0KCcO3LpdfrVXwU+sogkraq4JfC2ltNb6M3FErZG4
+NdG18EEVWdqeabE7fdzDVSGgMCxxSCQbXroGRB9BlaD0KHDp3iWnRH0X3NKZfMW
JMgMhXFVYp0UYL82xKkZ7fEQM3xugUfde6r17VUiel6MG5pIapUEs5DWM2IjyP1r
CZfgB/3ufg6VTaX2kVxa1RQaQwjbO4+7DGRz4eN+qIuJ74h+cnXEH1adM4YWmxs/
W7H436w3SPfVopMhjd4aMepXtho4gNoHKMUmQko4FiHtYEMHYKfu/W5E4opPyauU
/AmnLE9v9wC3y3tpQnzK0lvzjj5R9+3yexvjDmOht6z4Q9b33Bf4nGG0k/y1N6Cp
4pUuAc0Bbm4AG26yVsQKrDgssEgtmCT+DMDx1B01OYZnw1QJGa138AgmLm0ts5Kj
5TWvpIAwz2oHuKqRX+ZZ9mYGzJadxUEnLZQEBxfpgQ1QjjULxAHp8ZKlxbAIQPbX
NLCnZ9Rs83Ppoai2wNeagQTZMeRnHB5vXrZlEetrw9Q33em8HmRLNyyWkMwC+PGc
XtNe66W1Oum+75pz1+WN7kvhaZ24xAYWJQFkubDMZ+YfIvVsIZVIZnWdK96Tzutg
swZz9tHctm3KP+I+9hpRCdqaUhDPFwuZbRgHhxuO4MurDBozWS3R6Kn8fvo4Hnfd
Yae5peY6txovOwTjrV60Ph2rSMUVOiFTeb6VHzFk+CD/nvOKuAy1GkQToPgTh6Rq
A8Mwc7voOFaCHC2is/mdA1M3j4L6otHFVsX2Dn24AHVLeXrLcyx2d/+LGbjqmi7U
Pr5mTpXAgl+MGV0P3f0+r6Jt+4hC+Z/6zRkdJ1ZqDV93B0Ed42kyIQ42Zcd5Hgxt
laGIcdBHIYdubR1VIUgx1TIRziHZM2OTNfsGx62dj+OunqRDnmFBzMj2iSX1bQly
p2PAwwQ+XgIeSJIMCpMk3pz8+EjddJyH0P8EhowGl73b000hTSQsgg9do2TCBBey
YiEHbduJV5S7oXXtkQe3faAG5zCyT5oC+eiB8vREL6ocItDbL4KcrrhRuv8/Bxlf
MjgCAnmrE7+pe7vwd1PkMMbHvtsPwvqHoAktAmb6L7kT0nmg5dBnc5GSUfu1d1wp
el9ehlAAslhgIMe3svoCxzyoQE1XpujMZ4QGtP7nQJVV60zih4UAxf65hdHxEFcZ
MXbtTx5/Nyv/Lpzv/dWt/sK8iJoOgI21r7RQLrfHBBX5fs+h3N8y7+HRL7ycTkW2
GxL3ksosCuAR+sUAX2WdrKqUtC45UAbcsBsC1c2gBflQ8g3tJdAJcJe2wGQF/u02
298ScI6ddymMGZYXqoyDuUJdaACXq1fb3evMrNLknVyYpssEQT55nS2g9R4QQaaV
bEOpw5cjRY6MLs8nqhxcKwrXnV5Dc1HQykH2DXlysBHONBEndQVEpISpgGkWbaed
Pm19n2ra5YwWRD8E+x7srNk9tbaz4NvZ5TNXdNvX+dgK5lUZunDH6L+y/D+W92uF
ENCv8V7wClWIil2asOh8dO/nXCo0qIVWsNs4vVxKzJ7xK2nUes8NMYodVt4GmPeo
l1sAgN2wLVaim+zqaP8QK69z6YHM7tX/5xueKlVc7blBigLDbQHM4tUDpa4g/FOb
8HlbA0dH+VyX2JjRE9//Ac2HTh9tcQ54wDL0k2SURE4RKcmWbhQY544A5XAL7MPY
ncDsOChPDHyRo+k3YyT2a1g5m5igitJi1RPaz5hCYo5OPslbGs4wjRW1HWfJnQUk
TIbh2esT4AFyOri9Y8y5ox2oRed15fjvHSVxbN9YprVz5wzHmt4zSsrMTKuw2r5d
+QItm3oddMp4AlDdBY5cSTrdXfGB4cioJUrms/VSDXPoW5xPS1kRK+adEk+XTle0
eX2TrXX53SZlx/2de2lftZPAnp8QMKtsD6Yzsi5DNGZ1B9cAMi4kq4DmPfOP8fQH
Vao4krqDz70P9dlFsSTdS8WEyMbcFbO9hF2P8wOwvIPjJGFl93uOeowqizD44/C6
DxeAIjiEd8rG1fJ8dZL9QYiAiY3xmMgfQJhySYcEHKSw7J+v1x0oir+W9aZHHMIc
TS8Tfq5acs+1TSf4Q0G/IXPgnyy1dwIgL8EJK+ASG71qASzOJQ4VZ5KEwENQbTfd
e4sHzPHjWtx4AFBsY4Mz6O54go/yeBYeqVpQ1sXK/eqPq9tZnO4ppBdvDNEM3tE1
3kDD4wGAHVPkPaCK3h+c8Zy8htKFD+qjLd2ZFvaf6CPvL6i/f1/GwT5SOjX3V3Cm
uwEk+vpPVK/jes5hoD9N7mj94xsFQDnm9YO0xh0N66es1yYJeqYecUVSQ9nu7Vuf
/ocOlK1Od2VhIzAqaVYOE3jzcx8F8PJlX8EBCSPzoAQ1VOAuRQhe1lYsPvoT2/JW
ZjUwRdAJKs4l0k1tSJrfQyhqDq5L3iTsbF/bbZ8cp5y/FEojYFaY/YaZ9C4Hy5al
+QOw+01s7Tb76pftozcED6zFdWoKouE/8yusHyfo6ld0I7fc2iu602iJWDWdcpui
p30t1EYXq1DLXelNZGj2Ky4j5cOmHAFqu8wfdSdpe1kHodxqmgjxpNBLuJ6lcL2K
g1IUwE4Bqo6qUWqgKdUt4XPUHQL6TTHLSdpKDKynQikZDcbtBAgqxHZSBDyJz0Ic
9GxY6rlArbc/Y+xs+4mvLFAkMKQ7O7Ib5mWv+O70B+KmU5ZqwdJjFPRQN2rfVPJq
/aBXA53r+v+F1MyqGfx9zp9BaAmdGICMNd94qE1xBYjMimLNxer7Fr/VkmLHXjVC
UYit4DkSRYejvipMvn1/sL2jOCak1aNg3ZRBNBRrvxv8Zi13yuzne/pUOH9C/Jmb
6aICkPMCeVA0gT6gjUgfK8TETqcn7XEtE4YvaQhGM1JzX++nEJBNwE3CyCOMXuGm
GIPfQ00tifvybGVh1srXeDRsGRWdnRb3dUlW2adSAawALl+86kJ2ot9bzjIesKml
A99nDr2TZTf/Ql3sQI1EgH5Hwdbd8jT/1fxRuRceLmGQX5aSHEKlfE/xemb3c8s+
G/MTW0tVR1PDk0NexjqLOftTAcchcrr3VqYupeFfBhL0PGwQwHuUVBaRreTV9ajo
5OuYz0gWd/NHs1bQwMD7KDPHg5Wwgu39cIEoWGEfz0ktCxvitfRAwc3uEnfPhoSm
TB7PIU5R0zIuZSJOmdn2biYf6wBgb9qqV18d+/EnV0Na4mLWeuj7urD/h2df3DiJ
KSAGlFFYfuuF+DOVTX1H4M8XFK4oCkb5IN37LlCzkr/PGU6xT4hGCMcX05zI9LnV
2s1tnV27Sv+B+kg3BL3X8efY3JAA1lIJkcPIaCYbmJ62zxhLIHcY2vh93ehW0cVf
aZiQZJyuLUm0crWloq/v1N1GjlKw2q2ZeVuaoBQpXpQlkvUI/45Q7p2pe8SynUQQ
0nSkFve1QWmlD4bJQ656nveH+BGEmRcTbg073il9q6skY3a+ptDdj1eA6PjeZznZ
Yp1OE0vDxBkwM3deLLSSSrKL1yUs/exUc0NF/j+FLRM5aMWXMrV0oRhhtP7TKdyJ
+MzrRRt2OGbRtyhnzFi69m4EAMxDMzLBGkFy0ag9nbEfy395hIqZwPv1JI4eKO9H
wpfpDdYgCdhJnPGOX0T+OW7Ow09AyR6XTEVtkpLdGnXd0+U7ZxXHvOBdsv+MNvTl
pwg2iOld78xCMSjpjpijwMpYqWO88CXtB2RRHSNqAIclzkvh+JYj2kKD7dAbqgmS
w4tqFa257MRQs65jbtDRGjeajRHx75R3wD0S3mLNnSLG0h4otZMYjCbS1wen763Z
oJuxPNF9gMy4mZvSZqvJw2XsDjuCmEwInu2QrUJT6wUmSYZYhCZtWUn9QQMlRe6e
aW9M/LBIb6YOhGfZi4ae1eO/ly6hjEywihciLcVSQwX1jKvHsppESt/h8sgrGRth
sPwZs0nKcuu1c82rJFbCwgCQlvR82K16Gx4OEBYT5Hd2mLU0taFxN+Lokz90hRuy
2KWGaFL8sky7u5w19QfRk8zLntAILkTDsiZEAJlmo9Xs8lFwwWhH+3EzkfZfYepV
Xw4bofuDUTMVc5rkqP47M8Pnc5PONYC3a+c7QFahoIqZZzyzQMVzwh73PxoatPD4
54EfvdtAcRILtykmITVkgrci4DaIlYvJJ0SbgSjwyqKr8vhSA0b2/DIZgjtlf7/t
NYnRfKy9vfmM2JpHqLI3/LGJgUHtMM9ClP69FZqqoQiak3PmhRsCHUwZ4I4tx38B
PUfigAu3igzFqlmBGMHAT97L0nsd+VbOjW/28RmvoG4p8e/9dssqDTl8N4zrWG0M
/8aGtFprYYLqSAN08or1uQnMqk3Wfp2f19ufzV295vX5M0iOENIO1TqgezoXjBpH
uqcoZwTGevepzqzyYdlEjnBJpnR9y1cD8a7I+JpgRA5SVCkEtmDZVNjary+ZkzKT
sYH5U8a9232ENkn+XjUtjjncYj0S4LzoVzGg04zF2Gy7GTlAXDZhiJedTrR/8KNS
pATAeEiJ8czGHrWllQLsDIYX/RZgT28g5rtXiIi5uXjANayQ0XPmRjPADAQb6LpB
npAb6YNCm6CTbDP+4CWp2gIGMoNi4mFVlmv9KIZb1d95q90yh+42xIIZIm8uGsfA
ldk7iGdd9mTRtX7+9q0kJqAd7BhJdRFUhld/7OL7TUqziXBIUAwUa3jJL8UiZj1o
lvnTSbBi0/u8WUWZNRn0C1Lr1EaKYzOFr92A/gXHPQudgt6EiE1WZ5F1eXhMTn9B
c3DdxR1figEKKKIpMVlMWdJ4Qm9TgEg7L5qkOoqe5vKFUJFaf1HYybQLMhq5HEgP
2YpNcBJHA3c0VM/FGzhWZOd6iWaxVu0tTA24gouXit42tCPU2H5BBsZNA7bSXgkB
t6kotLxvPOU9f5XoX8xOfPyyvdMlOBcttVAOkzMEo2hSDmMPLRDqEubkUXXDVvft
6aaBWRlz4ZSfaOUcScJKXf4cOG4t+6zzAegD0EDv+b4TWCI+ZAvhMCCbm8eN+Jtb
Gfvyda9EMSNpFUVXkbtCOst0/X8Xm3QVk47PSheT1/zKh7EZqV1i4/7Cn8uXBdMh
0eHQmH4eEoE4HGpo2GQ4e2KZ2rKPdH6JgZciy88mj/vwsyYld8VwXHqE2w90C8Ti
FUYaS/EyPOShX5RUBJ2ncxdUtH/0egPXlOSkh0AfT+suwGeX2omBRS6+KilIl0pH
eFOX8i79ArXRHFyQAVcHauQYBHvdrJlH/Q7vVAvpfKnGP79WH7z738XTAYLFPo5e
aYOaLf73zOmr3C4yEmbTgDiGs0bb80Y0wSldDhZ+/FPiFBMlo2dPd5qZxzggUh84
86xgwc6W25EwZw1UG9wpAH0LpZn2UfWgqT0X27RDVfqbrHosgONslMei5j8qOM2Z
zb6pkyHR30lgSFA5oGky+81M1VwCBwHq67x/VfmitVkcnR3EGtCwgQIY9Ccm84ds
B15JF615eBiGDgUrzV0MSbZGyd+ok0jSWSi9ggeJ1ckLR21rXBBD8Q7QhzDMUaXr
x/EH55oRvOnNWHuDH6OSb2QF7MyFmhUv4mon4FEHEnGFUnFI7zCqpLP+F6gp1gpd
kNJJvA88cHNSB1uiCit3DrRfFEQNvIENe2A4sGNhLEbFx//jwMPwmk9TXH1qjpmG
ioE1L7I9brDApoIVN7iOS4oQUhUQfGQ8EmSU2Be/i7WDaEBxViJ2askiGoOgVsIr
FHgSEOXK7bBNRhXf6iCfCTOTtDfjQmEs8WCYMMoX2h3U8+hp257YXzmBugwPL+UT
/ygWD+JJb8UKHnKdL7JgZ3K9QQCWGgWPMTaHl6pcBkaGUNmI0fLlXcxj1OUHdySV
z0YEusOXxBAlbx28HkKyNZQGqj+HFoUxii9xGV76EEorue0odL/i12MBaaik58Wz
kNnKzmqbiVVJl0bb3vezLe+XEGuEU611Ugae+dK1P/rctFPmIOW0jXRbEGzOsRz3
gb/6fKAjE9UsAB+RlH8xggDWyfYlN+CZtT46oq8i2+Susjjg0HdKZkUaZLEf3xkG
nBUhCf9tH/hRIucoTagRj1Refecoe5xQ27pQiSkyGuhZVzscFmWXI8kqZ9UdmpH6
ed1ANmf22Z6zU0W8kdfHLGv9/3EPfvZS+Lzcr0irnORt20SqQdnVv5kHh//NQmx5
UbDbgSc3pL15DUcdMzJqey9bfpW8JWoyo7pTwAq7xcKhZ8PEPH52hsb92hF+6hjg
kcRTM3reG/ePTObyFyet78aFxRT42jZ53mKSb1MW0E/kL8oYCw45OmQdqd7Eeito
nD2ttB7nbhJoSYUVh2EPtoxhK/OcDpbG+AmKPOBgZF+6HduIJLDDBFPkRLpqMEWU
46QaUr1YATZhrqGFvQMoE0SSI+YUgfvugrDNfYB0pdTDnDIZmW9eR4uVyZOK47YW
SAgRr1APXIgbBnt6CZh19Yz2huMrAIyVPauT3LniIPY8CNY4ysOVMIOnB41FRzdi
DuNG/YBOKkZsFls3V7gxv7hwjytrjxhL9ttJKWVRWnlK/HS4MW04BsIb5YBSIuLq
/7Wn+U6QbSzbMpZj4TYKFduVaF+FpLVZ5mRUGtXNloqxoxcB9qXJI3WYbbiwTpPt
QQtDQsw9ZRob/v5W5QTj+M1t+MzfEfHPnQPZDyCn1N1cc+nOqpYVHlo91Mjhp+ll
TjUYawyaS6NCCDPH06x8uysgGcVY1DLMXTukEIGa9paNUQLRk9U/vhQbZzb2+YKF
JoHX2T+/iQxmkgy+OafMD12okCyU1+N3uFTRSd+RV1AJUnvMOipKGBdr7uxQQwQg
pD78ePWfYcI15mPiIP9oCidZ/LYdual/1qfk40UYkkHluK8RBADAyU+6+6fHFiyM
bh5ipasvKd+07Q81Jp0n9UwfyKPDRFr4SPoCDCLbgCwQi4oYQ9/dZVlFlBGcNt0e
MiKMdahsba/YowGumosLRnmcLBnLuL8GPEWJmIib0nCZ/FgnyhAOGoxwCqvGU7No
vR9+lQg5+47CBEj6qrMoGG/OXNwROFCqWdr3u3wU66R9/1alkwIbnU1o3pqpXLoq
M/2vUzEmT1fLaSp6Z1Ietlmk51c49PRHTH/j2WTFqHnGYXpdg//kI28KHoG/wSZt
sA4WcVaZXqeQsWOS/0YNVmzK3jYXYO0+Uje/dWynGYNgUXZnamyq59avjBQOL0Qk
YhUhSbssWvC2e0CoRx4BZP0c9S99voyL0MX0dsvIFS4RfU8KgWTFsPlIGjLDl6yy
P75vEUGd1DadhnJFHfX/lVF0YNVVoB+A0fAsdbKxQapgHQbJ3Wl0RG9Y24lX0dlk
C5R/pDmPBat1Q4Y0aMf2QWGIjdKuAF8iW8tfu4EmdX0PQ/6R5UaQ7k+NLqcyXyFp
N7cPMqdkiUv8NCEVPQW+psZyoSeb6SJNKPpoXHfntvJKL04B23SL9s4sj3UQ4pM3
i5iAnxKjqcE3YRic3CKByqaJl4cN/GslMYsTfO3BR3BQ35Nb/Z64UkQTQII67mAk
ZzuxFnRUweo6Gw0huKglxTtz3RQ8WwizTCeu71dTf9hHQJTkL7XOYs/bWJrN8cN3
QgTbkCi5EOK7xmlSM4yt2nc9c5RrE2puG0P9/Po3TeyO5uF6Ox0ETlLaorUYLqPT
gkToeL8F6zBVvB0SyuABB1AL0Xw8aupZ0pMQcfmJJjnA5AiVsFju4WIl8cZ3FmVh
LOg+D7UYaCOWSpIYfT7B8pgRs7vgO13Yo5TlfnTReUeUnj0DgGGLoeNh9B2YWcx9
Ql3fVGieePqtvXtCAs+cwjsmQS3DvrZ2YsmnlWy3qmOCqkBHY2WNGUijJI/4K1dr
WJ4GlIXETaIVjFWaWMyEDwzMvpFi3KwEvDFA3eTzsduHGNjDolF+2ABKKfEw9I6o
t++f3moLNDV1shXw/GZMOzi7/VCif9jwxvnQ/d8B9MQ93wntSHLZvj5iiw0ES/Y5
J2u5/4YNKgerGVPAnwuOyxXT22hAInyqw7vIBf0V3HP9ATTHu4RCIyiKL5k2KrEQ
t39KxT+7luE3GcYNk/T1DFKf69xtJm18fJ0mC0mNf8X8ylrznw8UAe+sep4fM4EA
DpXfdr+x4JOoP6IbNQ5wohD9PIE38HDZNq0QhKEJqYZiZo6/r4stNGpfIElGQ4gW
Zsky3gp1jBJ8VtNywB8C+5YD54Ya8GjrEpRzQLCs8INXWhPKsqTEpAi0/Ts9huo0
EeysD3h5ELBJJqHL/KTjlMbIBLWlf1oeaDfStRqYaFnbKyZhjY43oHsp1xfpFtUu
F6oyW+5ReuzbSOlK96c5UR495s+zKN/eqtt4KU3gcEOaJGUQCa0yAR8yDvbFT7Fb
ywsEemE0yeIz4qiCssttEyijBDkQwEtX3zSoRnbsbo1T+d1cd5iZMHvcn/N5fr0m
UzY1LEOXPyfK5Z5UyPZS4kku4qN+Q6OqQRa9SDeF7vMyP7ctREFTZo1tMIgCqE7w
HQrPZgsbC+3XDKoT1W16AWhqXCGDTaRN2J+BTPVwLbSntoUZQH1EM5lvcmZ6b+QG
L/8Y0CbmHF/1KxxuHDlRWPUinUBZ8elGBTCB9Ch9xv1CoGPh3I/72i0dALH9Qwoj
5ZaQqtVvAXubkG5OYgiBWZUT18Gz2DrV8MdLMEKhw0kENzKXxZr6ZGsXfmU9x7sT
zMwRtSONa9ZhVJRcZlAaFGpJJ1VRRDRi/OZkm6l+LtznAAiCz5YfeiHNnZwjNp2l
h8y5bQAS45Bss00+BU65bPRc94NKkPzA+AsvUHjRv0FmWGMMijCB9OF62xihQ7fD
aEn+BWmCgbGh57mtZp/gKDffqUwCGF2/bqlcJ/VgR+zDCfZbXJFPy896VHOLxo5/
pHPgUp95Yvq33f/v0bgrgfB+kLy9F0uB3A+lsbB7luB2StTgsl3MZQ1oth8o0eos
l354dYlLVK9RpnctFTvv10U8B9UupAKH8YsAvK9kHuvpUiWwc2k5HpX8pWSUUdoW
eE3b0CXhWokdkLLkoBg2hXkKM3UiUPjAMkK9rxkUZFeATMZQ+n2DzKNvgEWJg4Wg
n/s4WQIP+URHdyGk9OaEdo3tQMUIIzcN+Fo4A7EPEbBOVAzNUDJSfLPSz3tDexhR
0w2Mkfgxg8k3ol1g7Hs0rZp/2e4VdQP7NIvc9eFoZ72UX/Q6yiYhE+WIAMAJPIk/
wGPh/TqX9zqndauN3OocAaOf4mhoHS1S0fZseeXa10PQAIj0V4t3/ZfpKNQbUmrI
cfQFBznRXcSeY6NgMA+DM4Uzzs5SPxr8+PgJgFyeNMIawz+BtOPcCQpKYVwKiK3d
r9QSoMX9DcOpvxIAosDMTLFlExolBLmTqfcoHI7zqlLAd16SOwSyEHV6mlVE/cj5
v9KTD/XGYA4yHXpk4HUu8ZKXK/Yp1pZ3iiWjIj6xkdIuWrGvrZlprqorUcGt/Zas
FNPUZwMEadeBKfvSIV8k+4QOcc+bcmtJVgxuYqlIlEImxIfaipaBThduB5UlSQB5
s56Wzz0q6p3cuwYun6lVw/5ncIaHkrFy3k1Wiem6AufV4HHYYYJWTJPtcFcV0QMx
TFEt3lhTznJCwJ1OtVZXErctM7KDRidFPxQUJbUznr+RNdPE0WlNq6Gh/qb/fYdh
lFYexclOz9UPp9s/bH4rcowjkCD6xnFHVTxQoBB0gaijuGNj96oBdNJJkGAtw+s9
oCqlb6P7tDhsPuczy15YKt2s1GiVyL7QoVXMXIOn2p8fJHVOWRqnK4hFzU/hw9qK
TivPaVDjE8QqYLxQIJzyWBvHXZ+bp1eOMeBLhzoInAAkyWy+lL3z5O5yNcwKY7wP
nkq7bsZsJ49AZ+RBDvsPB7RUG+zpRIm4ZdEG7yuKw/EHjAt8BOt5xsI7fNwKiWN0
8MjfdVRXPtcYAHm5ykCTPeoB8LMb0bOQMzyD1kQ+mAQgOm7eRdqGbaRD+odUHo8o
wfI0ASz4FWCUPCPCFPtCQBRI2R7aC74UicWw1pEWiVnp082zjGsWw/D78SBYtL58
JL0J87bAW9KYvvf6fbeN/U3fpqUMkXozzLOK7AKPutzx6kubEH0S781ftxUUjbNl
YdmonywneFdBExNKG5vyTeYpcjWY+23lPNjMqdyqK+36ddXGNQYBOpelo9a1d6Ug
4O+hpI20+yUGBJl4sl7f8ja9BiS4gazrhcRryv4eimoBHzBAK3Ir549w77jUtAJP
fWdm9gpY+uer83Ny+ek3OLDeMKINhbeYwrogA4xBJutcHlBwVEwDneGrOjVP0X6B
+rWnm+tGEIWUdKfg1erpQYDw276Cw23Up4uM3WvwinkAd/44sfHTqVrJeMjo/Soh
odiYD7/nvMj+ysvGJALX8A9rvktw4MY7hmnPgoYPVFiiWSvelBstwxs+NlprRLi/
gzqAcb1lsf7P+TbIOHGMyM50bZK5scYH0VFTTm2i4jLbyudDuMvvJ0Y953HEmGBK
gsHcVJjD3CKWVX7Q1rf+wk6W7f5Rft2V3CFYwHw6Vvu5P1vq68cCjTOgYYnrYbjK
yRBucDL33g8h2GTxDlo4le75WDgzJzP+hIimNHmQ/teGjbRdO2YQh6/E9rNfUurE
gRkI4mtISFy1vbuaK7lCxz95f4En3HCnGfz4P/sBt2UZwkOoXJPgTtwkeyUKEO/A
c6tdGIa8ZdS0hp75roB2mdYntpz33FjNqNSsye3ytnka5LcJj75OEgFp3EPQJU3n
BuDIHb+fNcrZwa6+ijKS0Qt5FrQrbyFs2xLPXZAInovjx6qRx9bqhG5HYOep09el
OV/9rhBlsBvjw20lK/ByHTUg/DxDKXHXoodgKVRhEgsA7MnyeEjoR1wRqX1b4wwO
NnlhhoDdiy8TpR8axmHJjGuul6dPDby9w/fC5lOiUrgtcC+JbmWk5vUEr6pmhZlg
f7d8nhbZWUb5RS6E+RcW4uirrp/HJOZ+Q+C1MfrPhMTZ92nJA2/b9k5jgCjvgA7d
Tcf6qs0XO91S5vqkmgZ5/L3GcxrZopZtwpvt5lpkJgIM5NYNfbhtj/azJ5ZEUGDc
2YJ3chcLjVr+tGKywClGDgEtjhDSCD52BggOUYc9+BFOo4A9qe9KBeAwYjTj2rbJ
hX1bp8G141fqXXxkvjuXyCX6gE+nKVJOU1b8LaSEwkWoctKHz5fdfYt6RWlos02b
Np91X/aaaJdHrKRGyy+4KIp/+5aPzqlcC7AUX3wgScbxb9PteAsFfM+Pu0kDgoj1
AOQLYjOj57oo1j3Bb2aE7J61VMxucz7ewxPVNrsRjA6w57Et3vm92UjF1cMBIvxR
o6OcyY5DWVKWUIN8uc0mmDqdDZ1afMWVy+yBfYP8aje6HaML5VbpKrtNP0ehbUGC
Bi9RTs0b/QmTIL0x7AN5ZjFCcR841ZQCC29is/4h+FhGc6I+os51IeHWNU3AiBdi
DxaW7dQfQDFlRJOZ5WbFUQaj1iMtbJhrLRre+/6YmmctAmHII0mC0cdoajqN8AiU
FFuZA4SLiOQzSVDDdAggn5opR2bEMs0I/VfpXE5Ty1iKi0PzfoWbBhmRLQ+1v7bF
4+KmEaLOJkmJd2RiWrkHzzOkmaqM0xFXcmMqnowSj901zbw+8J7+EgpO/QaLOfUR
7HhNPSiLsdsKO66tDtnIsKpi9AcZYz+b0jMADdByD9HFM2iO+MAIxuB/qt15R4bd
Mmh8s8QVNT27QE5GgxYWb+tGwMF/wDlnF3VsmMpmoarO+bR1+Pa7eN5yyrcO1PZB
a5JRIKAQ8gkGDK/WF/3pmz+FgsRhmbD8wnHm2kmXbt+mxQnWGk6HetgWqU4F5wDJ
Ps1RCMLEP61aDKCg9qWohUXgvqI3deKUHhRlKqE3oJzRtOkpFGtCJ9nxMcNqJMux
Op/tkB9K7WBhxXumpZ1KTzhNJgMBMuOA5dWG9tK1E225WZKCq8+G8LtQWxdtC+Vi
AAw2iox/X47GIbpSwfGlE3wzHJhLnqCgpdxP3FDLozKg3v9JyVETsOcc7/y57+qE
RLNgm3Wt7P9N6kUVHhOs2ahZIiUzCij3P2MynICzI7hxcHYweEfnrsihKuM+MLq7
fpz4xsuR5SNAhLhfvjwUFX5B9+jgzzh7JK/s/JclObMcDDN57dIvaEWo2BYqgqt3
eSfE7z6hfBm1tqIekjPLLFbpdLFXBwk+i9adJEXTKDFWhsMW+ReaUXeZpHQj/4gw
S5Wqlsak32aggcDt2Rhm0zh9Ied2NHT2vbZGiI/PM8sZWNszPQaEDl+l+XFNK2nA
4qQB68y/iGeSy/9EG7rXHSgSVeiYft6EatJz/15VqpwWglvjkqiNFnQ1aPrVWp0L
BTWSKj3NqsokglnJaQBjQ7jseD+7g27RH5ke4YwzjPLZM/gFh1lNugZ1kto4Vyoo
pp5ZtewCtQCfDJhUBOpDLn1XqukoUQVpRffGo+AIedgwtbYQzU7tb9o0kMM9gshx
BgG7zysdpvs0drC1ZB9SUykzHhP14j4ghSNCC8dOmUBWJ4RQMOBGPu4Ul2wgHH4C
tcxHHpKbkvmjLiO99cWd6uvbDEi/AjbeTmexfJ6cxspWHDYFGYVdT3LSKKk4lC2b
9aLLqnJ6ppEKC1opasauQgmwdK3AdBXor3I12f02gnlC2J8/2P5KF7OEoNT8Qb3p
8/4qXXdgTfncHPXy1tKMrKtGDPf5vFnraU40RY1F8xAwL1seR1Ze8nk9XWt5jYyK
SP4ncGqj7Kv+/rBHtA9uKDrl70Y3upv5AnssJJazo8IHX5hI1SU2JJHpJJYf92DP
1rHPXvfZxMRqXQ4o1/44r7Gg+/LlybtK7hBh4rv1roGUXl6MinDC3fqn/ZFC3nZW
tb2sKhkpdnPGXlhq13T6AEuwE8J4EBcqDxOiiG9GDqvxYfr4/yUgUl+efwpP+R8N
h+DAInlEIC0XSW/J6/VkUsacALwoBUvPgL81jNLX1QK3wNMo3oNy6NwUAYI4jDzx
WtwsgAdz0QTvbw2S0iogjRMAWoZW6hcJk/FnYLXGG89JwGL0ByUdtzSc9fTELpaF
RV+JzIPcWOnrr162K19Dk2cU1NGxU+YcOdsog7dJ4pOkTxm7xODeB23DwEbeeSyU
v6cnhRNFETh7c0znTgY5mb5tzHSlQZ7364Wf3+MbYmXruMeT33PGkiEZEOpSxhJY
pdC5msDU5BkCMspvOINQLiyuhH25/KTaiaOPE9I6ryr400ZnIx/5jMx4Y9dZe1+O
u86hRtW6KA7CaXj05MQbYEfkhjmgPhm9ENja/Wbs83/p5qjANUjYLIEFr3aeJo0X
OO0ep7iKmcJysovx5Wn+xjbtEwkexU0r0zpKJXtRoBlMkchc+hMv0HhT7O/xp9bD
pAS5rPgWiy8RxJ2vSmqRRqO/rZFqxqWHswboi+GQ4RwAL44QDqUWV1dt2T2walg3
9HLPRn6yLy41PBt0E7BJhbH79LNkagvoQutXY2GnPJ0/4CQzSGHWHTbbj9AFuAvi
LpqgcPZnCo6jd/oOX65gUDCSUTMtv8RC3tb/mQtLR7ABE4hYUPeFV9TZTB/bhnEl
r5AKQNeWbSXS/zbPtz/wW31wDVC1WjVbY/ZLqan0XwP0EKfKVOIYZZGZAe92qQ3d
KoMpdR6IGWZaFlipIyJR1qRfKG9r6tpW3AzYa6qcCLRL5qQId1RydzmUN0Q1wtL+
Tr/p0Bhnmy8kT+x4Tn3C6P3LboFU0YfhJrGTI4LGRBHntgpFmgvGxLhqWQVzjP9p
eNAMHHXmib8Rt/bDten8OX7bHjrJEnLjxJvqGxaPXbJZDEaf+Qr8bBPOsvRtRk7n
JFCVoUFkAJikUG8Lr8rM47NhmoxyGKAYmLX+hgD+HllAB57FhTJQKPVali239Ys6
QiH06//PleRY2EyfRcESN9Uii18B5ujIOdZ0yA0hIS1kMvxlzu8pDH1sc99ETCqO
tmv2kMg5jJzOindLXZVUKc4VgItFXURkMnqeOVqn+K7gebL7nbfJkZSO6b2xwWp6
xyMSJ/MMMu0umK8fQKz/r6SQXOWO9+Ajn7ppyW5JJ9j7furmx1XctNPleK0p0hEz
OPJb+Gm+HtYpGNXS8PfuO4mUabhkY6odoCcykF+uO7fVgodhZWakXF7aT7d6dXG/
kDlX3lPY7LI5rhJAmeQMkYQ2rYJeAqfaz7aqyt53VeQnlrM4cbXGGkpPn77mqjQT
L/yb45UrYtaIdPcMNM+lNEfGZYbv3JC5IhyLCPlb5wvoNqRWvHOI1oZPZaDOxMww
4QEZd3CLvvDGUIdin1tbtz85kK45Cb/jDm5DRgWAFfSdTtQ6m9qRfkc26U2A+hKB
OWHdoTpowO/mmeDaj8zekj3bSqP4me9FpT5wFdZylsTjwuPrzC8/MNYMNVfKLRU3
QxLp2m3/Ss/BS9IQpJQHppCQAgFe0xPbfWm23mmQy/GPJsjb89ngIJsD4t1qEIk+
Ir7VUB0uNHUEmQIjTtpCQ7QXAGFp+sNfCVIIW8AXZo80oJ3jTehvFL/S4NULmkUR
zqwN4EsmPKx1V+zXWerKJXKutu4948ZTquydJZC/Ti32J29qTB7LFkHYWsmLJ0jZ
0eTQ4Oa2ARVLLY+JeUnSAGwxYsK0dYDojd0Fl7MKi8e88AS7CvAxbO+ZGhGu1Z6x
iAZFweirJ1AuQ2T4WQbPz93X7a0fwuD5aQu0ItYGK6E+PC4uHzT3xtRXzlBAEGoC
Gc9MK39agb73jpXmUojsL4H8oD+VegUJB4Hq71nZguOIlQ2O1Ql2jW4FSAkBwAkD
uX6+U1i8W3zQQOZROI6b4Cy9/qUY/RP8JYfAbqnhHDKTRiVgV2h4CUaH8fCLaR8t
Mp+3qpm0EFN5r6ht5/g5pcCuXCBO9GrN7+vFb/C3sOUOiphjDadAgVlH4YSL/WgP
eDX8/UlezLEu/vPtAyZ4lPAQZ+Mh35a8mmztCQzRHbvcBxBph1CPMtE1odBZFg5Y
9JhkaGEkj8dL3KqIgM8GBqBMEXm/Rxch/HcKBtXw/fiSika5z6BXCNXBqu29lIWE
cJPBGpJm1hfgCvGoHW45gIxP6Tti7uJ9PhwjhMWcWGALl+4AdAcZ0RoQrTo39q+s
Fcu+YkDp3lb5oDz6B4WAkCbnjSiyrFVJjVIpMvZPm/Agvt9IF4vzTHZpVFYjWwMq
yPRpya7zUUd/ojy1h1uSTUtGfU7XrAqv0hoKsKoGb947Up7T2NCoHPt7RQHStP3Z
k4U0Ovkp69PO5WfZr3kCquhRKH1oFUklwXvfEAL9W3eFjHKyVqFJc1bJJubZoBG1
j5tQqZFfM7wgL6hqYouthh6I47mm5en7PX4Xb95NEs25PzkLyTwOFlLhQ7sVNABO
8DeAk0xiECZm4o1NYf6Z5rwhw2KfKtu51a8UTE+dQzXF2ZY4EjsZ8kKCYAroGd8s
HWmh6neUQsy22Hi32uB8n9yCewU21UuxJkv7yd1FxcaODOyyEqIX9cgX0k8D9eH/
seENkCE/pcFF9zq+pCJBt4mLBc4rDnBdghdsC+yJutp4oaYhnfcttkYqO0fuPMwc
pqOglMBJMgeIPdp56qO/muXZ0i3rHSpQia4gMFEi3w+V9tricWoCHlXvdy1LuQoQ
4yOaU07fXuXekCIwBl2CIerhomnb6OgFH3/BBkCQr7bbtWWC/5KaVd5wLRB5+9jT
EzUHgL/t5Vd0GAjARekVE8wpkYEPVaUEBPzPIWSyxNJzoGo7faUGyb2X0ybJJQRa
EsuJqN4Xjgar3lIMxXJ0WmO0cTWI3ky+of8uW85CWMZIxOhCl0+hSg4Ho8Tt1mKt
v56GSq5OE8m3ZRIwFMlECexTHkb64FlwVeYzEvAMl6ymZrNj/bB09CiXDu76joLv
1Eegfio+L8f7KaTztOKKDpnJECjBrcQ01KZqmTOM1DWANTTjRpA0N4S5a3oHKbj/
JjaLDBl1hXOaYg+VuCFyviIHFEknqNHh29wC0+e3QbPCvS/SvTL9k/9xYEjpfV7T
3z7sgx5wZat9yxMs/qepWU4IlEzWP6E2sEJCD2YVooaz8qUxMRzi7Hmu9YRM1ITH
K4wAkk839RFb7KabjTpCnXLNDwxr2BSnfiJSggjmC2sb6/DgPGkj/3V0DivcZf0j
gpnTARHkooTmn6gf32aO/kuOk3ATm7NfF7bcI2ERYP1cYwUfTQedsZZYdvvlLdpp
zRbKLWXD5WVCwsJkYHZOxNHAJTtFT1y3LpgKpm7nKQCBiX5bql61bq2NVevPC/6n
i7EioxektPJmZiH2f3qrjWSBHboTOAv60wcw02czlwN4KW6B2EaW9kJ1jmGLDb7X
BXwaK09G4SYDgq/iKOtqRPUPSMRuKYoSSt4g8Mvb/lE0xL42s1qUej/VhtxupkRd
zvduZ1n9zc1sD+Bh54gXa4aPEnsauUdTfLcfEGllBpmP7Wg+wLIsrkiwBfAyFm8v
kW/Zan1IPEUcUsT6+8EWcIxiludfvIJTc0Se41B0OxH9p8ekrmtQPq/6o4T0JXI1
4tu77xEarEqCQYBRFCROLWg8ZOmlhI10nFTaIsHQlkpVo+hAerAzLMWFObCxprb2
4iQL2BvFBS8DY4+KbLf7yTocaEU4+wT25JONK7vssuwt1/NtdpIhEFZIKCyyH/Mk
NWEB7CtYIxLFREMVEN5e5eVi3hrBJ55V9Y34KmmmQ2Fi5COT6OX6B4woRkOLwnt5
X39ztTp8tCEH6Q6m42paBj6jR3JrNarp5ALjHZl/YktwrNUrbhOuMmVCcEBAiPEG
gPTxifHc318JTTtBMlSiujMfeqm5QRqk3KdvMsHbbzLLRHUasLh6CXLu4DGN0O1k
EvjIaq/m/+7og2ZqW5M1yVJO9jlPv9d27mtXbeqRrJKJHs9seBenWraw0wPIvyp/
7XAFn8/NXrD/CqZgEqz9cURIWxdlfad/amXpYiQYqSgwp+b8uSF2+uFSP8z+3aEG
BQQyeiUcxJrBSgHgatmYm5POGle7DKAmcVtBEk3o/o1aId1mCu9npGd3JTHxfkRP
bCkYXsTBxI827HKLtiGXuWLl3L5GoJ9m9cEUOFUbIdmgXpIT48Hk/LnVUv3zFWo5
KB2+5auSRnsCS18dR6bCiQ80r0H44wXk7SZT5CBzWaoGgQA9u3LKTz0ELD9ljzfV
6v9LKZEFLe/mRUMfcREC4BCXED5qIwLlzkk59/WkatVFPy4tRtxd56KtArs8CWZh
/NBzqwxt9HqJCLIJIFFyMsFz65TRIhdtrzyvbN2QieVx25sLFILT0ZE/rN4y7iIa
/C2papsF1i6NcSCnjQuJKkI27JgMfA+LxT/IUsnEOGL9UsVAzhzRTDORng8X1XEm
xN1WMHaOleJRWpz27H/d1wCv2l+2aBpDDHV4N0doKgojKuawEIb/7I6y36IryACr
jkf9UAxAV1bgYzF6fEvBhTqdR6JXqxeff6ar7/RFgpWycinSMwG6R5dLIBQztaCO
SwsoE9ZJaCzSBTqvBv7c5HkrDDNy1oASP4CIqeVn6kljv1z/Do7Jgq8GKojTY/z1
8EAwRL2hRh1hseEZOmeIitnTP0StRCmJqVc/wqjS3yLKKGjCELuKYnzBIvJbat44
xmYR9fmW7sPGthfsX1AoLF75A8EIgPHihrGxT7qNMcyj2SIUt+abJCfCbyfRsLaV
FVQKGja2WLEXFMU1hUMF1gk7nkFeALvA17ej2fikB+bqcSPUg3Kecuwkc6W2A+FV
3axdxrWHIyH5eqEPmqiCg2mds5SzGMiPBX2DjxlS1FZ87ox9oczm2XqCY6vrodoI
r7M8SHwRdgD1uQxdcmVOUmI2tNKh35DXtC8ujMwo+Se+ujRBLCSJAu/Ok3mmD2st
R5a6nURHkS/Mz9HAd4Uf+sgHhdsRXZoLU35wMIOrqTs/MvAwcpc9y2rOH3gl4v6r
uxCXbSOdKXKBqW5m98kFysZvAIx9PLQSmNnUVDeBLiiefVEk9WFiiTQiVTJf9LJp
uzjOw6U/3/VN7sCa80zMmsj8atCySMHeRsDKVYUUYuLJ9Cv4tKNukCCVO6CLMLfK
26tjdWy2WcOXDK87w3j+C+WzZm+MMtfHfEXA1eF6My9IZ45yqhmd7GVB+1g61LBc
DdBWrHKuk3UjSayJvw12grDWt8dhDYdPbKbPu0qv3VfeuG854zaKdN2fnHFgv40A
Ca1uqFiCVHl37rFrbKgiSasgiTufjWUB06B0dp7Laxis8ksx/pjEpF+DrzLxd+9I
jJ/zOQIVrELG8pU3CJTdkUX1n65COMLeSNi4nhhRuP4vMe/Uh6FrC4dNF/aJQdUp
hzTgk7v+XX2bpS7TXNV87hrL36Nl9gY6tjs2IT/SqC5rff1K1N/jRSzetJDISX41
8XMIp9l7opz618He0KtJOkIQATf6LL2BCOegoGl8BAzztI/6M0d4GWD+y3znTKPJ
1fA+2oKHhr2pDDGoKA4vCcPZjclJFsWo0VIETtIJzaoG0FukkpcVNoU2A/vZKj3E
uKtKo23wsNgzjtvOnRy8UeexdANKdOPRgyBFQmfYlYilHjOqH4T1+qAIjYmive06
t0cSprKtMo8rRxdiig/nhaA2BV99FOIslrjKGUhZmUOjfm1BoP2G+fnqWf1GEUoe
UkezEYRItH1wI+ig7i33r1QwvVDAQK7V3wMIjHdV+G3QomQp+ST5IrizZWKJiwl/
p9vqwezRCVDQXgvk/meStf40bdmCwcKl3PBdeSNCDUmL3yffOcf1qMf/rP+ojgOH
kcE/wgRNPx3RGdOeLlOeTuCG7pfwme8WtHfnRCsTnjAw2uRBNn5UXFWQ6wwxLOzp
aDi/Ao3dcVnVz6UmLPxDRMMhQo8etctRO2RhIGwPiBevMFgg3auP+2+odMFqZBRg
6UZmGw9LF27Gx/8H66Dxi0lT0RyFFqUB1Rhxx7TZEeFa5e4zDEm4UiunMtqEKfRG
+JzDyRI8RE5Qp+ITLYOVLICFmMw+Zt+CL1z/vQhYK9hLBW3twgYjAiGrz3F8U98n
OOTXpyJa9wpBlVdh3iUwjiDuPH1YlPt47O1Pa6BP0LG2xFbuzNCZYLWxuMTW0oG8
Ry+MkmT56H7BYnRfPMGiQBYrou2PxZliFsnRPebNO+OXd45/sSpAKj831RlEW8lQ
D4YuRqmSztlHv00IpGajN5a23+2Tr6dyJGbO4NiMMoP+M4LGpmks7rZ10DxC2CY0
L+82XzklSGK2YAsDlvvvzaRLpulXLiNdKGyCipB9yD9kfHFz1k+uwVXzoAtBdsgR
KzcEL4SA5osQbgC/dQRYKb0PxJRgPSofHm3LkDpsnHKW3/3lnARaAWQqRHfHHM6L
XuxZ3fjhUD5Sgn5HbNN707FRR2OXkCz9qOvermQaucNU9cctG3QpzalwUeYUKCgJ
Fou3ICAAFMpBZCpfkAXS676CzXLk5VBs8v3FZu0Sgp8YvKF3uZZoGt8CRtfX2SPb
Pu2Q9Nw8Agabp7XYQ6VpgsrC17sX0a81gsBni6uZHhkMNkxp7ptSFvSvf/OFYxhO
eIbYxeVvcCeGsLuJ5B30QwzLENj3OuHl+a0EG+pFu1SsBYqwpY9qGw44ftPCv0Lx
sRSX5GahmoT2zRYlkuZqK95CaR7dIKu1uxxDb1AxZlmJc47mZUoDDgJMQwKiJeOm
w9DCUMZ9U12WIv/nrskvnprudozzmO+ATEsB37TRsMML8OwV6tYToiZpdCWyuIeN
Ki2uph6E/ox67750jclY3TG0I8gBXos6ITrzoBisAB0/Q6924QIDtCUR2PlpGaq9
vN6Z+WUmDL6cBgfkVgNJcU6ncBAZYhl7VoIEyvbdjrIPW/LbXvJBGxifD34sMMpm
Ql8nAtKUW6k/HS9QfD3zIfrVFv+lxS2wfb/QKKcWT8Q5gFOyzSi8WLpnEtX6OoaQ
t87EHyKPxxMitOgJObjQim8qRkkeW0TjfNXP8odAEXZ3g3YQZLmClMMv+Hqi+TfX
qGUvxdKL7YMK7SLNEXgSY8YStmcX33qE/3YXBg9YbwWuASR1qWv01498PIcpODTC
iX3DiXr2ZRpCePQKsy/36S816AVOQsmE35GMRF5G5on6RtpNYpJJZLmuY0WjUi3T
+GyYRMeRxaG73pb1xL14UetQFztz5jE27X621Z8nKFo5qjzEqhr0lvT/xVMkohh9
9G9DLwrWTydV+DII4cfIBM9tyfM8juxjVmPLJqsXHsoQNCVlAW6BkVN3Rb/UPswC
9ak5PptDtECpyLAEu6D/9D8BsmwLRO6yTmoymDp6r5Mm6OGZ/ayBZJgzWoKWbiUC
QFhoDDlvz8Xzfu0LUSURyURtzbP3Q8esb+L3jjkdEtsabQEH8KIs62k9bG7hp/Iv
JLygEBjFGjXaum1qWQpOykatzcyB9k/hUTLoB5wZw/rQ6N82hHqLkRaGf1ua4uZp
7DSstfjiPOrGo1W/OfQ+mZNfJKS1oDBMt0u9OplARxOYJXsQs6JcJ4j96gQwWPJX
ahyMmLnGINcQvsFcUAYMytY7ngBcQLt99oir0x/1idKsz55fiLdUMWD9K49TletB
MIX0SKsdo6wGNGKHqrhYS9UXxJjtBO4rN0PClMnZoTQ08l5AfBUvopMpuzdYteWd
GRKWXasq6WeC2DrLmGWuK/1zZ5fezvx6CooaYDNYnCSeEXDP3c2wBTFe2/9HGjyU
HNmdn0vpzVPpWzkPzx3DC+yKZqNnuT7gkhIX97gbMjOp/6Xqm/5MtmqzTFwH2Mqv
awrBscca8ehGEfW0n1TedUcIu9E5mlAOoGjxA6rnk/50olBHFVWf0hCq5Gj81ftd
XhhwkuiQHs7KNqO0YEuKmTL3YCJVtAunRmWCYtoq8QFIiNq2edVPbZg9QT4wNVq/
Fi5rKEYNZaWzfRTL6bhMw649e8luE2iOZeEbvp5UD84vkV9FcWLLpmeqwNj4fbvl
D5E+kATUvgLMLVHUSm57JJmx19frMygp05YWES3RRQpBLhQDag8djYOxXOMMmcJj
c51x14UNtf/HTjK9Vgsxeghp1epkR8hgSEMRHRuzP+FU3+SIlt2o4+KN+tiKqpiI
JAELViDBR3XRR1BRL25yezOokmxtxawULnhtZycBYYkx7R15DptManZsY8K3JFav
dndc8bg9Ag2qRIelBy54QTKHe/UOpWifnF9uFNjhDNbPpCZEGmgOggydYR8r0V88
HS7CfbzJ8CK7DYIuUgCs3W4Pd20eD0BhikpkmLIU5YrWDY+xIMJ9R8QoiadvAhB8
TAXQxT0JVjMks1Yc/DmYToOKLlLEKKQbQ/6d4Y+cezO4kOPAUFcdcTUSq5km/Foo
1sMhwAuPciACQJZT9AP0HnrDLOAYs2VD/8TXBPI+nd18R7ZVhuMh39ZJAznV8XE0
ZpELCAV0oYCTUzqXi556Xf9LFrm1CeoQhxztNg2DUMCI1NLIwWMZSfCLEELXCjy5
H/aJJSmtkDKECPWHlq59FDkG15m3m7YZbXdrGyuohUZeFftk/5uWbm+jt2MDkdp/
6ofrsTyoDU0yq/jyoI7WpEQlpU1hUjFdcUBXggObTk+lJ7p5Y4G90F1twNcP7ymP
yQpRfYcnJHzU8O7rnBy7eTNlNYzUH7ZX5Vdg/HxelTXuKEVy5BO5T8M8a5fgg9cb
ceGOBK3F1mo0xQLvjFEgjLADUcs2UStZzYUKEFIHsH0eqEeMySUe8ffbk+xfSUNF
0htG098CPGXVPiw1jkm0OZKwF89y6hmFjBUUiNXeb+dZfweBk5maIMxYXzA4fGbY
Zj/zXmApLHY6wYIHYMRRT1Rm/P0/MtFwC41eNEzukpP97IQ4fiSPpOWqK6vwWHHv
DCz3YaGYJSV/85xfbTXYasRFREiIDP54+lJUWYTMkebGbmM4tToJzzRfVWgWU8/o
LijSmTPT7eTZ+P3ESFKcQy4VL4gkrVMDUvm6UuXiIa8ubsmOsV0WR99HYxO1Ou9r
1enQWff+xdt/4LXYr1WuctPELg/BxGowiZJ0jpiGmFgWo9Gf/tZF751t7W2a91/j
9cD1mDjBdWStWiC+2YYf59RsYe9wuLwnLuzWhWA8FCkJjGXiYEymHAROpI2oPvX7
KDq5zwKMXlXOK8giR8aJJv2UZWFljn5TgtFfGmXAVTN7tcrm1O8Snzxf5VqJujHX
SJn7HxF3ghFsPrpgWF9c5/CyaIp8kjCvLA3LVKEInPfvKhgXmgsfPXJCm1WlFoWp
2Ttkhq5idgYR3oFmDihid4FcrKczIT71zS6wTrsWNTXD0h+hfuSOZsTY9DvdOLU+
G1rqh7teZIpepp3P8EVKHCXj9DA90PjISvmKb071HnhPPbH0DyQMG89BV1M7d/s6
upAQaOohFjNzwaIj5vJ5V7GbzB92/fm+eZPJ2205JKPUkR9iB7I9uzv1uXL1DmjB
huE3QDXGPRLMGw+PVIELluXUylbEWESuopjGGKWzSlMZC+dtBXI/+CXVkBLjcta0
L+moUydPzqWsLPr4sByH+oh37PYKDiha9SQu3FN12eK5iYlibhMhUpg2oeMQZA7Y
aGHWcSPeGRHv+De6o9hxWPa2XOhcmJ35wpIBeotTl7KSDTbIdNaQLr12tsHaN68K
B+aBBGxW2cQHVSv779de+K3LWbq97EGUeYgjR0iKsZifwA3ygMhVqurtgWshTQ1Z
tmQLRKpLnH2VWRhXvgy0/DqPnmrXCCj/QDlEtzINKZfLB07du1VaHomm3KKLY+P5
9ky7FFug4lR62PrNptmSrYCxHwMVJON9wFQv0ZTECBXhboRPz1AZELCvzM4q39r5
p2WyRIUWMwaEt6YBA8Gb/x2oHFnNKh/AYPVKHURlBSqjDwKX9aQGzNvekT70O1xD
iDCq0YWL/uSVyYwkq/wBhXoO1+sUIkq8rV5VOJThfSQtN5n9SHU9fuLKt+1jJuZl
69Q9Mw+m06k15a94wIQM5KG7c/NMYbAP/zCRIY8ZUJykaczbT/P/hc1fFjqQ1xpH
/ZANTpVjxDemmzfx1GP/pU8TvYHNjjQCRu77UfLD7O3Bk2IplsoNpaMRJWZjjmBn
vsZkc7jUujn9jk7WCe/9LsnvL5K4gpy7aBPydIQx13R8AKdyKvmujuDwsiXKEmUW
gCFlA76vB0fRzbEWux98CYm8aP/ewcFstJmi6N22nvnSW9JHD74EQhVEHyz1WVAa
ewospxa2NT4xFtH7sKK1tW/Kd72Iv+FxQWWkLk6mydNR92j6StaFTJ+pAv35YQJv
u3P/yXV02dfR/UhuIHVmhaNaRlCSh9AdaK81iMPtCBgCR5lIoy+sGVL2Dx9/Bz4K
5RikGExRsGR2OT9ZXiboZjhARIgfTdP/5HH7OUbFxExhlctUlgdWHgGqfsxA2v5Q
ZSKphlBJrUlsQ8idVtZ7w7E0xXXHNTo5Yuc4f1E7yKRD6e3yxiaBhyuH6NruD21b
KFcu0iq+J/Ps7SwydamPYQQ3kFg4vuy6HdYizIUrhYyLbbBMusg1Ru+D/EI5hYQ6
kPPB9cLXtX3G+9+ZQXoXvL6DjyHRxPXZQAX4HyZU8JSKVlkHdYWy0F5Hcj51RFjJ
zwiS0AZiZJOXLz8alTli36kkNAt6Gihv4lwpYkQ5CglykuGsImGRKIh5tIanh8dI
Lie/jVa8iMDtlfsiIuBk/jJjuOp9pP3s8HzQJjec0GYG/islEpgyvPg+mcDFAcRl
No2IeqGYrtSib5ghtQOR7idPaypRwyLxFatf8R+Ql9ym+PK+a2cLF/ttrsPeQN77
MqSoGf1nCFd7k1jikZQaGDL4DkQiEmZJiDbBpMK+HpcmqLJOm12npkINSWH6bcaC
1AzpNn1cMgtmcKTWD2Oc3Wi6UPpxdqyznTTNVyLQtfKSIRy2Uhn4o+oz/rOwLx7M
azTdsn97XfUqwXe6YiZOmpjynhOnz8CMX32e1TE33/CMbSPAa8yQsI4JG8penTh1
aJ6d+Iwzw/uG4ubizUiWWfjTx0r3X+kgzq09aQYYLRT34tcuK2r2Hc4sxsy1HiY5
e64jbcjPfjCPcSxrj3R5fKRHEDdHumpLL2H2P0uIROXPVXRR1O8b4Ws53K+6PEXp
lxxBNDVTCdBhj7Uo5n2bflJZlJzdFPVurpI6frBBexIvEZ6vN15603VgHm+UhFkF
L2AcODXmT00DM81FqtMe0MsHd8pWnJeoo3SCKcUw5+SWRq+gfaeH2J+KtW3uwB4X
jWZcySr9jwfsSY+jHTcFy96cr/ZcOpqfaq+c2aYHjIDo96uzT01G24TWvnIoUI2A
jibkn6RfUdb2IMEm9UjDfY7y7PtdNx4XLRjyde8USGaVJzRSRP5BLke6Lme8yhVT
0cuVUKkyH1WgXXNsFQrsds9ipbH26zYxzeDU8x//8TsuWYZv32XxOKZs+0x0FOoq
GRaPqTyzltgaGKvGk9dGTfhzJ20rZpu1o74jMYXzOwu2vexeCDo99cceddz5kPTO
nxD96cQVG3PHxkXphyZukL49mmuXDdv1HTETOTO38qPDyU4mFZbrTyNqercBYso1
zyrvmMzWEVBGvSYOlllH+RY2qJ0JD7mPP3fQYijpP26iu/lxfByvYOwmksyujli3
8RRmvUd+zwry0CPgQklq8NRu/4tqnbVotrTQkqQcyh5FU/SEkWB3R2arm1uK5z70
B+XFeO87jRAoRN6JJxfopOs+8MHsH7LzUBn1qYFdvvzifekEYDmPbz7AgL7MtKUa
fnnFQA1zclZohrp0I3BuC18KA6Nb+oHV7hdmBlzy4+n3Ut/SJVg53Krgm5ZJlk6J
0BqHxXCxTck0Hy+zcdfM3/GdyfRcRjuHJYZXI4zR3Oallwwy6YhAcxdCqg9LnAbM
Lfllfg8OLRS0elotZGyHa4+DI4IM8tUPmtI9VvO2sg57YxZFeFMg8Xe3y+0Z7CXb
KODy9eU03z0bjo02eU6LQLg2OmiWJ/bRtxI6VcelOa6bwN07lNpqWAztSVkKB6Gc
ItDXIf8XqNnLf8NxMg8Xkp0LhexJ4nqDAfJBmYl7Bjx6Nc7HrkBRIlUjzP/lZHwF
p7MF9HLr3uaWJrbZ2fidEdwv5CzDyBkjzOp5/XhfJuTTsOKVcQp551NOJk83ETqM
gJSi+H8uyBNgS5ikv8XAt8Sel49Nz5tU2Qj3vYa7q2QTnc/FyuPbDa9eOLPpZvE6
VuIGwVnWN4ul79PK1C102Fc4+3j1L2yhJDEMFXpK2GskhCkdGLrGR3zFv1AFL0fM
EpSjaGDa9y9YZ9d8m0sY0O9ZvBGlk6QdzrUQ4zahRdFYiOgJ24CSEQ6OkYJPwzIz
zZVns5pY/LMOyti9ZgttrlKG0Zj0ZI0Hj/ta2Aa2aOSZIY1BaeBIKW7uoZ9X7U7y
nQ55zSOJkdTZJlQMBe7SkZKw990SeOP5hoicRmFXNITx3HKHoSSTogyETHqm0/jV
jWBoSNijfa2C9eGvJfsUe1dwjlqJv5uD36+OYE8OcaIRLstVfSP0xCuRqgU0PQrB
AwNOj2EanZdGqXvAfpNABHowlXSJEy2W9TIOK3P7oNwOg5e1lu+OvkSaCkPJczec
wCp4tgA2KdiCOvEbz7AvrQLK4KDMDJw7ym0wyp55yC1tS8mhOVhdi7xoHRpH1rHW
9RKhermlJtm+l+Yc9LnNe+FnPJhzs5TIMHgcljn2ILKtCpwyjqm8FUPwvGr0Gmd8
qoS7C27RtQrUDBsxiC+FIifKs5FuaoiMlGiH0VPMboRl2+oYA6RUuVo7nFvnQP+X
OZot8Qh1ISvfONkaWk4gHTnKCD/Vz5BnbjJP/Kl9arcYRipHQYuumdXKExY2EoDk
CdLt1V/h7uHbYQjhhAuhb6bMS7zLQn8BW8mVhsdAgMrh4hpEZuh07+krNk3IAI6L
CFpE6gnyYWY74TQt12l6WmSoBbMfaQRVXRzniefrLf3R/sseoQZfpNpaub/VD9rP
CTLWzTFyryQX5S+0XsGUZh+EX0zID8pIpEjbtEVV2fUselORK56MWHN7RBhHdmA4
rcSq78SBr9ZH/9zdaIlyQbOwx7b+Wx9SvFw05P94iMXrN3iTqCZaUIPqA/T33VPV
1oDOSB2Se9a+bgvvLju3PXiTYBkwoEBPJ/m68ue8k7WNEqg6NN4dCv/Mdjfo8ctY
SjT8jtEsI66KSOxbTOtYIatreLYJj4Ur2RAoKGtAGyRSHdsn5zTAQ+XLbDrhL0yf
8M24FweUkYtSNe07KeKQhyuxvuy2Ez7XQJofYeg+78vKV/Cq9xi0ynAAHKUh/QBW
1Jx1/b/CQ4lhLYHhc5VnU36mYY1aZLXeCLBdVnugszzpsbqy+/ZvECCtSVnoxZKm
+8owiyoDA+w4f0RqYpVAIdprq8P3d55QX2tmu6ZXJl+jNGujcDUj4yMLRK9E+3Go
sZc7xY9ahc6nVTIocuIm174Yz5iI4mfbyphbMl3lJpaz7Sx+/tlBv2zcPOUTDPyo
M4O1VxCx7UfERBsAo4oS/8f+ggWABQs3YbHVs7U8AWDCF1BoTIfofejrOH/Nm/pf
cBXMkjvNVOd6ZAZVNQn814yEkvrdDk5rNMm6Q8ngvDlUfVe9kfKJB7EKJrzLGXqt
1HNDUTbpCXgr67teKozRu/JSMJ/yl9TtMmVnulgkF6ws/wUKF1zkRuPXxwXJwObJ
aoth7I4GUIyIj4Hcxz3EIpAvM6VYcV1ggj3xdvTkPBuEsVL+GvIGShodszFXyxyU
1i0ZPcAmBMzkMxnJAI6H1XQy9P+fQL9cMUfGfsPvNalpofN+mfvEmCIPtZXfXKOu
xvU1dchgBAjRA7/JFnEdN3qVG7Im+3AfBhALpluDvSnpfZMkme4JqakAfhHsK7P+
RhUHzPA42JixBf7rkz70Wgq07GTb706ot6AUVaE2QKZTZCMeYlaTxloFJ6xfo2Mm
XnWnK+ZbKtirsCEOibEtfpFITD2V8PHjIFX+tri85YKAzF26Z/FHi10VY8k3MME3
oCPPZMgeosHtBOemHeWs/mYz3k0ReQW0w0J3MX4LSKLAwex6onfoMEmccp/GUSvO
iVk7h0h717Tkj6eOuwkMVgup3SXQAdM7JzKBHrhnMJfIXWPWkh03vtAoln56lQOB
cEiOU0FeSJLgc6KDp7QO4MUEouHwFPqfM90+oFXfevkZ/Fs1MFD4poD3XZOLV/5Z
Tu+kPHXI2b90wR9Jzu0jeH1hU/QONFnVpi0pHjX0OkNMhouJyazIIiEgIfUbwWxc
Qc/P0j/R69YM7qkpJrVm9TJl+UBpSaC2EYFY6PzzLUz3whe5Bm655dJfQmZPqtLI
cUOrRrnUGX/pNu5A2vmBkE55AQnc+LTdFXa5ngJqV+gnrL/B3atS33Q7qoewH+Cr
2Fpx+q0zgoCACgK1avMRGxj5h0Vbq811bwaBA5fFA1VQv9XiRbHSXSh6xOWuJYJy
HN+N308Q8BZlCMAVRIjSf0AzcdLQkz5nkBREzKaw7yrRiAk+5U24Bb2oZ7CwTZKv
xwdUzSlpgmiK23XDGgHmkVSAODLdijD4Xe8kBHUUDgd/35eaoP3K/HnDdmASpn15
aB8f6iO8xKyZLanXGm3ikCDCaTcYoKr+ZIP0KafCZWkzTFqMKhdXt6G7erc+Mme5
wKzQAhPrZbRKQlsmz958B+UsIXX//xsuE5hhdzLgmYsqg7gBL5Q+Z6A1egZXy15B
7YTg/ZH4trlRyEcI3ij5ulDGxXd3GJlHsZOlaxAqXm3ITgMpp3+7YCI96+1EYc8g
gXHTlRB8WgHYjTpDrDJpfgp5pZ+Ur409xDqLj2VWTIiU0IVHbIkMWuKgLXDR+FwA
qAAdA5rQ56/lCWD7wam6675fODO0JwPCDb5gns/MJFSJSi+C4devnxfMMX6WOikl
jxoYV7FGjm285jURD4H8xCS+JA3uE4vvheJwfp6GW1oQEaathzUUrkc+yGLIrB/r
7IUUERMptYdP3EQkbjy2qvOmOYwewBn6WbicD0f6P5I9v5ptYgc8Grgitir2tL8Y
Ri3j6UvwWpVuDuVXHnHJ3+ZOEYSuVES69iQ4g1nIjLTeyNBjRFKquUeMXceWxw7u
3D1D3Khl+h07I5//lO4WBsufv7VV/DA8AfrNUkeyHkh7jOdVlvFS1xdek39LHB2+
/yOpLYyi7R2LVnVIEowqjW6O+GxCC64dUnwS0EP+el12q2BFFa28m999y1Dg1MsO
XKBbkpoVNOIF+kIHOWADh1FCFv62a2k8tZiKKnkEvpNejdSOxffqoi0jDZFh8pvl
/uuyhmLFzZW7x5IT4QA//BjLSFtm5nuixCje7CB4jjM05AztwGpxcFkTGQtBdtw/
HFZWT4sZ8bZc1tVnrQoVs3sSBYxm+Yd7tTQV9yOMsFvebx9Dm4zqEh2UY2B56/vE
W0ONPhTZIhqwGvxLIhx6BZEO5D2MLZzdwl6nQXqMOlJZAfXXxbLKuqaIoHCdZ+UI
fqJIRc7wfAPiXMZSkJrFCTx+Mma7lw0rvactwOcVN5GmK2IO2mUnIl3rPsWSfL/I
Ui1etxI4GCt42ye8VqDqdSQu0lz9IhFOFQgFpaObUp5LqYsF06j83q0E2oRcPXOD
2cV+4lV0HCi8dP4pOsIwwH0Gr7Td05b4c56Aucg9zZF8RM6w99UQAOxar1s2ijs3
prx7i7tCNVQ/rbJP38IuTY0SlEegjiALiHnigmzy5Iqojuww/IpJ/x4qtnfw54qq
T3omRSLgM9ctskAictPsZJyB/BhCLewlGBnUBgLLNw9qwuM5lkhmyIf2pU3wgnzS
hFLkHujfHm7d8D70KFtC/uEkG8GyD1YA2ehDNpK/4EZJxzqTPX6Ct6D5RnKE6G/O
WbwZPXHfIZu3t5toJKFMcnL7kPnPuCiRwIN34VuUjzXfz72swpSqpC+1A9qPHdzp
fs8OhDxVai6xMhvSSueDA/zF2DG6G8Tkuj90+73GjJ0qmQqWNLFN0L6iAx0+s2sA
2GaUPvsOL0VpafVSgI3ou1uQIGUQhlKqHE1ZYXevl1WrkDxpJnspHLSwt8DJWALN
MVspFL6ZSuoRnUhvWw6vgYTlciken26Vn3NxaSWP8uTKFzBlORc080yrEm9Ft2+d
ZYL4DJ8WXw+AJvWtKOV6i4VW3f7M09C6crrl33OdwE0J/H6csV9kH68yR3btIjhx
mN/RbHG/iZCWiFD6sDmPOoge1LbEa7+IwbaTcUJZkSdj0DkwWGtqezC2LxBQh52e
GTLkn2mrLeryCPraQynA9V2rcD+4Xs2acNXxOHv644qHT3Um5uGPIRNiicSRlfX5
JbhFRuiUCsKzihq+SsJLE0iqWJsAFD+Xlivh8AZCjUXMRDMLTPE1zCdlsqNPGU2o
PCilbtzD6ZC5JfxegqLErAbeyphujG6QNs6U/IylFNlPT0mmxnmkIPt5mbKMUBNC
PLS7ONkwlwTEZTzMsQQXuF+eDXEb9+hHv2eMtFAKONR9SKNZcJNTBB4Vx3fFHM4B
xzpsIqJg/Cgkl5V5DZgXHVVL3U6jY9ScBGD1tmcvHXNW7ekDTOeYGQSrdsYTjmOd
nO1kyiCySvQaV+oMkE6Q7Rv61Q3Sjurhs5lveJMCy4pGRQwVHof8Z7IgwlO5iMJH
LqkSORF2gYmenh4QMuougIHYxvsl+VyAi8ZCmfKfB7V6JiVXd9fksbctTysgb3HR
lorSLj3fhaXMyYu1m/4s2HUGlCtifjXeOBT3/uGBmXlW5j5Jb8eqTKlTT/5jr513
DkHzAYUaWYZzGpDGywC4b90RIq7wYAgzRV771tU31WVDpf0SndXfCKLxxTFhVdD8
VozgO8CgvmXjj8bmuhetoREf4pKIqoTG0EfAY1gNgPpPJD3P3zkAg4J9XAZ3oGoG
g4Qmj5LhM92ioFl6yiAMVv8zL3qhyjmcNAI4vTVwGm75DBJl/cmoK3EsveS8cYg3
GmfD9h3eKa4o0TG7o6pdojd9lTkwySbCJyqcf0/+qp7ekjnto2FsvSMBaJSDkhWI
AV2Jj+B2nMYVfsNw41Rck4vLXN473LAzIdVjyFxpWmh7z8xrpjcdt+vOp7bPf9qS
lTlWYbYF7wO0N8wCcdYit94xxmMX+g4Je8NK2G/+ytt1bkma98FF8//ooRu3M0xX
7Qu2BBx3uuB0LZxZwXKjbfaILRC/Rwkq3zEiWAkuzJcGXe6Cf3WQyfhbMRg5//0w
vIHCnc7AY1eE3Q8gv79DvOHWyvLy5vQb0o6ajTf6n2mLdTOLqjew57YpB5kaFxMY
MMewxqHtQL9WNzRo8Xjs248Ziy6uOh4SUdNo75tCCoPQA9lhtruIHle2DXdTFt47
ggoc6/ePp0+AXTgwfG/JNvm3NKxCpt4qUtrCwyf3n5Z1CpJjHYddgM8ligpCDNfn
uXDwT1FLjLL93Z9/W8QEjWYuzv6/P3khS+TpwbmaPq6omivnTdfoBcKSjC4v6TgE
HjMXfNCo66YPTyFnwORQRdEb9eIA9M3STGpH1g6YT/WM0jIQJ84cA8mDwmcb0ey6
FU+xC+L9b1uapGiw4l6fwwr6lsN2/JSzog9Mh6Z6AzeieSpooCpUil2ZS4tnzBjr
ezPxswUvtH8p5Ol49IGykidh1fH9XZAmm5qUH20w7qriXnQZG8hAay7Z/eaRqJ0f
OqTE6Mb02+OoG0/Wj9FDjQBHDrOdwG1DtnyFbBMLdxetxo90CxmoJo+lPHcT0Xrw
Khgov3alvppxsL2F+doQaPzG8Mj59p31IukQ4NQ7sQH9nblSI9GqInRpiARPsnZc
Y3IUTTUFWsDkES0f31RSpqd4yIqW6tATMMelW/dz7MQIB3U3/F019YAYbViF77vr
Bg1AX22tskFvMj4C9xQAGXAa+FGP/patuvWe62PVS0AxgLHXM1UJWGuV8xQJQ3EI
gcSUze5CuO8oGgpHi3LubeIumKgazLatcK3CtTxfmFR53EZe/m4h4tMcNP6yioje
A4KIMuNTd9ANAvP4kuCjGcuUZQqBkrfE6DM1wTpYlGppK7iLy6vSYvt2/f66qVDi
IpT5GwGWyrxO7GtohKuBuvfKJ+D0rwmpe+Y/q9VxZLBtVxYXcxx4IKhBTnt/k+9x
/QoJ/HFgOYL03BiQoq31e/cCwHQVB7+94YjR7xspMxUuinYhvSgtgs+8mYoPixuV
N9jC3HpW4NUbDv7piXd4j0HrWHT7nEidcILuVoqC+VqTPp8UkjsLTNIjxcRoRssH
vFrSiX2sFbl2ZnCWt0XjrZNdRNAbYas9CXCoCnkRsyGdWGtf9Vx+hM2n49svumDE
SuRTTcr0RsULcvL7mYe4bMEma5tA3EgdZ9hXnt3gW7W3pTzW5v2XfgWqzRPyvJ5z
TN4LrfWL4PK6xzGZzZr5WiFzVtuydoEFVaS5lEzS7ZUCu5/6Te81WXj1On4UvyHQ
p4cjNWVzEDl68pQB6p1RJCE5rExWTm67PDBU/iqSCUFXIu/e6I3Tdc2pgfApL2wc
6wOBRCXdSflkANcrLmJ5JPpbl538QbVuDWrY2n70wPqzmHYXNiCA+WmjGAUySRnA
VLoAmVUXGKNxZRpRxzL/ZbBNXEWGLAzZ/EnJ7a69q7tDRr0zTgG6pP21WEyUoKZ+
Q89Rrhuaxq+DCgN22CoC7IWrK88A157BdXKE3JtxyPmolcTVF1NjU4ZMkHJqncH7
QSxtCLlcfTwAMxbD6AjoZd8IxgN/XDz4dPALV96SyGkl6sNgKWr83sLeglW+uYEp
SrLw+ANyH/+t760xefnHt/7+S0R+WlCZSNhYmotlRKfOUtCk0MelAHlpkEOwBmuh
62gjw43LBk7zxVXfaECKWa1M1w2Fz6x0ujMCoJ1aWOIO3LvRf9i0DCVrtm3R/266
zBO/rwa6cxnQOw6gGZFwGse7fCsu6IBj0ofobjmoXtn2o9QrovrxdCsCBfVr4xg+
1vTo9fJKqA7WhsABjHZEkWJmzfTq6534G5bktveqEMbU3WWcL05Q2jBxFcVrO/Pd
NRJ163lSO70DxzfysrgtZil9lVt+1VnWDDb9htgacC2na5pTWw/vK2SZlkN/gEQH
U0bEuy3TBYihBG4gIzgSU07zOLw1iUx070DuPemWh1Yu62YvWIony2bVv7kXET5e
lhWiRVsFb1bfOsxSW4T1ebENh3yMtvpMj7wTfjJT7S9Wf3YodHmodC11qQ2M+5LT
dK9SHvXRs6yQa/p7zl70kZQzG/JiUzS2PojtGD1yc17wlqLGG0Guc3LHRE28l95y
IGpC8JY5mFOsSnPcHRyA6OtSrn8d0YbVsVW/c9NzhZYnHRImNTcfsFu2v1lubq3y
kh7lLBDTF5DTYdZJSkCSVS7z13JUXic9ZhKMaxEoNGL+23vnwoVszXfCL/xZ8gfj
pkFjUUfIOwz22bwGC629MGxiNTKybC6drkUihwXfke5uWdieWcRY1+is8h5eN9h4
IqiKkWtjN6iOUkF48XDp4HJ3IUqIDF+T2fglgpwSeAR3xEJcbYSKWyUZD3Yr3agh
ZsoviRx6a6wb3bJTcaajyIWLFobywFjUgW89LnNXIe7ySr0kgxs55AW0ROSqUzqS
q62AT0BmW7UgdJYMXbbDT/xoaA58YXXiFM9KIanVWygtUZrSBa0SIZZnAkHPi6bF
rqZ/mRo9/+53s6Sx1zNOfIGPog+5rb6aP6QyFQzC/9a3d1MOTjrdv9ELVWCZ3zXz
jrkM7Zdf5hQCBc4cxdw9TNR/WLTQt1TYpTanBuU4NtaYa7TzG0Fhx8TT8K2oHJzR
Pq14NV7vvkdWLAtvJNhz3oV6pfKhgdMcnRr1dq+O5bST+qBGPWWe4XRxxcOGSowz
Ed55HUISa9I+I52FZ/REYKHEr82rtD4hx09BZwnv+PzMOzm0Pvu3M0HU5XKEfgQp
ozMSt4s4DTFC+PzgJJYFahAlPM6UHg+XNo8APjXB9G7fBWxQstQ59aKnsB8cd9Mf
B79ptqFfXjyYS69CgHoWlZPlsua1j8EmFgC/qbX7CG8+T1+zJRFv8t83uY4whXLT
DfYoOQDhl9Vbi/HZhCPFKTlAN0LH8isl6vnq7ogSBHq4iaeN054gkb4Zxy6eYwzG
6YkoyHnFc/pcI5Qz0XilUYZ43V4kjpUhWPVrvGXrWSnzF/xiXoCd3Bd9cgMPsR2m
I0v0vz7hFaNKJgiS5Cd7SYqIvW62l2fVry1mYpNfwJbL1bwntXs6XTQrOLbTo8NX
rALXqs0bHG9GWQWXnQd1OTOkXorjaBZdz1zD04X8VX3vUxhYLbnTVPIjQct+3lrc
7HzvHMWau+oKjV5CXlwdc1oslHfUe3fC7tizHxVIxbLguhZYZu/f7/VyeTG5RXzH
09uvCspKtKaCqpicaDEQCUg2ibHT+5hJ4qckiy65oI3OK77GwWph3d2BkmVhoOO3
mj3RPPJ30JoxJ4+wq0JxxKcS5HPwCQVjJQr1TP+hRpXbNuP9ZAQtttj/DiULFqdn
Wg93yXhZGqtAxAxpFByeFje99Bn4fAsmxQtHaWnh87QFdcebLk3BlRaVztOI0IF1
HJADwPfGaFVgJ5KgrtdGoPsp4W8ZYOIZHAWKzUfaAvB/BdO5aUY3YE9d5x7cdUrx
z7wIE5MOOVvUBr5L7b8gflQNME01GlHl8hgis4nKwqtsSO36iQDOCSQaJsTHrrW3
tq+eajHXsAVdWWc6extMOgybO/OCpzzDTWlckNXZahwureVVpAFVPir+dJQkZTkI
V8jJesluTsThskljVwLRuTmwiMiP8igBCPnbY5NeSD6YMgaqg3z2pm6oiGK97T/M
e7aW2SAyl+RISPOnOE7U+NtprXkAWsgBFbQEbltHz4yD62/a1Mvl+JbXvK4r7w61
JRpPdDfYBfMlKrIvhl0j7utwTan3itB68dc2JjGISB2y40PAzFEPew3TBEr2id8I
36F7M7voppxRld4WrDuCDzpQzwnA222bCl6shUuG93037lkqZnAMYFZ+hDjnakQF
fQU9Viw2a63q+si6WH7u/BackAdk1slMMDgagLCa4GAFPXwifkQBwUEK9vJHgfg/
QIiBeAJEerCE4w+YQ8+r6+KnGNkNqwnVVQC33CAOeK6p/IAn6jnIVGOixDEDgNs0
WDXNqsWSdJuawKD95xDzF6Q8MOaHwft0Ia6G9tL/aAbhQfsUnuBP5h89Zp3L8UHp
5Q+RttOUfuswezMTUmwWv5f3foBvMhPokHWU1QXGocNlBDsW6V4PtD7i1bhR1NO3
kjWsA+68HJop2JhGRCsGPoxEKd26ssqhAjCtmBcJOYHKfuT+Dcd2OAquCigkXZ7F
0IVKQZAPjpFlCdu7meB9zYwRL9x3JBOv5Ie2Si1jVlj/6DGz+3NiHo0fgJXdpXV8
NrDO/HH5cjN3D/7I/Y13P1AVGMrZnDfJgNcNQJqhyaHDgDK9jD4R2RIDwpwBpeWr
uBkw6eTIHnePBPvwABksjcHzz01kWSlfel/caRFM80Ab2mMtKeHBVJtYlyuLGHmU
O+X3eV2f/NpvkWjKZHl5M9VuckyTxIma2uwRNKHw213c3o2CyY/rl5RPJ6w9XVNL
X1odSldxoT6XyxpwFigbqOzSW7uIBEMSi+Qhn9n29BwNIePi4wxCo3eYgLLNLhXU
rLgz6GcqiNlEKAW7ZsrSW+DQGzZIQlpIPKVA+szyWloqFnEjL1P+LEJixNdCkHv9
RXz1Pzb8QuDIR6we9D//gxXEoTJ95i/tqcOHoA3XNg2WEIPR2kWKHnZoJVuP3vlp
ZPwN4ArQ3qbUMgWcR6f8j/I7BFMKNpUtwmkHOa3X75MRKrJGVpfrfxAnESLE8zDl
EcZ8DcRHmyznjhRC4uAjsgpWTOtM3cB5zdHTRCOkaa+vcQzN3eFAn8/hpaod+Tqt
zkLeeJ+0Vk5N2eEU+Lfbdw0MzBX2xHAxJN/yZjQksDPUY0lc6yWRLeTd6tdwlf9H
CdnHJmqrIvYJq+TC4kX2oN79ElJTedKXK+6ABWisjhJdE8EFIeff5LrFb9iOMiAE
nXq6NxjknJ8RGyt3vx0SvzQy9ldn0MZRYFpLVkG7pV4mXyUT152zNsgj/1WA22sH
z+/u+u7yTZhm1R7GTk8AXErE8OJ60VBHdsb4Z//gVki2XSqkk5DexTjfm9GSAu5h
0E2r171Q5PDPtAH2FiddH2kMalY1SXIq2AeCj/LXF5B9oYV+dsOFysBekdcCVKJj
ZqhAZMOk+uty26Q1EqfNZJpnBetGa4U4D1cZjlAAKxq+uE4RQqNc3zzYOBJW7WUB
WdmoviQ9JrcrBfLWyhEJ3Oh6tr6f0OU39VYxcca9XLuTb/NCa+7r7S+eN82xVqUC
ZFQFFkGFvpSY5nNuSqW/DeyaUoa15B+pmicjV3jw29Z+TUkw1UBaKdC9BsKBuyL6
K2j7aVQIk1zFpL3IoMhMH8AtPLLAhMQig6pkJ9lmKlyXdRSdURVcg+80NFyONQBc
lUSVHS89TprNYydW5CZtoPQUqW/SklJbL2uoW027Y0j5wqK5VAShzunlDq3rBos8
Sc1Nbzj9EN+ESy5OYiKEjiPoMk1MIC7TB1zJZfrFRLPd1li0uLJ2VO6j7F7Tc5J5
v2gNtgj+lncAX+yW05bE4bKDCr9MWCuIGiYFNL5G6NUqTk7L9Qtx3YHRpLIFPT9x
borkFwjqARs0AvvHYYEME4bOoZ4t+prdoJHJ++KTRkPQHpSvllI7IByDHmKJTS/E
qsYqDHL/VRH2go+thpom0NbaESa8lb4CsgWrP1MobcPUpf+GWN2RMzuLgVA/gKTr
7RV3bgIXlBwkGdqG3hqm7RajfxgGNSqR+JloH3fUxVlfizW+t9PYVdcD/Xdt3BtI
FVas/F3BW1ajhi2zbJ52KLdMR7D+jbag3SWoeHfNEYSwPjEPeKHBddnNKH7+uEBV
J7tuz3cZriW8sY85GtZcHWz8h0ZFatpj7IJEMSgNehvbhzpkfHGeuapVRkEa2ab8
/ScapBeqj5PYAoTtCqOTcvpor/xxIJBBXhRtgL/txMwbZGIafYhqozjC9dbkSHVj
5KeSOprkGcHd18rw7I1WlO0XE3mN2ilhVzSPFClSYGWjczJ59+455T31PHNIobj/
/NSIYTrKKUIGyVZxTnzrolfeQsa7FXXyY6e1nVfapx1o/yUbXBjNxnbTJDO35RFh
Ob3BITo/lhvMdcOarjAODfzxK8eWoDSUcj5w9qJ/5NAJ8WqmrHoHu8VaUYWtBiHP
Lovg2Nivn7yiLmevfK74wWYEDDLebFTyPO6MsXIxJ8wg+T45tetAxBlmpeNxMG1u
+QIYjz7VPyX/4C06KQ/C+jiBfbZ1FYDyaAKvO4/VTT5YQyHcjv7y5CofBQyTd40b
Pg+u92YwduMYsf3R30c4Bvaahdl4Yz3g79YZwrys0cxeywAsuFb3cazYwTw+IyPT
nIB1YpDLPBCjERLjfSYRtdtxr2rosK057+nfOUw59zsGZ1NazI3vyu73IyF43xge
JYDfrPxPreRCKAZ+Dt0gYCDCQljqbkBd+EL0Lld/QXpswT20H0q7YSTx+dugFc2N
LfjmeXRcloL8/6Rlm8NsAviN9vx8YTLy+YxTfZAObxg1PWu+t1rrhhe87Xj5xS4o
lieJ98Y1dri8BHm4eGZbHkLGfD9gyUE5xEVJEN3vrWnFGSLMgXjlubMZ1a9He04w
kqJe9QA9EBVKhSnBV3vgWxuRPURlLk/yMs5BMFL8U/OkYPSAvGfw7VLU46IkmhcT
0D2VFC6YjmqZgBl9ttTru7RTxh4hYMg38TMITwar2a7rInpZ/ZrorPXNE4gAtk6k
DMMp6dMUcYHqYfUnOXRSOxv/c+R/HHwPnn6h5YGZhpXt/w4veR7VOZBsqOAyOeOU
EbItXSzcnmT+s3r2BKhmu3kXbMggiFoRi2H7owLOeR5LyoUNlVDsMiP4NrMA9F5g
4mQCA8Pd5AdH3PxAcdM3x/bhRDzvjmY9K5fDU6krpKo3vhuzr3xV3f7Mf8nnw5L3
UN+6Dor/dqCFZX/4AzVETN7C00bIPirwSh05wM5+6PDxsve+8MlVaAJL3Qz11e0I
jAbzb9dkrGQyMfzBZpy+C/gNzEN5KJOG7sHHBIRKCFDLO1cAleYEJg35xWUwhnCE
EV4QTsDoGdT3t4A4di4pSYKY7TYJOGVJunIWmKXdZOlG+MXhwhUbFBYkobMjrAzr
k2vRAZkcUHQQfyDtJMaeacxrfFL4ndMuICGbzKFUS2gyespy8QgbD/XvSUOah/eN
YYZnWy7c/NolWbh+kpcpba4dDLC73BqyY1cj7b9ipPgYIiuPIlCMEDQJlzUtm6Id
Aw2CCvjg0fe5SRspwYtYUy2uItVl168xN6wPt+DWIWjDQwjzvbW6bAPi5gUoVhzd
L1vVMbokbyFOOUxb6+DaS4Oia3Ghtws40ti+iPOtjJjvHDjkWniVhBMUMbS7KUJl
lUtzmPc0vRBaiFZ6jwl5MXQ9+U7LQj6VHIKv8da7Y7995D+SZF+mJBt8uLWc8HGd
hOyIgR5MSKM1k9NWmRGKAsK2pJe82eMboMpUAYHShiksGdbPO/Gjqdq3NVdo9bom
MdhJdDIP90vAVI+nR8pFDgLDLFoiQxYgNiT2bbU1uNr/JK0v+qMJHa5cZw9X+RS8
0xgsT2QaMHF+PuNghnSUxqWew3PUtyhMTYvRuz9qCLo59HZ0dsxdCqRIgdqWLwL0
p9Hnu6KaXK6kXGzhB0F3wyJoRdaCcq371aIxVNEOU+S2Y+gnp803yie8u99bTGSr
TvtVVA6K/eMzycQQZGzx9+3YiiWbEBonoynWaQtkO1+DJoH0h9M0Jco/2rq/f51i
iUvpkyUOyOP63M1PC1e1H/kOHpPTJ2znUibjbY7rXq5NCbSGni0AuH0dlT6+UOmQ
qDwjxkhFZ31A/K9lfxMiszmk2ZcvJYKJWIc7ESY9rI2rgs+XNGN7Z0C1N/hZOgbP
Siyhi3f6wsX3FjA96xBdS5J2/ta5Avlk9gY0+VogFWA8nJCXZZHcTO1KV1f1nSFa
gN+x/LZkLfhfdtKu+fzvwBj93lJs+C4gbcuhKCi7+cpJ0DHFxjYcmiLJmvpK/OHp
MzYELfaObBZLCxm6s40oxEINoZZ4WDESBbrzX0sRjIVqHmUMR9VECxC7QcdWPebj
nvlTcfRTHtosxSv5Z6KBEcqq/BtCtw48I4CG5AfI3U5dyKzI6FY7jubV3/frUJuV
9yvsMwQGL2SZWFOsCVYPNmsb0KKt5sEwViLy3S3Z07lXO1Gi4SiXsvGsVEOKOOPq
0ML+lgd3KP8iEA1e5+fJjNCh8GNteQfyQlxvqTF72oB14cFnT1/pxooWEsEjpz5c
EozsaCrrI/CHbysXFKI9vakGQi4JAmDXMx/uAsCk64kEbOscJ6XOwyddxW5mA5+y
Wa0pYKX9xSraPj1PVAto3gTQxSARPaYP7NDuhGYNKYutr0/pXSlNus8/FvkqRa/B
Four6YMndmcQQSbRyacDLhmpDiM2bfktKR2OTGgrm+AGCwYlbPSroEm2SdMnqeGr
GpWUHHsEvNxV/e74TPv4mAXfpWflc2Cj7Y8OU6r6ohzrJ3JXevZSQCcOhhFseShi
02eL8NAbDgINRb+OVAqhNB4mCXGyEEguaXXJixOMBiYM+J5c4ENKPqtLrgQCkgTx
skAaFJBZ7z1sUx2Z+R46Qq8+BfNR3y1YpTmxgPdOCZBoCbSQh2Tra6qPII6v6JGG
glPf99Ofs5h2iMzpi5uvH4ChcAejBWd4QE3bsiR1nBD8i0vQh8WVYGcQl++LgP6K
1YUUIZ3In791o2WnyjfzWCQ2FuDHltAPjQdumx+e7PrVMGsg9i2a8f1Jn4AG8hzk
Gqhg6BFbAtw/UmO1H2bCPRHUVF7/PzAOSkFxmxTt1Jji6/G3TBiYjR6C1CJ60NGT
Ol8FolYklhBIwG/gk32bZ4H5xhAuEon1+1cIygEnm4xwmjJ+mkxajKz6KEe0BRjj
g3Szkjq02FmkXrIwUGBiK2Ofch/X7diUezBdK10BZAN0U8VpVjH0PUpr5DzIsBpD
uj7Op+Ct6gglXuhGiqEaDOVY0WtqTYbeFCkMz3Rqj9PGYZaBAwnZuJE/cV3Q+6Ch
aVl7ILHfhs6Q/FVgzLdpCzQ7u0vnMffGRtI98eSACRcQLUkASx6FgD6f+xoujUDn
iTB+N4KHnBZETz/DkZ91AIlDmoRNRkebyio3M1lCkQnPf/yx375/lP3/eKgJd2IZ
bl5kg67hrpWomQsxG9eQABnNX2VQ6dkP1r+BwOGSO7u9foMhH+mrTwTsH5clDVUs
HTO/prqhddz3UJWcMVBMQiVF0aj3gyvrTwuehWI/NyUDm5+ke9HlTQ8tzu+DEKw3
/TAB1q9EyY54utjD/asPfWUt3kHv2JWkbFlGu1cL/FNPJ73qxarE5Gn+5MKAygTU
eqc6K8gs20VTN3VeL9jghLPm8CyqVBOnNRL0hHhoxE/Ylr6muxmRBUX0n6lqw/jN
Ho8xBLmJMzftX8/SB3M8RvyLWrSIRUmVr5Q3ooc1qgvich/tqqzotYE0GFfUtzpf
iPKlmEkte19r+SgIbXZN/R5SkLN0BaMXQHdh+tFXcAf1rJOuAfQvvwp28xWMk+17
+ryabhOFjEjrSmAmzJTZz5To+5aVWSG11BHSg5QIa/gZMzLcZbSkM8da/spmM2/0
SlIvFdWMThkjU/X6fPPahcwDvWHb4aZPLV9dcC3KWUChUwQ5OSveYV0XxTPkuk8B
2dk6mlNsKlR1VavbnsjLQKa3KFAHUrrZ0UhKLD4fL3+m2ARZI1fkdwHIEfAJ3efn
jZCNN3BHH7ry2Miy+2ytjUncEaS+7Fsaolt141PBdIVL1fBeuoS75ebHdTwSOGiL
j4mERhsl3WbB6wm7VZX3GRkagLTg+7ZjYcATEBmA+HXBHhzDhWkHF19thMt+86SW
5yDwYlanus5HApzbwvlNTv5QxEftXh5665bWgMcppOjONk9snlgQysdoGlLmgEjl
Tq82Xrm/aX02paluLiutqomRtNKg21OImbD4PLbSxGkH61JqBgOQ9n39qylHujXe
o17JhHiJflqGD8Z7T4byzlB79mN7GPtybRH/P722geI/OADWm1vq2lQnJDgyNqMA
V0r7ucTVKzuP0ddJH6P3wsG0UCmSPKV9tHnaMBJ8dJxoVw10WM2ZXnOUTYafxvNR
i82p/dayT3CSp01L/mqvZun474Po+xin9YFZlsIf0YOZhfQQV7AL9WQHBGbFaNSg
n2NobPBUxGcixWOZqANqHMnJHO6weqmwy9PoJxHj4dJL9kNLuQSmPB8I1lMG/Bxo
fvvkrsuDKDWtfylXBiCWt+MY+WFpJ7s/hay8L+CXiNZpb9E6ecQyxY4tzNXJOoyY
bki7r7pEXrLKTMc7o4UWKz6yCxhLM3/tF9tdGWbae7sFvylcMc9wX21b/MmuGE0q
fvY9EG/39VkuVkFmDtE8uWgmpc4Jxw+u3YZA/TpIiZLSOKbKgyomx2IUIMhcw9ym
kuHoKIH4FPaaX6wPE3D7GKWy7jHgjadz3AIFcfgPm1V69Tls358exqoQqEDTolcx
LOZZd9donmfJrxgfDRhLBYJOU0gCRcIwwNenffv7hAChvvVFQk7rzpaANmxnxpMS
qa165jbpLaPLyzcRBOKTeAzbrsWvWYMP6NItQPRM+ph8s3a1ZWv0XY1k97/05cZp
vwAOMOMd/Nl7iT1RBSEHoEqtB04kxhzvawRzjPAYMik7xDbdNFQA+m7/2Zi1YC9h
m82BNhv4gV3j+v8b7IEh6Dijk5A+3XZNH4rk4hKIENT4CLJULx22S6B0aOCaLoEX
bKCN19KjlL19RAdkQznouW1tclFmm2uYhrX9ajyfY9YLaEFkbcnV3K2twHi7RxXM
8tWrCcZ+Ck8oGDgWUINwqXp0vH0WAWdEx95P8SkXNOMJbO7TXcRa2y8wT4UtKT8d
u4PibxkNcNfPt1tYmjDykMykb/+/YVgDs7EwTgTbr7UL3b22VM3AHf17G4gWDBP2
DQTpQsrBZRSLSU9O9abzfXA4VTi02n8ZoamgKNJQ6S6PLSJ5c3yc5Bakd9Cwl1sR
wN/RSRpm0ZrpZtiT4gNGj+zRJ5rL42cjtdgCuuiARRHt1Z6T32wZ3yYOD7RXfCAZ
YmTubTkqw6OJyo9/bRjnmpeiZMQCM7NpDkOOyDt+p2NtrsWKxsmzxYg5P90f+5pe
wHx548vBMZAEjwpQ+cV4+Y/KLAzMtt0ogdVAxMVLuOo8QCHsGsk/nbR2G6LlwK3O
U7mdK+g9XOGSrQP2RWhD0mIZIArtHdQMARdfeI5Nk3vlplAwhgTSmePXg/2trJi7
c/+qtrNJGB1o/NXV18LSN6/mT8gujf5BHi5yrFcViULUqzgU0V4wBaPwuos9CaIB
8Tns1vptVgnNkhY5H4hjD4AsQNx6D9CIAiruwufz+5JbU6+8N9Ab3UjTzzHAxh7o
/A2A1TDuXY8fZx/ThSDxa3NwIYLqC+x8E12/TGNy4MEhiSH/JRn0HVro5n/ht+hQ
JIRyQ4LJj+nMix4TYOIYTOhSjjAhXB+QmMOXQWAET+dajITYeK5RWRGraCTKKl1r
6YWVpUlFOZ3+SZVg0SYojnE+Y8ylFUshhT+n941Es1Tg1EpqnOx1QOaKl/LwzDGY
/q2hU+xMVBlQehF+tSwVGAePxrmpb914lKeRASOCJ1mvRgJtnHXat0tDikm50TYL
OLROu26/Z/sGUXqfTgwiMX9YW+IoBe1xr+HZFx6rNEoBteTtFsqQEmPjqBob1U7V
0nlPtvEWBqLetKTYE3HOcx+D5som2OhnkgGDo0T7WVg0Xos3DubiN79RdiOniawg
7cswCt4ugJtmcWa+hIethBTWMbKS8aNN1G6LuZWWo4g0BQ7gzwf/AF3SUuEt/xul
d9inLyC/zzQggaQbrPdhRcUcHrPeCCpKNfTbsom7zmlSecciW9ju4mNKPvEAadN1
i6HBpra3dLLgpdUKn9IRngFz6sqa9YiNa3KYzwNqW22+Z8zYmms2a0FjQJNh8uBa
H0LntgrJsA8CNx7z9Y7bwTLojoGhtZWOcqB1h/6zI7D8EIhv30iWSa+V7T33vHuI
MdXHhB2aCNrxAqdFyG9+TazSocKNjKtcPRZOQMA0JiPB/q6PU+dWrq4hm+dxYNWs
JLfV1FrTsZY2AoB8U8ibqK2xdGs3OR5fAx1UzNMCuRyvvozgbRaQS3s1z3H816RY
wwM18Nkkodlb2cBNibXPtiE+iN0C4NkVdAa10waSaP5soxdieN2cVAojdivQtwrR
PACD4Zod14aCmlM96X1gBb4FV/ct+l/nm4fOZJUUzFhEgfRh08G/WW6U3hGYnD+g
IQwczR5XR60Mg1JcaryDlrWAWQos15mYe80IKqzhLVIkvqzY1T02XJGJL5R/52Kz
KyhXejReTJzOh/FC8VR2/nhH7gEyU2YHKNhun4uP3mcqx77LgV/K8j9kSJVXHNQr
Be6JOOx8drB07LFOxV3e+wu86u4ZsGVCSSd3EMar0ZwT69DopkJ85mMyybieCCfD
xbKMmBL3/1wdqS9OxFT76p+k1hR16rWRvf0sdsyspPl6XEcz5vDcfxzVGawUg6he
nHRKMo8YUQJY19T0SheyZt9O/EQPhOMnAZb/WhdF83Jskns4mmSHnmG4N9m1Ie/X
kojs6cZKQ/HZrvE/c7fihjl7twAfFz2YHQHiW0BAYDHNT/+my2ZtEdSuRCimFKmv
ITbQ/E7DrM2SGCmxdAvq7YIxvNwzrWGkSQhvdQKqsgd1I1EjopSUF4PDTv8aiRuW
Vur38ck756CENfzeVc3rc5cpv56/pj/p1XNTzUTOXj1MB16Mf9WMCx/sJXSjriT6
tu8bW4T5q0ypEdoIE6XFhf6tM8awhGqX41mMU+Airf4jGbCHMr4BFgIgtLDoyPBY
RGinxOQ57f7GVp0YXSYEmlLgzmKxPa4D++jQQEf9Iq9DayA58e+USIIjRbzMH+9V
LCPW+qRiDDB+qH9pWe18fi0BqBOBqZVKe1oxPq+qmvD+f94Vr/ZNM8jkr4wJFXU/
QXRxu2NO8+3fpTmTeKharIpVl0ClvMFbxE/G4FHBodk/3RBm58r/th8BLSJwdmyu
iLFEcbujOCwgaX4Je9TIbgvS/gRNQBaTxBQcSEAa91zSKGQqkl2il0tAOmMBOgQ5
cGp+tbmLrz17sc6VwkVCQNx3mjnPDs682CJcUMGoVYUS3f/AeXRSbFXZ3l0VqAwc
vAAQDD6idrfW3IohTqYad7leAqZf7Yj0NSHpnBWAWwaS/AIFRpIJS4mAnhIM98wa
GyLnSv/HU1gw6v3HyAyaaYCBY9hskXwbWKDleUDlBHFj3mAUzh905k0cpa6CLrQQ
6EJRxb1qumZdRMOoZMeG7a8l30DHC0oJNV1OkRaSW4d8/vcgA70lDyqvgOV2vRkt
whSXp4iVP/aaixCPhLpAfk/wE9G9kj5BQAiaXNgAS7QVWKMjPhgTdWF3oN9bc6ts
AzQlA3JJckztsN+IU+DhDIIyKMSAv6GGrQ9mhOpehn0VAu+XymephKsERpdIW7Y+
uvUXzHcea1sjfmBR+ZCTD/6CicprGGKSIHzCHb3Pju6n146uNnalTDWy2EEFoX5H
Z16cndmofdotBaOPXNVIenpW3fvZuZpiQ/k79KcqXNz6ziUQKy3zbRN1KqMxu5da
XhrHsTOOzRVNYj9OKY/1CKmFqUvmdMpPqzONCMLXLIXXLF7CTOr3UeVg8BOr+jVg
k+YldPnQgLIodozOE836MT8217iP/LsWUslPFOvJA34pA83/wAt8qK+BnaoRpkz2
4+FeNuYt1p76hKepfrd1hzW56Qrr2vYfaMubN4miZy6p++nKt1rA28YGJi1NIz/w
1YWECtRmG90fqTZxToGZW24a416O7iFHgrMlnDPpHj5THv0nOXZDrW7qSc8DKsxl
SetoWntIyDuZMMItl54aegW5qo/ueXqvU1H53gQnZEq0PAn3iQHUcOKHDs4XnmFi
nnMRso04mS2XS+qQeYuQnwjRm2LwzGxpEU08Zquj9ESZq8FNc6fLquNQ8niXO2wO
/YLhueWMksj+jF9AfIOxLag/BlAGp0wWPWU01YadY1f+6I55fAgGf+REPS4tScul
uti151JkkT4D9dYalaqHoAcH/kJtRuAgZUuh8NXn7EEh/hsWcDsX3sMAWvyZbRa5
3/g28Ay5UQDsKJhJHxdLN0vYMpdoTp9IxZgn3BDpRbpgdvJmSaJrEZixpsXzYP7J
xb4fyR4NYiI5jTIWv1xDuHmsmqIMMcAuxI9LjctPghygPvvQ9oCu16q014sg6aJh
BVY+SdFfr3hI6kZ0BfQHJK1YIuxNLxIyeiBO5zgYYTx0DMW+ljzKx9Mc4dPGynoC
DJsIddySr4ANCKJMu0cSVIrQ3HAzMKpYbeOp2/Efbk5nS3ZmoKKNrdbrKlBaUkDZ
R+0Pdtcak+oY/K5Xbe1DIJ7sNdLAGqv++NDmmXFhua2X58JLO5Unf9j2RDt5QDyi
fO3sl5arUYfVcfRF7c+9gDC7kU/GRKkcrJby6ghXrLMQFywtR6ixOb5LfRMcAzdA
wZ+DDJ1xbrKu6YILDPtwEvaVtn3wTeGnMPeayU7tMvNQpbWDrrMQpUaFXtLddgnQ
/EfG7rsnuHPXhDOcAVTiWvZxinkBynP2txCuFnFXEo4Uz1FKXfp1Y9YotfOiM2YK
YeC2BSI/ykTWM+WIZ3pVvK7ULq4j4/Z9KT/0b/euumv758ZRqUmYjXoh3fLzQgXT
yJLD7w1KYjlJYez1GwOZqiwxYx/9Tqi/toz2nHhuF+vIs4EvTk+u2b+c+JypwOou
gUuVNcGHb0mSf1VrGdhihPK4f3q46K0RzBZwC4D5G0FHsa+cv/XNgFWVRl2ACNA1
+BKp/WR4iw0ZiJsBtvL3wGrl/XX4b4kenTd12KCDP8dxrnyt66Q1diSA3w6GIAD1
9/nJgMmxUBHFtocC8bIbCJBi+Gf5Z4DQgEPOgjNnRb9RfZg2H8OR7l85Ei7H8ymp
wiT7P353jO+UAvD4uGecfC+uo/Hmrp5wO0BU514fbv4X6qZ4cu7t0IgASnCCKaip
m//fBXUN/htY/WtyGLSGB3zkJSu0AxLi2+Z4GqIMU/mB6fualfQen/z5C/bcpffZ
z1nXxf1RPd1wVffzLdAlijIHeRyW2sbLkailtulkNUR3i5yFLjB3hK1xx6MLPgyX
gktvbLEEL4DSvgeKLahsmttiReR/6zk8HtNdk8a82LJG3GdxFAGHlo6t3CFguv9/
ad4pmwYFPlu5SfCixTeluuZlEIN4g5YU4AWMmIKSzpLExAy7FWiWJDqBuPPFGk90
pl2hOraWba8/V+r/TWbKmXuM6uPzq5wRdUh85I/584fL7x9QDowx7G4r0fYeNajH
gB+2IqzT2pBqAuOB/o3bZuo3XnvPuGNQVIGzqB2dfkl3rkbL71PySyfBwH8/CnRU
8h91gxYDZelkMMgiBmsKl+k48EioARcwri6Pw/o2W9efbS5h4e/aOTbNvVs8QpsW
Z8dThBaTqPJ0nCfVGJG/h6X4OfXUMtdTHmW4f5lXs5q9n3nz7by1rzlIqPb3pAAm
+RRJmRo42boU2gKuY9rBUMV0NRJbje+/k+ArCea/zYgWoJ9z4g9+qfP+mmLG+Xvc
YfMY8k6S+pHYlGi1C4QzpZVf19sWKEJerGxvrb+pnItYScOk180c400fxvZbByOo
fX+k9HoqK5TDxdbfa7n+jzvCPOATe3vnLDbTCibNr7STJbC6G+CoPs8MjTG1WP+L
AOkZH9JpS0kDXkTS0GknIk5EwSUpEeECVt9T1UKxYt78psSak8hNFUHDWeYu660g
MNN4ywU38msVMJklBzSIWzUS31If5IQjnU5Xgs6HpvWTeIbpHSW7z7jToh34l1Lz
qZ2/qtUp/xU3TC/SaCrhrQhH94ngsIZXBcIVSLPvj2KFNf86UutJsWPLtXXEe8qj
y7Cy/w7tmS6DOUDoJFG5oA7TCCaTsOvU1kiOf5GEaZq4BKpdUqJtd59QlYB3jzQP
FBN2QXF3k0MoaEhB23jXorp3dhfYXSgMpO/2LjQApzKvVVZxcaqLENPPf9P58Opm
hrvk9uOgflTnC/KCJl+DxcbAhiEwdZvYqP+dbX/9ErzuUz4CaZuYQyrgzrb48iAS
RuIX5b70rgRGXP5Ovvam5LNQiFwpg9zGq8n7ueB/8apfAQ6I5qIlIDZxdN9XhUUk
yIpI3BuLOV/YvMSDcbXBwjrTHjl71r9yqb1hxSWPypZXmHveED13xbgQb5Sn2RUb
r9Ik3cgTgO3J8kjmi2nwnbUjCJLKZ4JuWWokdK0ADLGk2dfaqthseXrDb3G2qL9c
niYUoW1oLH4CWuKJ6DpxI5NN2mdIOGvEnG8nbjJEMrgGj01E5ZcfMoKtpMT4lXyU
Hyd83yhn12wfsuCYiRBrf7AHybc7kDGtzjpQXMQdFLFzhEj/ujFO4kDkIEQVsQMQ
lElo+omMKQ0cJ5+7lFrly1ijcV5jjUT25mMOaAW7dLIb/4U7TB72RdKD/NEDxddI
aQK5mFWfmsvIuQ3+iwZ5nWLJQCu3m4lhEbwsHWFSm+KHSyTwcMZPZBrX4LlxvbuE
5zQmsmyCVHIwwhU/D5C/ISAn77jOvTRI9+QbL2tXoXF6o9oBKFEPbDbotRRnVs34
gU+qJNizdbM6eVs1n19F+p+R+IJeGK4N49P6TqYZmiCsQNJgAdCcB9nz0xlV3qbE
2HcA8klWo3w/T5gZkG7JHUxhyUeHxu/zvAF/MjqKRs2+zEOCzjBauUppz4PsZ1qQ
x4ZuPb0g5Y00hdTXn85QATdtCCfMOnt/zQEGogDBX/z0OVeQ2qSXQc/I15PUz3nF
+QxMmyA4yJci0SbmBAEUOgW2sR1ITDZL6iudqNWRfXzVh/NHrHbcch/plUhoqp6D
EJPcjrPf/NKwHlsz6pd1cPyrs87biM0qZzZwkSAnLDmKSmj8WE3IRG0/h1pYVYoG
UPimdTqe52KA5RDGATVr9yE7vTylXx5Ioh199QtjlS++IYDOQAiMYjTF8VZgbUDB
nDQMksfXCXVoOfWgPgrTjvPktlq/542HKhP8abu5/2F5399sS0h0WCLpEVJowR/c
M/dHxw2kU1R+chMkEGpMy1iJPKGElN4fJg+lJgpnQ2Ms1+vLt102ZpQLkO7OjRvk
/i9A2ntdz6whiCfH9Y0y9RxQMH1RxIr5vjasKeOxW3Xw7Cnfr9sxvyYPwCmvPKcG
qhoNHZT31+5xDauW+/Cm1lrqJuYaUMuMdX9fyoa+HmkFLRFHlSV1YlJTKgyV4q1k
0GaJPizRdN1yhgu1D7UhlaKEyNwdZFcylCK/ZDgsrz7M38Lh2i2RA1j3tWYzpeU8
G1J1j5Pnn3j9tc4sYgS6HhiS5MWdc5RPL2DrdFUrqNrbCB7lEykgMEjrJsnDkfXF
lrnAvJ9soS09eKgAPJsAwhf7NEc3+C8qXq2cWf6ZLJtoWXqjb4imiTRzsa7Oh9Hg
TfmeyjOoaJt5ZPPzT0N2hIw/siTP3Aj8PwizNv/o38U26CbshXhwZIeiHJTMbpI5
vhOIpBjURfh7e53XJKoiHrVkcc9hLmSSQnqwd5NniuV/UCMIGCYUdwx73o7Qe+fs
uXvMppN3aMSaVSFAhvQpcLIqNxDjsT0FRyZxTMcwwDdc34liTQFpmKrrs5Ppta9s
bqhHQr9mwOR01oRU1t9U11bnyNDU1GSuDGryNnyXd6O2b4FqwUfHwPc/DJforGk2
oL5TsDwO360A0V9gpOdFgErKXmA0GBdYVFovV3PTlb9/kKnJeSddKlMsLNUhuvY6
Vt2wdjGVX7kerXZv/S0Afw6pRBLKEfZcTQu/BfQDKK7P1x1Bs70ZRw8Tkr6/YSei
TQu5g/tFZ4P9olVbWK0GPUMv6acemqazBvkRI3AODxlnhPdB94xK7tndH6UuSS9P
klI3dx1giPVFWu5MJpnBND8tbMIfXv1zoZUtHR7AfmzFDdWaj7Dyd4UWGlHeJ2gY
bTFbmNxPCzPFicJRQ/g1VXhDIgkLYP/PKjfNZQLBQ02Sc+YZH3QZLi+jf3T9GWOF
sdIrJr2+AoOBnbaKnqbPZMHiDfA1T6igtseQZAtR23K9W+Sbi2VJ/5cnnwRXV0TN
RXDn8HGZ/FZqxxgUH+3urjJypgH/FGoyBNT8eTJMwk8tOFQcvbrLC4VKrW84q2Yh
siMbsrmgC1yyoyMMwUjOturctyvWqM42m+v9Rf+igk5JFU0jGDILIgrxyIbfnH1t
3WSXeMWZ9VPePjB8dx5Y3asX0EN/70VC3nLW2nOeO4msTjrQ0bosH8gFRX0xS666
YlAemkNrT1TrPDy6poZZvEeOTW5ERL8yLPr68xwcw9N1tHwGQ31E5gS6Ze4y//C+
hFtKtFHSyRzdq6hJUT5Pl7KlzlZLrJPmiNs1LkuSZtBkxspzPm33kDhtVn19Zmqo
8hOmGpzM8v1V2N2ce4/47Lm0zQbQwE08pjg8Ps9QfEX8DTGxPfTA7ccq/x0X03jJ
XZ93NzhtGNLAFuMv2QGFc5AlqwArlX6bQsEcKR8vatZjsGvfUU3/gEF4cCW2g7tl
qBlZzI32UwfR9WgojhHo1VCgW18hWdN3q95IHMxRMUnX/2IU5nw1sSrqgQIzSzUo
AbLTWcbzU7KArG6b3lB2krPN4bwHpP54gj+q/1XDceSr/q1cVYM3QTiiM2ifS5jR
dSxGrDisr1iWrZ7v3lmfCC2AUFykq0L8YN8cdTn4XxHzOL1HBxBYdp5aP2DYMXxC
3umpalv5rs0xItFytaYLFcAKvB+MQLTfrfE+VmjgZzAe3B7OQVS8E5JR/qsfMSH/
giNaEAawTDfyeSZqLSpSUKN/aub3FkTT4d7lBahx+/Vz+LXiktIWsC7easdfJWLX
ubk3pbyKnXUOTZQXplUAQIfF/NgpO2RPhpGTy8YYovkG9zbvKScLkvHBYg6Z/jf7
tIktkJ/mS79GXXGPZFAexDRX95XaxAIuJgQryT8cHOX6m9lVw8GBumXvbipgsKZL
VnnX27hFnsVvXC4a01IDjdmumjX7SrV7n6DQ+pT/noXEQMMmzuaEtLNS/aAmUPy4
Px0XBC2z/A19Wxg71gpAmm9bqw6j8CtiMONrFCLTWVRlFAkt/P/BOgqrkiFQiSSl
YYcYRdHE/P0ou6CrRGKYEVaKMyTGfa2BqXgMqB46LDmIDycliQ97eTdbdWvAKEbf
ogkUPNVNliGlAHRfa41fEg7VNUVjcZjILpeer5WicdtRyGhF5oBKeRw3tQNDza5s
hfcQTfOUc0r70YMNobE9F91wgHuvMFG5RdGFHjY4Zq3oGU76WCnE72nM1ISp2PsT
ozG/4e6NDUTwx5/phEw8n0o1QK4PnUpseFrJAEWnaLxgXqwZbiYPw3k27sSBf2KM
83b78gsf1EPdhrRPck6WNZw3D3jggGvYUl2txOuSbcAGp3z6m6QCFL5avK1GWPYo
ky0uS/rSC+KJqQA9Xc2z9H6t+wyO4PnMIhOIbHJEWGMDS52Pfu86p8StuacvSr3M
z+t1KbLFc+bdYC7E486rN/IW1VAjVpRF+Y3Qib/34P+Ww+ufzY/fK/GAz9qtByPh
mjTDcUaNrn1m19kfKpBMQpzuEWZbWGgCA9LYc8t6lA1BulPuY34XQv7KGFfzswmt
FaLXivht3dH6GiMNv+DcXenSD2E69oO6Q2wxPaL9KADuS4FdMLOeB02f7DjoIGPR
aNfD1ojuTd5tpsDrB4mUfyKfCSGhdhubh65lv+1d1ZUh91XZyAzrSnrRL8ELlAeQ
4+H32sFLBk4hnBMAbatgDWp+mri3FS/a87gFFu5HQbG5IUM0G6D7LuoJBKs5Zu2B
Pb4ZxKHMvhB0r0wcyDFd1dHlf9oHpFcwhzwwb9x/hCT6kiXe+Imo6L3D5SqLpVa7
S6UJ/DDOxxo3vBZLFhd7MQFOS9JQJnAfQ52k1KjsyU+UuzwlWIOp7VugxA+TS1ib
txPHZHDb+NM5jMkMZnnnLco0v1gcb15KTMZ/4xWGqw66y/c6N/e5TJ9XNiVEGxLS
5yc0xsOg21rDluPaG49iCMtCWus44umKdkk/SVEgklQ85Pg70OcwV3K6hHnSvC8E
y/E+SuXVlWuWtqskFbOFz8hEQtAfltTJtem9PUdWNRKUeYdBQkKcLkJwo+6dmlRl
GOZBFgHX3EgJRwc5mC7v+8m906ZaJKjMl6o3eCnyTO9a9Hzs6Qh8KeIKhO5CoqLn
nEZY4GutB2Pf2vJbj7Y8dOqSj5JXv/7Xa2QOVfoq1Pj9dYniE87vMGNSZ6I6qHLO
lCe/EmW81PftrgbW7QewLRxK9qGi0dFfekYFJ+qpNE86XdoecZHDpcAmKp/w5uIr
0Q99W+RukvI9hxScHOMZn+sLcL9sypDT6qgmgwu1oTD3IqZmGzFS4UY8GrlZHywM
f8ecIYa/du9dJ2JE761csAby+Qzw6ZGjDV+l37oykwD7fQFgvRzCVfu9OnvUcydm
hCC1piG3ZcJwFZtE2xGcqEa021PsV4st1o1bIQNFm5nn2lyIUmdjV2v8ja5qAYvc
x2Aqpph+X4TBDNyYTVLkRTUvdbhD2mFUd6EopcfUhYY1r3JmDQYFSYfmqY/dzrF1
kN/yGH7tu12EGiX/lvdCDH9tE1FAexGfWUPITwxcTs+pp9xZ68RiRVIRsqwmQZkw
zAoIBlTiEHhoODMuBRqptFhJta/RNLO7S1t7ve11mGnTPRSGi6h+6BZU5tJ+y3DS
uG7l5io66VraiYF6+3YUkFAQu1pXzaiHpmzHhDBDQ0PwkWzXcxiDMMQXa74mDrhh
DyKK7XWaWvLiiCxXKDDlM1IEPKoU/Ta+mshhRoSl7TTfKVpuzgW/MIvtMfnOMW5p
C6Ir4GMN6v1i4ihNjsGJzEI6hboJuyMBpcHXnZdCEDqucRKBqR/y6lB3psLuGqA5
nQS3erHonPZ5rWGNJrZDxvcJjaV5IjFyoYULz1f9l14Hyhlu6CyWmYBmkBZzk2ZZ
6mlgXOnbBPl9TK2KE7VZ7PnNRQOZ8trXAdsaCkeddYteT9NhbpZirmO8RB4AArEO
Aw+xBcBOM1V26Q/rx6B98Dd5V67jLP7ex+TarUPBelqgZxbXyWEiPxZMPjvkfZmg
W7KIK3WFmLPi9itG7lDd8F4n7saO9ck16ADRnuAZ8LTboCi/SOuzehxiLJ845AU/
hwH9d+Y62XIw1ZofEy2fBy4ipFDEbIkh8jKFlCao/KrUQcl71n96FC9uEb9AW/us
EpalyIMvVwJxCWJ3WF8q4wBvqN7kBEj3ghEl8crFZvWf+6D2g6qqu2TR8fhD9v76
cyet/FsKLZUJ43Rwitl6bSuP2a+k5dCpEm0fyANw8H45b1FGCqd8pYffgB+fN1DQ
pNskNdcKM5qLgYQUhkIkQApKcN16Fi02qxKdL8R2pyOzrRt0VRtuIzvGmAHNQHW+
49IY+RclR3rQa7IDk59Sy9YFs19vsSygXvuFs1e/f8qedOoB/sVBSz2FLkQPFMlx
lnbD3sKmUwT/Le0n5Of70rB17y5qKjYhGMJIC4vubE26JsVSD3kiwe+aRFmMYPHp
M/t9BrrhdXBO/+D5/H9jKgj0AP4gE2P42H/SYRqJ0Iu3KAkN2mF+DNSyKDt+uYhv
sejBRS+yxJ8LawBOd3RH5bAsQPjTYFY+H//XLMcq++iN2ds3HaNRzDy0QwF/L0FB
fCjEW9xeb+8huYDLOPTCquzjB+SXxqVsNmB96cEbDWuzLoBjFY6qKeET7Zw/nVAK
xhfMILKrQV5ZLemp5+Kouqt3+dGab1kCVYTmM1kB6BZhy3eIdXZAkVvJ11t2LGJb
OEIfO2dQ05i2E6bjc/xfeF30dp5cmTuNcpOgmlIdGipx4N2ej3ib1JZ1nMot3eoG
m8iyoCORcK8GybuK75OrKUBAxgoSgei3mkLaFlTl7Z8H4bpbJETwRtI15/L1HcMP
JtY9OqFdlbB4SxUYTNhArbNbN7YQbKJl71piROt36KI1uhpG9T+dKmjcU/Y8xqBn
RFeKKP/LEANtFlR/HArs6bt2w8L/I8BtIKMdhiouSW7QC874CNSJseHs1XUcudLj
0KEnnGoIkFaP+VXiNXib/nJDoHXd3aIbloGLtjGrmp52SbS6pPqJmhKy5J7Cds1z
eFsPbueE7taNnc88Wx8ffUyXO7K3CqWs94hSQoaWcLHq0o9pNDfJGhtbYlpeMpCo
UGBW8uRgO8yAB4+npJ6jKb50lrFHKZbOPdGu6/LFSWc050TXwyWjo9IPQcH9WPls
n/Ebv5jhemO3NRuy8EVEnegqbalICaHahuTYiWz/QYcSflyLWvPdDwl/zRGDI+0q
sS6pPoWjkjFf4sSFdOgryQX53R65T4Laaarp63kC363EkPgtLCJ8uuE06koQGtID
jdlgWPkg/CcexXj5JqsKfgojN27DExf3nQ/empMU6dDGsI8GW+MHSqZGnWYr5xcm
EZWv+dCaOPgRuNlJRKLISEkn2BrvGFwODKvnudRnh0dZVWaN/veAgFSLWUVlNqbq
29m7jCmm4g0/049EDxSPzcga8v5po9p1c2q7zo92lPmyOJQTwHljXlA5+UsV8Wvr
Xoe9RU6suJN2+mZtSdgp5j3pCTX8bs0I/ocvdzqnuLqiMpSxve0Vhw+VELeeNdsU
pdKZmEOOmAgR8FIJ5vLvm8np2c6eqKOQvnVugiC3SB32qMFoIlNdcUqSVRjQqc6O
GvFvUs0pOVtm8qB2k9PcZ3Y6hXQTfSjfeWS/TqE3DjIpcMLYHhC2VlrmgZHq3BsV
trh9rofT1zp9Zk0PMuqyuvS6f0c3ftV0amDSXRbXz4dg+6mdDCyApY81L0Sc+/NS
OJw/VWtlBOOwH/tiJ4ed6SqHnWDZQzgat6/UOBwQYPFr93ab1NdjekEcwkUvUP7d
JwHveFDpgqc7j70yfN57+UrXaDqvaH4jKSL9v/X4nqOyLYiWQs5ghiKdGFRiJR7g
DtbAaiMf6jDBDMKHPno+Jr8a5v+9270bq4Yyjh4CgpwJPxHqPkUw4ehOeUHjRYX0
hay0575x7pLD4pec9eWpg36yhwR7BnjVrw49yD7ocC/uAwn+c5PnUnGfhgQelz32
ddM5L4R7RUN895sTTujMMJ0j8SgmG9E1ICqGFa4hMvfiqNXyJPZZwyVomrdVBAtN
8xDQ12HL/srtXiodx3pj60vQsO+XzIDzpHoNOVtWW/PLJUK7kSX0zOQbHSy6n9oh
0puGVqLETtszzWp6eyffm6NLTIww/2qC9hX7DVhnNQGjmZhayGefeq2Zufjwv0fh
ek19uvb0rwSJI0qKOWBVs0RwZEO/r3kZz8kWccksOs7fT9Q9I31iMIGS5iBWAJdy
6jFIzlxn4JNQV1GfPuSghhvDiZhETAZlBiwPHnsoOke31TLB35xJYov0QlBy99mZ
iMNoWBcnaK+6QMQ/YWDUkBXERJnkFpSLuMUZwKUbKf58MzeoWaT3L5f06dGNhEHI
K60bwgjNabdDU6QT6iwZV7M7ij3AN9i8QpSZwPT+6e3XG2PDAWX8ygFXljqEyNzA
bllwnmGKP1f1rMqar6ihsT0RgnlQhupqvs/9Qathet9P88jOMAp3UgiH5cA0wWv0
04dasLzoXS6oC5hIgN3C9qYWb4xfQDVcrm64QEV9WJfYKk1IsFHP071rgpWEmLWG
JHISNucwTqKj+CzQT92kgxtjjZDwH84GvwpKF1Vql5h9KUn0Xo5GmCs+1k0bb4z/
ejWpO+kAM3MIe3oaNUY0sGGFXNHz/ma4qQUWeF1AuA3LUCyqOBKl5C7lPSeH5dBF
dB550RRoswLH2mElEP7HsIGWSKp3uOvEsy/3Ij/O+xOGEeqWikmN0AaUBHg1dafg
aWuUNPbakC5b5kD5N7XHs62OUPAdtPdwpHj4fC8KU+hn0ZFcy65GUI0feIMguJlk
LeKWJas54lAdtraNcVbcEWsUrATjsYe+4+R9d4faiwMO0gSPapSToaBgpicjjvyV
szHImozwyqq0ru2wORSnMZH10yhMHovM4RQtMmJU9c89ihOLFJ6PhrYjduT7J0j5
p0Zrc88JPOVJuUuEKtk1+Yzkc/VVcaN8gEmFXgfXolUVTMGbWT0YaQFIGXCHKLPu
CuI8In1VGT6XSI3++pVPYCPk/6Exy4yHZQ8doSlhBkVKhY6DDxFrNCF+7R5djdhl
/ZqdU2QqKLsuzo8kZS6yxKIqCX0Xr+kmWJczwrAoX6HUZGbCJb7U/XVgFXrxGzpJ
HE3eSuZ6FPECeHsN/Um4pIwsUnzA34rpvIgCBDEWEc+kwTUIUeXewbbW7oYt5CwQ
r8MPi3STA8PyBgK0AYpxGe0TanP+3hw1mqmGlFWSw6TDv8FXu3U4nbDnKVdHK7mK
M5ag+gcQG+ngab2uU6t7yeKwu0Q6mEqcGQZV7YnWJM7axuZQ2MAbyaNbCkPeVckB
+QRzby7kKN98hjpw+eK6SH3kUALbG9auz2ub+JvVEwEQ3Ruri/R8Qcs6Vp5nS54A
s5aRJk1xVRhfxjIeiH81UK2VJPW4FomJo9WXRtNKxJI0RD7wkFONLGMuQDoERUla
OxO+7Usj36W7Slwx50hp2pC2kLudmthc6CzDFrYAtrWw4riCyxeYTPmGr1seSy6S
uMw3ds5N0shFTrKV6evWMzW9XwrYMgGNtYdxL1DAu2fyCmmGYzLh8+OIZ8oz9I5A
/pPkCtOsfsz+Qdqd//9ylLYs4stT/4wAzJzwp786IxNY3Adap0Iv/6hFqnIwYLYB
Q6siwP28r8ZUXj/V/Y8GqeuVvLkpatpqyZ02bCNkLMG/UL6aoHYMU14iuyuMzPLp
I5QXPPZ4LVK0XrUVYf3jbKgfm4Rki/UBZW74hiVxUSklFH7/mTsZ6SfG7s3qSUil
bxIYoEJ61g54ZHsF44K+TBeXirk06Lm8XafoULvoIlaFgx+cclFcO4WRGcMaACgW
u6AiednPm/NLXzzGuLp9YxZRLb4vNrzjQ+qNu+J4ykjk9K1psfDY/YwJzq3DH2GG
2NW+661vHC0QEhhhKZ9AIUpQY26V/1OKy3F07gNd1oq2ehCb5UPi2eLlf+fKvWHr
KMj+yaUFQve03UlaCf3BurYPx+OdT1uHlroG5hlbtIcSxxuk5isliE2xM3J7MOO/
2hbdalRMrRRWEYP+NbfxmWzSRVrsYX3C2ocL87i9e+88KkwTNJykR3ZEph0S1htM
56Gl/baymJii4JIVeum2S61hLPzL1Pdy7YMNbpDEo/xuZi18szVOCkH9ubNFsNa+
IrxtoBVHBji8JUpYLxc0Z9D/CRPBkez3CI657J/WjGYEkoV+JEAAfQaPlSQ4s39a
sQ8sH9zj97A40SbIyBmr49PR+PTI+Ag4+HPBtG1gz6UXK5rTV4lb2HFzqjZ4+2EB
DwX/3A8uXwFbWJ4dz4tgD1x789dAWF4b6wkLCVFxjThycfThUFqQisOqsno3/Fd/
ayMnoRJpwxWiHm1IPz4BKXA2en+mrQ/RJTEkhLCq+HxrJs57jz5D2QGbChFJvuIn
kqg6NzJV/Awt/uwyaNfHuKaYNxdHzCxB9/gGhyicCRl6dHutb3ycMYFyZGZ+siBI
3Fm/4rINOyb0+HuulMy0CsMZuo+H7airsKMmJ3C4z9jGDlXQsaY33A1fOEtLceK7
MqCzzYO3vyqkIBNZxPpMXSR+bPa5TLB8cJ89ArwYWA/9Pj946yBimqwkFleJYs3X
VHh6bfnDu8gVEWWmarWkWebFupAFxtqnPtVyCUZc60+wbhvj2mSUHfC4ft0EaOR+
6tBZHEguct3wlGTafU+mAofnNvIgcrUcVrh7v3sgLS/nC15NSHORAB/m0yW6OpOT
ayyZiFKnSV12KgR/E8jPeqJWiu+fT9dM9pk/+0GQIDhapttleUYPX3UC/cB4y2XI
zMP4xoL33nt+jkQOC0l5UpUHBpRww51pjZNiqkQNpU0pFeHkhXb7GwEcf5pGnKUS
NwEsaGlr3znqBoiOW6OE1nSJQVEp3Aqi6LAQrsXhNhkmw/sSX53avkF88XFHIgxY
SkDa+8G6XTkVuQW+Y6P4qvc+ImKGTHQhTud39O4Ye27eHuh6NDAbvliUeL6nWFHH
Dmqb++tZJzfcsULVNTSEx5R9WSow8qu/fpSSFsprxEcU3IryvnS+gXhhCcKRJEZW
JbeFDQhJT2lGcgRWATQIQ7tkOWc2MKff0j4MpHTFMXaLksTQzY3s94wQo2bA/XpW
++inCqgUkIVvqsKfFpiWaLBrwprV953IikQXY+2nSzYtRpq/es6LmHcw5AeyeNqR
lXGekobXWzipdhr/IlkcDIUVLmQnsSckHH5QGG0FmTJ14lNx7zt7It/rN5wFBFjb
soanHdK8BthzuGArPKprgmd0eddbMHysAsS88/i2AxuWtZALlfP4+QOxRQAf4WsH
NehK6zG5Utvsukqgf7i34C+ODrcWYrE1cA7o+0n2GY+yaqV/5Fnoj3gnZWS3g71+
Em+24aYPPIBGtVCv4VN2LSDJnSgoOhyc8cTb+mvqne9v9gMem/e15Ms2ei9xCpj6
D6Kl8cf5pgrzmh+Jzvrq9Tpwb35vtFLibGkIxaS+7TUyhfAQGiwGHtNstA0sji+6
rYxTrAVF3KvtW5OnJq4cjeUtE4uy4PqYC3+nAumcZkvpy6kMyYb174RafyjltpCZ
cXRQRrwC4zeP6yUxD4lxde0PqcRprgYv/eBkxDN+/TW24/tYSQJSqVBrkKtI2N3o
LnTCJGMagYRzeHmyYcqiAjcKFDoPxruEd09wEc7L4Pb6BhDp1mXwziFn7x7b+p6F
HkPi36iI7vqs39Z/YdHRFZknY6x52+ehlOXaG0zWAZjY3hiq9gU8CSNIvPHe7DmL
/z5ccbgYhc3Vz8H5pomANOsEk70NVSC6biWc6kSNfvjc2etrsIysO7A712RsG1TQ
aQP81FPqRyXH17rmeUrG9RrfTgJ9mMkXlsjiwVjno/t71x7Hk7C3nISUMBbooB6z
5UiwaM+JOIzqMmZcB/pA1UHYNKDjVxl00D7IiwsAltVlOVvX/o1+jUaNdjIzC8Vp
v9ah8E8/yLz2hukDTPYc2vU6DDb2/EW+eugLHHnVElWPpGFw3WaBEMMmKOEszEHR
39GoyZiy7CPOf2/gtCdx41oB/xh6MPOrZJs/bDU5vm2H7unAsUfwZnRSvvbq8oPR
dTU7yOVLXf+hD0UeVDA+7YKBiVatTuo+qae8e3ap3qkGGsFpBJH00LoB4IN/xDk+
lUZgRtElMB8+MrSw8/ZrDd5Twoti06uJnSc0NN8NWlEPA3om2ViyMLHgfFLIihd9
KfsW16ThbgvGVvZW87IueDcssqMJhnL1pSO+Ptp54eW1zYgqyRx1dqz91qxaRQK6
Wnd7dULVwzr+VtwbAEDQ13E3KFHyoJ8fz0wDaZpX+V6tKb8FzDxcATb3Sfp2baNY
q/2cfHadDQ2M/igsS7BjTLb7IYTnYCQaT+iODhu9X8t3Qn0bhbrtffVU02DKQYYt
qojGVHH8hTbNhZcj715yCGq3qGrmrlUDSXJrDTRZrrIVSYa+cWEFELKamoHICnyK
3JlgKXMX7XnuGuB7rm8jIjgHagi1XWIkK2JfCNTvAtj60VZ9f+4/tqYNYr8wyJ4c
qe8fWk1quC7kg7R/s6qKvWjNfRQHx+hUpCtr5SVnV5wzqI3eCdgUDGaAYdxtOgLb
tpvpUcoY2qNWiPzmPlQ6Svog/hrqkHULBxYs20AVQC4YM54/5BZvxmXOgVN0wErs
SEXFhaCXSOh0JAHL319gHgCAtx5Nx958FxHeCPQpfb6YJNYoraYLNoKvZdn71fEq
UJYkzxEWs/U/DRa9J4SZIXZVoPL8Jcb3sNzWNJxylLMQJxNY6IRpYx8Pij8rKGps
PjV1NmLut2GErTY22f41i8ENptOBpyZLoXpdOqt5F/64aiRenQCcMpW/EkKjucJF
elyNuVkbmJviJOxRzCYSWG9PvjvhOeucNPfsvzxmMDgm2d1LG5g2Zud6bC87Xs+t
K7YpYuIWAlHcW1aYDu9cJw8mnMS0OudiSsFnQXWxH5XwKSVKWnNVawRZodkmvgt6
2jtJFjDeWEKZmUiC7MLN7eZZ5x9MknmtzMQEefY/1yJFIK6CGpvSfh3loTUBDpCt
CJ74qJ5dK0cFBQMkPFichRPU4KyKkVm/rR4cea64mT8j5ZiXELtQRjecXFMHUKtz
+/mHUKVBk03WtnI2eFFBXvyl60/5ktw720rHK/R3Wo4Eo+0b4TnyLggWh6pXKkH5
Ax2otBolhcN4ZCXT4UBvc/qI12YdlKb2zaRvqF03eg/IUFhQmoaqxChO1A/J4ZMe
LjQTadNyQHGxpZ1D9v+GxOvptJKYT79XQSLKreeW/3/6m9VKk0IPVpdBSMOohDnd
sJ0WgNTbgzrnttYeTChvpd08g8oKwSG7I5jcJLLJ3OpN7sEfvubcXtb1iRkAovkq
8j5RMEC87u/Gi2/JKSvCWFCZ5knoJ7edmlOraNGIftebP9SVq+EJFSyW7i+sg6Fb
guMJVOb3CrWxvxIRvKYXNQFOpXWYqlZNYYbuxapVXvZfZ/WNbScVrto+uYgO/VLR
Gc2cP8SDuEN9ee0AS4yOGtKD8BC/JrkE/CMx5PT75sSUpw8H5/JGEhUqujFvS2mc
PxQBt7QvBxtC8RcP7+TKP7F3jYyKeSngT9nwNDEXjoZMJ98BDmhTjjd2+pgkDf+Z
wKFfCxIHytZUk/FSasFBHJudiGbYPY7MVdXl/HgKWgvfoE5+DDm6wizhXsujda0s
wfIcJdlGsWFqiEyLSb9XEVTILw33IZdbnl+OOG0/DHpx9c1xbLCissRAZsunLyBM
/PxSb10qKb5tFm8zLli2w5q6Vjxac5g4xInuQFkHDlyXbv9PPNN7qUTi7aOIkfYq
1EU/7CzUhfsgBK1VqpVnk5oQxz0bqBadSB2E/0UmS09RjnOsKi77SziutlR5Ns1B
zXlySV6Nx9pKlax4bJHs/RLPL3cDvibpqRhsI9nMNUAek1dTRHy5MYueRbzPbN0f
+g95zxwLi3dwGnUHzSjdgVeCEtZQNRFlcrRAURX6CgxGuaM3s13+m1YiDj76EScA
wODNdG7w7aawCFXpD0C//VztM3o3yY2Rb7ohFPgwR+Fsq6N2G3XURvt+/35xZwZp
tjzE1r0s0H1ID22L3oteO4lGvb6yT4MyiGEh1WuInKsz3EO33rN8sQHVBAUTSRyL
B/WVKZVfDwf7pdh5Bpg68LjfjNUL500Y7I7YjgWLxEx4n9VAgM+tvMade7/nqtLY
6l+3OfqAhmIINoJX+Wzy+/YD6Hev2L12I1vRUsIF4EBaPpPo0AvgomwQvgTMyqnl
Ho3WpQaDW+TShp11cFhjpCUEQH35+BbiaKucDGHu2rO4JzyRR1L/SK21nlfLZRv8
Hag135wt7YkAaGYBqar5VhCQ9HuRPtV8TEaHBGb7qp7bMBj2/26GFv1e3C5l24lJ
7bsHXnxu8+0zKTfEy/sCfPCjnFHXySzdgUqcjiHYmJqckBVEpfgVin30yrLELQvk
RxaRYBqy6kW1m/Sym9Pxb4SvctKcebHOj0WVc6UgXi88K0lCmJrbdWc0MTOGkYVo
wxM/7lZ5Ue+a9olgAI2ZD/yXApTHnUIPk4Msq7BIuvdFQvzSYsFbsVM8UO44M//E
tJPzFvP+uV6lmTSQxyDNWUzeKN4tE0Z6D/ECYU5kP+VHV5ebQeuLUvzPfYAalOji
sMTkwnqXZ3SxESdS6/0ZUQJKOhG3NuZFR7k0cOtK+4Dj975hBNw3nmjztM5yj500
mF6MNDf0D7hoqweQNN1NgM+121SssUS3IxK71lkuAVQNeD23JG/YtqlKNI9rcV5I
m5AXX80th+P7J8MZBDeV7WAhT9lTKMqy0un5l5K2EUdtNx0vJIJvhGPoImhqhmeY
JYGBMDgcO7LoKwTXNBjPgfozRLZshrFKYYtyVEmGezrKr9sc6OtBBPKAZlF2ibFR
PZvgVO5AYs9sW4ul3tcxQlQKv7NZn+E89HN7fRl8CCXwvznQ0mD43aq9PQkhJQ6j
qd3AzPVrdPru8PwL+JCviKWFZrE8Oc0o5clMsMJ0MPjHe2sV86NPJfBup67aD5NE
ibhgq+BZocI40Nb+W2Ui7F65ol69D2T/TbVMCh2bltWjPqxnWOGvmbySmoIoULcD
iQpAcUN21JppqwZYa4+s9EqLMa/mX1Zds3J2I4nH6eh8buJomNmIHuf5Uv6fWgbj
tn4kxYU3TAqa+6vG7TavA9SHzCwsu5xDXiMDxdo9E4nMnjW6PxxclFfxz7c8Hz5w
VkwGiAIVZCggNzGV59FiR3NEs0xcdLSnzmiwqjFCNuUxWCy+Fev33oGLmreusDwo
qmpf0EGoNuPWwjYghQQTH8Kgtv2avIjhbOpxn9JzrnKM0Ezarv8tFBJZru+CsVLe
/NQAHqMO3cLzg1+ZGrJgQe3AOqngq218Hzhl/xRM+R/ZqxC4cpyw7bbWaqI/05OP
dqnf34ElYe6HC+SiNtr867h4G95d3PCIgx69L+ZifafW3gTxduEpmI5+833LJOTA
QsLSiSvRfx5fRLv1tDcOZkaWE9FwAAmsLJ/jothsHW7EwJA78DieCMj86aU3ehGk
hHprIXF1SSKZt5L+X4VVAd8u+KyvzGo5qqSIqwnhJbd+gNJLxER4YV/SE04ZF20x
hezSG2pEQv2Rjjp2DU4OiF283F3wPoXJL/SSUYvPrZ2Bi2EnE0SlUoUyJol8VxIn
/UB7ukE70L9SqI+bSUpewVLba+pLGBvmkZu3I4ONn5GgOgM3AjF1Bvnf7DCd/rg3
rX8fBfq2lNdwkiVo9SnGJCKjrqr4QA9gxbgOtHNPQZ4ANJqEUBb7DTgKrQ3uOwqf
A4omb32jbNnFmbQ8AyONAV779usExwcxyc7ABfj6qd0TRHB7x5Yss1lWArci+zxn
nGfOrOZTu5XTp4O+CkqF0RaXhTIT3YnI0e/jOUz+qWBe+opuHokFoAsJhDdasFRm
cGvtn7BGTR7AEDLHR8KuHUkPxKvARCmmAaU4rw1zfeSHR+HPWcdd980OpJbKP+lx
NDmnrVh2zTIlsRMzmi7Yq3iKB+pLNg80+2amCs3vu6cw0dOpSo52r08hKtMe4EQc
Ac+6oER1CXoaNGsLmdREgMOMTpdh/2z0uqIgdNoQ/RLJ0Ftk4bTDb03Lm7ICNlYT
YifyyNWKIx7gr3jUMS3HJPrRZjAAYKFBBqXYy0YcE6kHASee+udhSgnUWgHU3mXA
YsGve9YDhyzY6EuncvjXmyPp2dlEKM74zaetMawW9ui00Knfn8QlsJB4P5aXkGNq
Rqai5YYszvfJoVUkyXfpw1/tAOm8RhDA1p9E3gvWwIIjE9vLRbbBSUKCCFx2XANI
icIBjxQKsFvxjhS73QGpI7G4qyBEfyixYnlrLwgOi6EdQ7MD/yo3eoq02RaSLvEl
pUDW3O3LLwrqBbmJGPWl9o0z/o/yrhcpCWyfX6eNDjq1CgEoWgWR+kuNyNkZfSWQ
XFnZLl0RuQPiXP0zNCM9ExgL+Cgmr/2rZpgnSEHCmoiXKaRBY1th3zAVhRYTWCfQ
n5Og7GzWtvPq8ltrebm1mFNmbSBZ5woBZRA6WhQ+phSiTAQdydFesyJP6BGCaefA
ytRSKH7PmoKhX+7cGB3OWqLTXsyyWbvNTNUy6U71ewjzfYDGoQcvqtHnSDrEbGI4
WHEYrK869VRzu/0oTuYR0VhML7qAFZDHrPUO1eFA87pnRuJiWPmtbcF8krQwzI2i
QfBIGof+OJSz8wa2Emosi087/vXGv4RXQk57UMiZuoGlQVXW2YUXrYxiiU6IpYv+
7CcPZLO4HgEf96NYggEWmpSJVB/JJZ/qbNHyTqqcAaZVwCwuClOdhnwpczzQpIMy
dQc4TjpQdbsQjLHjvXkMKMI4+ewYgXuAYwLBLPwg9a3nijYQ39yBgFNnCidpBDly
OlxAXJLDPJHnYXHn5L/w47MGyEoTZafqMFoK3/FFa+DX4XyaajcYZsN9/yIGMnp5
XkvfYWWvrCfd8nFBHfBXGlysyO0Zo9uN6PEvyPl6TwtEJkbiR43OFdpd97FAUxOA
s5dAO+vCyLcvOH2ib2hoxMo+BDTACCLjgPB3f2XE+OhJ9GNXdtD/IMze6rsof5ai
uZ8WiEe7qVMZU0Ijg1G9hml9PG2jVFMPduK3c/JA4c7bLV3mZ3ggyvkWkQ0+H37D
+YT+ql2OyG0m9SmoykdHQz1Fs/DuNlBWmBL0OdvWS3CFROdSWy4VJ4asiiyZXEcX
IXhdEgv5EynhSpknPyqpmSn28Ll2zWqucU92tztSCQP4XvZYLYki/2znBIZWCnUZ
P8GOej15NcwcQUXFD3U4izVrbkxNX2HfIK7qgBBl/Lf9RlQr42EhrCEL5pAn3uVG
BK2wACIB5ydQsl3KKRT1I8Nc2wkeFUa9/I94wrFhDOTFIgm1vo78L55OjqSGrHT4
F791JqI23PoYVDBNGs1I0VTAaULlEJe/NWc6Af2hVzocd1Z4/0KlvfXl1pbb9WmK
HwcUyyxsvaUohjZZMqbguMmNmlw+ZCZUfWjFZ/ArPTwMqKYWPTahKWKdl/amlqDg
u16DQPKFqIPmD06OxY/OMZH4jxqtjqk+T03nj+EtH7lTV6wc9+1QsXjHf9VkiTgR
S6iNkxP3F2jC/hC8ed45VFFCVsbjsg/uLqNwkFzG2GC+GY2S1zMdmz9tpk7x9V7l
vg3GBlkKzI1FAcNJumJH0VOTLLOHlGRTcGRCPjm2q8Ht3fCBh4gIqp8X5QZ9xBd0
/n5I1lsc7hjsEJk5up3wm99MXBCdCFjc9NhLPvvIFI0Gipd7QJxU7U93rIYzvmjZ
KdQCsAbqDcri4r0SDJ2Xnm3mqnnoTgZlsjojRxGqd7BVPmZh9As15WLbDx5sxGVo
NodUd9rEzvqP4NGkFwl2QwCyUmvxPb7vMg+mcoskDMBeXiH1BhdmQPSYH4jzjXXx
1ZdDwat5PlMka7WIs9vkQrVFoqXZ+pJEYCGH+UGaKqJAZs+vTVxNHYiarWziL3nA
wd9pwWuLNr77W6cdLyKaf4AzRwoJfxfeIb3VjHK2p+qdszZsriF2DYzGEpAejPkz
OssQWkWTHzJ3Rg4MPZzvLz8ndZq0eNv7OnqUQzAeBMcUcoNygyLmlt7hjTKDCkQp
kRZ9SZAXjHmn/KUqFi+3a6TllYnoTjSpTtNty8kzGML0/CM4fgqmv4XhpmTXn5Z5
X8LstIlPG9i0ylqF1BS6NdvjT+agLK5rsXBeUqbvdc6thsZEcvV2neF6+q41V17u
w88jxvOS4z9Io8B9ywlXb2Wsbhc5xcTNDqT2jgC/u/oRAHuD0O2L92TRgJEznHKd
5Azz8Sgy9PvAA04o7T/x5FoXrTTMVRl5ijMRWy7356ua6YhRcBxQgFkFZhsV2MVr
q3vr2Autj2PEkURPfBu7sXLel5JQu9nqZoGC6+LXqfXbdyJRwOvAI7JY/XtD3m+1
x3zlXve092L3eCTOrcO2SY8ZWUMyeea31NJzmzRxvwFd7xqQyTdK/VkwS3/vyQmp
fRHp7SHKLiYDhnemhuVKJ3y+Eolpq3TmPeeThnpCQdHiCiOUCXDSrrsnC7wY1iwG
K5nC/khr5suigD2eAOtc2T4IDS1S2WGPN6ELoIZasT4eZaoWfbKLELpKdGoK/Wqp
nO/ic1G+LgQQrHVN/FFpZz6YUIzdo3CQL9cqatw3TbCmD3Ex1hd73X4oPCFF8jxp
e/J6fc5Nhijjqn7AlI2/sdOoIrwFyHUrbb88GYmHl5BaAq0t7rTIJnnTE9i+v74O
ijPgZD/ke283n6x+QaQZNwZtGmvrYhDvD1zAKkOGxv4DqJ47az8hJ8mRL+gNDhxH
Z2xjVKuCdmxJaWMzfUSmd+eHSciwVDkKpRe4M6Q0LCtEQjO/i5CkL6JghyTY4eX8
T2tyuwdfFntQQohilVOcfZromRPCYGpNo6qfFOPwXFbCBE1QscWwCKAwuLLioww9
JG8GjxGR/uFzDP1RY/e7qPX73M2orwxWaU7eIBpqqjT6bWHm0n5plbrg4sB/LdNC
sSVbVtWK/KjysVZ6zuXgkYXAHpSq2IGehWWiDYgRWnYgInqN9gHZCbkChfwggnPq
fePHSpj8aHJro9FQ7V5PmudwMlkkUMWBCr0vBCyqNHzPWqB1rC/rioF2HW/ktACo
9lguv2OEnoI96sXYfnCoCY52z5SUnLe7+QS+93ia5VJN/bxnxglevYD5TllMxZ6b
+j5U1YCkRvGa19lxy4c0B9hHp81cSRsL5BwPc2IpquRI/TzCiZgBj36uMF79Bx5R
vfLz2p6eY+mwKly4SgXQBPdC+w4u/W14hWLDuq3r07EhT4lChA9OCCoTbgp5BuAq
bCcWZ2NELE5WN7DxB8gCYfmuNrsfkHmozVloDYcvuowqm2s5DlkpygruPNbYMGJ7
aTdyJ63OkCGVrGw1rbQeu3xnrMNItme6NOt2S8/lJ4gzmhFUn72cRd3uBiEBuqS9
fMKDfpjSmje2/jj1+Qi3H41WPXuawoTTnCNcwe5PZa50NtP3mOt16Ayoe38pb7SP
zkyUiltsvF7ObadJld/7opFiCBcYUWI1fEHpOT4BbK1cInHIT/AWHvild2zJZiJJ
oqOAxykry7kinqb7MZhdIZ7incYMDAyV0GY+vtyN8x5+ohC+rqgJlNcjPpQ9By4I
dbjRH4J39hQbSI0gekfaUIBqlu5bdTYbHLg8DNCpnAxbyFukzneqOMPLiTOIOFVU
VX4pJy9lB1sIiYYdMb/jqTYgXJjAO8Pisnan0xGsWJSbd/lhDEZaH8r3CjSKNouf
/AkgJcl71Q1Yo4es0/7SIkegRI4kYMGOnZy9+LbLpsKdDsc7u+XyO1MT+ag3QtOc
P0jSgrPeRIkBo61jvkEWPrsl46gGxmu6/eCVSHSrbAfaBhjT5HYzPOOJ09Way0g+
GmcNVSkU1NumaWnC8Ale28HGe+Ug4wYUiV1UIRIFD4GhgVrdJ0ZdVBAaxf2kQCsl
9OBgwT6ZDSRT/AdLmHq+lTmvrekyRcdhGMnFHldOozpYfTGwjYUCagxnuwM2fRKK
czEhRYY2vhXGrV/J+1mCIR6PNsBIyBR+XZ0v/G0xuVbHP45clvMewckDC3I1NXQO
qpzr+z8Azua8A/bmejAepK4q3RdQpiiD6KVidtfJrchXc+lDqnglYttmle34it/p
BLqDAPyBrk304erMXxraTXUUp9Djbl+VvXHO2Jt2qftOK/PZ7WpsX83htNrNEEol
r6GByPWNksKmIbeYjVhwOU9kohv+l71S3NGV+AVnKw95Iglosn8B8yFMtfw/RfW/
jWotJtO9Zi19z9Z0TsK3wpXiw8x8A+VD9DlpLAVHmdkckPead3XHxH7kdRiNVid/
RSXQtUZpcDeJsznGZ7ZnglJ9DWMC43fwkkyEV2S1BrKf/ZlIG1PyFKNXE5tX88NY
/W4YejXW1WKSC+vPnya/ZW21vvhNEjZzM5Cn1KBBCLh7YIGZvOLt5Wq4JY1vaZvl
NHewzaqJLl6cgvD1Rr1ubnUZH24lmOj/pvsEcG7jvGbHh4BIyQeUHP72V2SA0ZpV
QBRWVIEIuPOF65rV1tXKoMcinz7Mj/EBh3fwo+28qVDS1Ng0FlyGaovh4oAF18bC
iHMJKH5L4snRJze9/7KCPmDWcxtKztSUqhEBY9IxMBs0ua2h8OvAOU1glqI5XEmB
dJF2jZOELYcw+13eAsiz+B0MOA4uutokHWXEEccuks34lapyvF65vgqW7Inet5pt
idIvK/d0yJGEaeR9MFfwPjQS3OJipmSv9K013pBpS68nkj1MzwuFwR7x7/Onp83Z
T+WukIEm8gsL1n+jGHRAbTy8ASyCO99QqQMohIlJDwTOeXeEBpBtOxVNoaHR1km+
fubUHoPPOS/fNzI7F540WxUhNzVHAaSvdPNvdHS4eZzF08Tu9I2vWTwd3OKZJ0UN
9kiwcALoM60UVPvEChu0AYDI8SO7YvDO0vncDOvMfVbbdnrFFhrWocI/RJ2V6MXM
QU3MdtHbhcoivZvSMpupHkQjYAOMC2ML429dbpOEWG8jAXatuNrYlFrKfhiEn3mm
eHrtRQtcfMAriCPtE9WYfiVGcTXAMiTcX8/B7lakIlTFbMRW2MtbG02Xc5u3d3az
ENvWD+eZS21YOP99AoWkW5jsoXgNeFSwQgS+XahZT8iNk2hlduQGgDH+tgUAhsNc
j9o8J0OCcxQgmbY4UOGRx6/10NdsSFpTSBbY0YmCDYh3gnVt73fIunBPiQzelS+1
OTuGJQKjtheNnndwYKAxwCqQYMQQjNOScervUQUb6d6S+8jbvHD2lEuaZwXItMut
GTGQw9w5uDrqEyWd5+qQpEQcW6Gs7Y4QCNC7e+ocIh2OXELluj+As66gZmnEoRHy
l/UgjgVLbRzRycCFb3zweYO0Qm9Dn4gfvnOUy7FZv9531pkjm05CjkNld7G8Fa4d
eMEVMsQ1jtFNE3J/+IdSN223yTbyqWIzTkT7b+LESt6QsUqmCn2Wdm7AQV9GFKed
WaCxrJVPWMUO1IiJIZQyjYz5uJ4CYscEVaDET+yFUXLmNKdXwMrCh5cdSH5CrnR9
vTypZaw8h8cUp1ZZTCwATlvo7yE5R49K3Q2tcYQC462otlgYzx2seeLEJJtL+36F
F4W8hWp02/Z4MLy3hAEoCrMa6jAr0hNe6Ge1u8YaLlNHoIXSxdv1AJ9/fwopMIl4
u9wlWgEtyo+tXZ5iTGAPM004Q9U2u49Glo0dZmWEbyE1rKyNlNOUbLCVquWj+HEs
eme7D9+r06WtuTVJzgIIxEAU16/u4O8b49O/iMIxCx3PY6GSRXaNbovTz/gYaOo1
9iIoUxc7hqNFUaqrxpw3n7stIA7ccMYjqHocZb6bDhsC4y/N74ByS8R1Fo+SjACj
6kN55iJgaAk/vdC9TNHLItSYlh9QnYaxa+i5VHQaC2+WCht44FUggGBucNddtwiJ
gvOPL9kXQEISINVt9WQIA4y/6jj1DeaLdQ2JHHD42mUV7j51H5FeKDjtwRPz4rN+
eTGmaxWEczBXkHEuwTCTL8gt4zSnAk7x4npWHuzuUbySadQJNxxVNEqdPpD8gdZF
Ef1hO9OShCr7wzRWvPTFWjbQcTSJlCFKaTQz4vp2H8FKAXmwi8qlRBhlkwT5WDjS
5UJVrYkJCJCR15SdFSRu9beeKfEaj5GkRi97xHb1+Hov94vBb6EkqkWc1LUYhlcJ
Brqc2V3/szGL5fr4kjkcqRrt8upZrNdMzzSu5CTG1m6PCVoDX6+JPm7LvWnO9HAy
QyI8rZfMPCYP177dMKIdFxmUiHFndvLyhS076kIowzr4grxFARB8I4ByYo/gA7wB
OeRpEyE1JauVFCPfRyjipSazaf892UhZsCQ9bemRYr+zpS8YDMD1ACR0DcR7DfiC
zBznHNG3UBQYCyhbTsXVKTD1aN9b5VVa5LeMhtIMNlO636TTCwDZnHCuCdd/CIX0
EudD4BmrqF999fqJ3ePaqdSckkx/t/MyiT9yI4hzMoDN6Czx0oVHtUQN2EuZecVx
IUNMku2mljGHr0PE3PVmoLRE39/HC0gDezsAUC1IHTXPlb3hrNymgKVf4Wqxt53w
/wEL0dV07mNX+355lvRP7hxf/xrQ3IXpsGb/1pqueBDmltn/ivzUdG5f+29BKmCX
zhFgPnuq2fe5xGNWrpM08GehiXl1xav+8RI1qH1IFBdsz2qe38pR1B9thM5LWmy4
NPX/WDTNvOS1qhQjHf1pplrVNRObFeDe1AgiQGK1ikffWAVLMTY0mr1Rq5iOcA8G
Azk46kIEchXdlnNrLswBGgkSpyL7hSymZrg581C/RI5qEfd73RSj3Iro85VaRiAG
tH+0tr6dRNDpUlEdlEcwtgvGM6QCajv29NWPggPkET3j7aT0BefN8o6oAfuHdTUY
XGumOy+7zaHuLLOnYCEodQJr+6yBVo/lV6sCCrifrgMkTBVBbHN5bJdDOx6R1iXH
sf648/HyWckNTnehPRMkGNbP6Of0dpoFGo1v0r7i9VQRTOMlIAC8/I3WJammtB/2
gcFRx85unAr8KbIh9WgwRoRsnkCTx9UlXxEHuuNxWH4cFoOVq5zM52fMVeg+CqZx
es572+MLWtTV0OgVobSvq7Krx/ZnTaoJsaB4QdcE+Z6c+j0mWV5HT0Rs5eiBueJn
v0093x2/U3Mj6RXD+uvrmmVLe+vZ8LIZR4/pBjfA51fjFEOUf0THaibxzCeDNpvQ
T7h3P/pRswscSzyt8Gcfs8GlvQTBjzSgHSS8WTOSi4x/M55mJxoagiSEaJmuoF4f
XV3M/qFIfpO3+HGTiwFVrcVL3P37H/ntZNszMraDuXh8I0QYq3vvte8EBgfMIVPU
alpSeTuxt8ZhUmFcOgvbNFfvsjIZQ8s1lWa1k73lTNH4/Awj46TLoSXvbhUEOZ4z
m977VSLpGkzt+80QZOsfyhVfa8exOREJ9RjEO4ZwMK93of0iQmk0F/a/Aq8Q2ToD
kbz7dpZ0N/fFkfEv/FXncpnW9/JBSvOUsZNv3Mv07B/+VFc/xgXi18ERmdtD8+cp
bbi5jjLv3Dv6fVmW8eo5jbanxmIZHJtVTMc+OBbPmvqXL1ckakMZJiS9ky0LKqPV
pWX+D4t177lpcoZnyZFN2kz0LIel/VSGX8xAqjDWjXAFIZVImzwjUZlYIVkM7vaf
tMwTDuz8WxZcMskFyjw8CCunUwpYmyq/MK3rb3cMhUKrx1X5ORT7b5hMmnZDlpL0
lYz2r6pAHIoJylidYaxVW9SyVkKvuDGfzN6TQf5pWnHh56DrO8G5p5oh/YSPMnBX
FNcuR8/clKdi5/9DMwWQDvDXhjhPtZLjC5lByNr79n2ofL5uhfOGmFChk0j150Mv
Pl6XfLO1KDA/tJSdZsA3hwUqI985CCGFvTqgnqq5vFCO78jZUsaiUrPEkbP+Upea
l+l1N5E9Y15srZ2mz6Uy3weOvYHqsmtvmpCaGvD24wuipipUWLDQxW4UCgwLeV0G
39kc6LK68dT97zcqD66kLEQ8Z3Oerk3//XdBctLPidYHqetzQAxEemOkwqvUnYgU
SRqaHcwVpJxTu6Fxf9QGvSkZQaJn5FTUMIIIUzNAAjc8WIw2i2zJaf0pgwtqahbp
BVF/UWg+bbOd13Z1PFwwpJ+6YzmHWFG+prWID2OuPUuEgNMM3XwvZ6Xo9vW2RoIJ
Tg7cf8CyrIzX7bx6FT4yBUogOQoAIh6LiszcEbp1Dyv4PLNUQ249ZSvo/ob5DTws
A0pQXi6fFGswhNpvxFqBjw726/InLcuLI3I0KE3iZ7f5BUEAlbpAEQl8BKH1wRx3
H4zd3gyajPFuQVDjyBUCzh65xvIQpbBBMP2SIcy0B+Mzpheb/94V4VjhW9gDDo9W
Tp7HOSwULim2gB3VWJNkGWNtZFL7wmQNL7KZYz+UNdTPKLlzsge7OfVobTRuHR9x
Pu+H86eXD+dBQGpMg9ozQWuBSfPky5vI0uX0YqZ41vGKEQuJTY+OdVz0efsV7ODm
QEKuFn0wMP4rq4Q6mlzT/cx57w+KsVumrwP+EYytH/n6Db4PClxsaIUW6utUdjmy
852OJuTmbGULfSVab4bWXJlz7Hljn/ypmQAuSGKILtTangPP9UVXrgTFw10zAbAH
RAtlBYS8WwkUUOcTyXNNk9GkkabEzidmw6+K22glQn79tWchb+ggLWYlL3SzesoX
3PIkojCGlaRUpK2FjSOYEhx03101R1Fk4cjHW47BjR7vTPgGm0IOTi5NOTmjLRfj
oaAfolXt+rxoaWs4ikigm/SbyXuSRoEnd5ah90c0VV2SwpjpN/+UyNl5GvfBqs3H
4uH4sUJ+MYJe8S2Tw5Tp/rKdxIpG6KGzsVzAsq/hAYz/+RJ7NXeP3de4nx+Ph4QO
fY5FQI6KcLcxfyjw5a0ZeH2ao7YrR7dXqIBNu3jsA6qvXLd5MjLJlx427c5nJEaK
Qtt+DoOqkrFLyEnR3RhNcSbIeOkrG/x1cWOegJXjc83yObnqUxJAYz4doa5Sg77e
KDjrPl0bBbXYqr9FJnCpGOal5ZyDXdHU+cOipI7XYB/+uU9yqrnlA++RZmVNypvY
DSV/ICkKkJZYu8PbfNa/zH9OBsbeIAPBt4vYSWimjo8mv+u26WW24n+fbsKwZI3s
a4sUpAzkmk6ZonO/EfTZ41WBS3crBaaN7bhAOr8wG5uf0mCFoagVaJ0JJbT53TST
0GaRzz7zLBdbgZjerPq/Eel9WfoWE5poXES63ALGwJtK92Tai9H+ATcyufMZwS25
tENqhcyTcZE8VAFzNGBwj/V1tPoto4KgPWtPoVDfU6otTEzx9dRR8IG39/KtYfyS
bupEBRNG0risj3Q7ap3sqpPWnicvibu+pgmpOQGGa44WLe7mh5FRNyV8NcwI0HX/
SUQPL37EbpjJByqnHSX3M/x3WhHGXxjZl5dJBMcx+TEhlbHhuYGalyjz/uJilXxh
ZRiSDV69rlwGfwEZQHIak5TGOCoXz1k1vhdwT0SXAVf0rwdFxDp+tWX9kuQMYGpB
lEYuv1vwzLQKvnLcFSHZ9BdGqZz5bRX6UP4yqpsB2VhtutBfiEHIKvcYQeZETtxW
i1Sq2jVwi0mxKy/VIJsFOmCB3I9c3E1VjySaJxawtamZf/34QV1n7AgmA3vywIdU
7LroNSdFDgUvQGs+b29oIZ5CF/uxPbqfU4mIIxWY6koFYrbMS0QOgMJWRtIyqEDS
YwhioU9mM9yKEIlk9mPyM2lRvhfI5f18Qx4MAnbfEDhAhqhMOAeDdSxJu//VsJxf
DOd0eS7jGsgooLUacImhZt1nedU40DeXG7haTZE0mVOzi8qbMB+CVlLrHKnSyH+C
aTILhZF8R8VdLBcOcSSy924H8k8AxCN3r18lsDe3NLOJgI5vsKg3Ya4ldypdgCMQ
81k5/d2tkK3b9C9aasGOFzv/YCqQuE2qVE8Kcjrk5DCAKCEi44P/OzuYRQkQQ7gg
egK+D/FstCuXbfHB0A9D0irP+bikKktbhuZW5GgCCTFxRzG1b1R1qgZqhxlHFjja
c3syAevo3zxBE9mxoIfqC7KV17eJpixIdOsko0ivgPWMfh+E9yg6Lmsy/r//4FRh
jVfxdZeHGbYlctHTwlr5mt++PaCgm5dDLWj+ArfKYjU5foyxeRVzmFeU75p64hNJ
dcagdOyD9s44r1MzADs5ub7rhHoa4cAHwu7DqSjKVAXrMiH9tYJBPpEZxBjzm3Kl
if6DPTYvR3MlAJ1bUmgoWN50YuVfkGRkSSrJkKJ/ERzzMlBsv1OVFLR+3CwVtWy9
TGvaD6zfw8OVTOjc6l2j0+v5nMWUxYCM9Lr/Th5DoDbanO1eh24YZe/f7p6gWOZe
1rtPSq7i+qrqDmA9zrc/RMsXqhKfl3KTxoTrqPSHBTEjH6+P52JkVoNhhtVbaZKZ
quCQxh09RaSYO1agMRKwNKLM7Wi6vV0wQVVsQL9/sbMs37j9D9WEcTW0Qab6jrza
0/ZmO7gj9Hn7+Gb4TUQL72nki/22I00uLY0GArfSgXytA91Ygc8TaWvHYOhzvFef
8ZcTDwiKVL1Wfc/LXLtH1y7WzUv3pCi9PcFWXG00HqaNtk5r5G/aRMzCeWlkQoA3
RqOw6Eb6McIe6aRzedgdFcB4BJqfjU1NdKI7xEW5ByUa42GgdZV+ShpefdEzOqUf
BfrC/mLuI++WFOGjrzAm6F+kD73HW2+290X90tRacLvHAt5l7JOwPm0YMMZWrECB
osbdgMK7eW/oyXB4wzPgere9tcw+ZpKrGxgR9cc/JPXJ+CsGNTUZLRlrVcdOYetP
md8TF8BZqR6ZSZoFbfKo4PaPrN9AHEdPGYIfqimNYw9vo5BHeobhSS0zEXBl3bHS
BN2mOISUcDNY+qz8CJl05xxFgJL/Mgx3oF2w34nh6xwi/UYizXe3/LByUjWZLDsU
guLR+tdojFDSno36Tipwfk2iMuUgZGfKayuLzqcp9iErIDQPDQduUAMcN0S0LHE7
h+NQ1XrS3z8fJS8SXDek0FgHDqKvnd3DhwmL8q1VtUZgpWpN5NNQMq3jcmAlOo2h
Vtf0nC4nmWJxK7X4qJtVXqgyLU+FxXhb6oijdyqKg4NAu6KD+9oYJquNIcevClCo
ZJam13K7oGerHRhrs0hYDUv4bPZyPk0FgqhHaM9oEfolB2L1iFyHdVxp7A+J9rcS
X76OcBXlnjCGMhIN1SezwnUa0u2fElhLMN51g1TinFyOr4RT0OEN1H22K/txV2Yn
Uij6hAMxHD9DUMteqq3n7ncAPUCcAE96ISm9Dn157WaT4UV54Y0Mqfqy/iKbOsUS
dxz5zuWf86gKsWFb4uv6oMXdPMMNK2g+5uNzDJKD3HBSLE1LjH+VGZPO6DNfXg1w
32uzIrvnPE3tPOZat5GNt4RtYkZCQmXiJSDn+ljxcvtcTTyy9w+Eh3hLL3QyOxlc
V0YxohLB+oaailDWalSJXYLM2d6O6UylUPGYaGFd3L6C9Pgmv0eD/CA5nJwxL/1h
NKEybUIhOqGlog9YGqxl54p7/gYpZpWHx4kkbT8+JLZjQdFq4DVOFKy0Nsff03BJ
wPWCrG4U6BJhPMdflPMgOj+psqdqb0iplUtV3FLmf7SthpZ6SYul230lHiRYiKpf
LXL6h8UUOYmckIM/KcfMUEPlWR3S3xQPhyiYmXRTXYuLkHo/xC987m+sXFQ4E+vm
J3hSFoP9iW+vizXHx9SIfJiYhnJzbiVxLOtwpq7DO5REmlXNQQ4sDb++dqi1z+be
Ms/s3Y93ssIr5utjfNWTrPiIUezvGTpV4AXefjjJqrzGIU2j2iVP0dOTkhLwVMXT
UQoPsEQIOqF+kQyAumm0b013u3o7h+2iBg7gjmy52Rxz7z9a7mpmwTFHEtDDEeJN
9/kVO+8cpRpayxjDFIn18vK3BqF7sp6gZJN/2RS5tAxNPKJmOBQhjcxSeFqoqX7a
FWilvaR6FXGxHleq4GQWsewdSL5RoGQ0aekXgxBNDYVfvnBRDQCy0IbBfQnS7BzN
+jPV9ozOPPQied6GThsvoSzEsFote21fYK6uvaEAI3zhqIrzn1BkRg0fq+gueUfM
+1SAJDWVvGwi65sd9feoFxxXRUmkFtqGGRZEbyYqGnpJ6DWQ/KTP07wuyn3Fques
6coirfj7jLCdFkO/fEOvimxDoLc6f6Wfq09ZQlOM+JrxzGu4CECepQmv8QGFBJPp
Ar4wYtWeJdPTppYqRE6krevCI42dUAHMRlJbRTFi+PF/LCPjrdPDNVA7Bbfy06fa
ZjAbM3VZ2WIIbmW2G4JnGnVgBB3g/2NYXE1n5wUt3Dk32e1awXsou34VOvzlPP2B
EGo6K5lGZa1xl+6GKA0SluszY8/jBfunVIga5eu+u06Q5JpGXG5WSnBNO6eDZ/Ye
Rr0VqKBGOPPlw4XI44tMUJCDCkywjcxdv4XMiyg5He128TF6GZvLMwb1lAjgLho3
PQTWZnGa6wMfmkdl7qPG6IYcpoKkTvoqzh4g62lCHiHmrfH88F26ouq4rexWe7nb
exgsC3o8NwbYo/7NZj9ovnjQ95oWf+Dc7wKS8ipPUsJBwLJ7TrXfWYevwQgFxQnt
ppIozU7IfxzWPOIh7U/ugl7uhmNiUHzeyDNWMeFaIo4k4+2/yv8hHmL1vrRrxEdp
pz07w+qh2xWr1YAtHtonM/V3fQFvB9ymLx7woLfVIPV+kxAdgsVUkAtc7w3sC0Lp
d+lWDIQYRSWS94TR3vdKdbQdULEmjbXpnsjnhBQRygJsW0LfB6kqBF9QMnPD9WOY
EgVSd0If/m0Fq7yP2ru2jc5hdsdd8J6ZgOo3219FGL/70AJkA2llMOjchJ+yJzlG
WcuVCoaoWI/baHByK7YKvElMjt3RX9nS6fkElbnn/b0KuAuICaHP5aMx7kp9STjt
j2HtAmMoLEUlCpKZwFncR0NVNDHOABQRc+Kioq6mYW2IVaAHtz9aS5/5IHMx2vB4
QYkKsw5T2IpsvFZbl55S+IrlYdKRehuwIHo+YzbQ0BRVc+BLPHkz6L1MKEeolv5C
xURWwpB7NqgGN1GmdKBwmpUtNIga4R8mtczjZVPHjRztxivu9yM6gzG/htaSbXGp
vWt7RKCm9RIhEH1s79M+PwtRXF0pFVCiVyFZ9jni2/Wh6s2rNTRiCW8RyLSo2j5S
L4vNNiwg5pFv92rkiL2BlG/EW5b8OKDJpSLClpZwFM5Wl5DT+bXwIWZlbmQQ6SKm
jnt1r0VxuEo7qROizY0EYZ03coLsQgeEoQKk+Ww+pPuAkOdG6WFgMYc2SJ8F4apG
VD2+k8iVmd4XO4qNukxGrUqyhYHLh4FuVKlcUEQWYcrP3t1YlbsdvmKdFCQl/iJg
aPapDMa6rTZ6k25xfpFojPWbVWGwXxGL1D/B+sRVFgWvGhEFnGMEuOkW9ibHMrGq
csOYWgAo3JYO6YNTBNBXDk5l51Unw5ckDAjvtvZHhO3xPsHUajf8B8qXLdK9MVOC
VpI6Sa82p9DAf3gRQUc52FOKBf5A2u/8aUX4sNhEbd04MKGEEeoAli+RNq/IEAIs
14QAvCXQuKywjMifVnSF5lV890K0kGi65F89A03TZogu1Z3DwP4QJdvQHHyNXMcw
817W+49kkxWldCMMDCs0LE+M738PZV4rleEMY2ODIUHVNvsKVhSKmqshBBtMYhg1
4Sfvp9V3GoKSS93k+uXXVPIhjn/5STqMdV9NXhBxgplkuVRClvRr2np2qXhvfifC
6F9JlKNrzJ38HVUeyMNXhoQPZcsRBEptqBDtuNwzrj+svkfUvujya2X7aJ5LAsyp
QyjvxzqfF07ZbN1DSi7Je3oMAcBXjPtn/YmBvgA337QYGg8I5Sbw1UNopFy9dKVL
lFaITlIiEahEGFg3I3pviRVW3hGI84oj2cro3iGLcVeRC9C8DdIq8tGu75kU1eCE
vviX4VqRuU6QXUp8v0QmPqU2oOw1WQLIG83IcGNVGikBhQalZ9pTNJew4UHh18/2
zbEqfps3s1wVa7WqaISX87AroW+BG88N9HK8gvlNBM7o5B0t5UJyp8jtFrKqvFUo
vpyVyM0gO2B/XxbXFy4JDlXpDOrBnP9quIUSIe5HcaJ7u7aRoEezVzJEES6Qdsci
tTh1RhgBCzlineslDqe67/ZL8NLy+uhjtmuJxtr/52Lnk54fBv5ZB6ijSoyZB/QT
9iwFUEEXsGjF2/1ri0iFsv/NfaN2xjS9Ruxy30iLfTBYaOV3h4kM1n28lK1FCtls
yESytjwfQzYlC2iYkhTvxW3g7v7hywDRQPeAic9j3ya4vYe/eAnlJ+Ja+QkRP9Q5
9R9alQ7vMx7yZCpw9LrOgmI2LzsYN5r1iTip4zy8QmPn7DRNkLcyXJ9fEXIyBX55
MTJbA/NF2EXcJZ9VXqqSnbXrHhsfHDprx0wexgVrR8zS1FTX9r1kMCvyqQycTZEp
43m+VR8l0sAKJyU4TNOvt0UywReMDekbn/2OXPStEG4VslvTk8By2ttnbtCxku7R
Dy/Qv06HV0fuysUImik2VJy9JP4FN8YcHhzq24/UGLCmY9B3ZXwv7uSnEoSisXHw
DJcIpRQBd8CvfIn7mljRdieQtlocS/UDRvFtHZVUTCA33+0v7YZlBPrrAKv+uRcu
W4uJ9ahF0DosujqeLWhzGqeMJ9RmizlUqWbZYOPUxk3ret5ICWhtimAXfwBfHtrs
EzHwb6n52zQFesn8bEGYJu8o6Fuxnl4cVWnzcqcbNAdZlfWeWE2lTlzqcYHda1tO
7UeX1UiVm7E+2HIuXSiF5zdP7EBKGIMDRbmPv6Fju6y9xp73iKMKQO6j6MPlhWKy
s+y2mmw5YFgeEhyQmSYqZ3G851Qz2Z5xsk+gGkC7Qp98/qkgkfddZ9v81Zq+PV3d
tEq2DLDZaC4JOPthLwinzLf5IntbQVg+s6B0yYMiu/w9t5Ht9PY3eRyVYw0AazBw
s7XPA75acGFKeBI5iJwv1dBM1HdteWL8tuSb3e5W0znVKwms5XU2INx6N68+AwTV
zd2gEAG5TNn83pBfCDj6xWPs4qq9qtbTVQvpEmBzjZvd+lfr0rWvGf6iLZNDbrv4
ehm2Fw6yVPODFaBUyeiW6qcZAP6w1/xjaru6NsKU8fws1XewGORruN0l8AJFLbB+
O2krSQFHxozpLeY7eRSjyT5XTMWbsfrMtWlZYI0SrDJchqGnKyu7OLXLuJbpGlO1
f0H/sXzDR7jeMioNEj1JYqM52MuYm/mQ/EG6I0FGDCpUocjPVtXzLmSoMOCBzMO/
VYUDPIdL3MPoET7ORRzieqqSKGe0rDDv0mHsZ+yDC6gMK2zJBvoB9empBHoFMx+F
toyDk22aOSJOk7CO2fHI9PEUd7hUJ7vZlT7U4xA9Ugsyhmr6Q3QhWfWFRdEefnZZ
RfPrlcq8Xsoub6/ubdLbQcr/hLBG+x6DILHxLv39fDfbaQWFl+BJ36YieKtuizwo
Zv+4nATpuZ56arUNEWs3QOclenYsXMvdt5Idrz6na35EevSxu/KkKXrYWGIy8zmh
qyDyWKIpq/88Vgw6bH1g2Bm8XlocwvG8Kdd4b0/J2eex79O44EMp0zG5unYTODw6
EgvMQkjf6tDgj8yz6MzG+oT5B0GOfBv5S206fFoG6LeCvf4V0cFpMcO4f57Xt6Vx
LhnlBR5lTAmBEU3E5Hu6LOvwidpsuAQxq/YmWa+hzlwN/24Wb3YtJ2oYydK9pG11
vRyvyGr63XeysSt+PRFqYbzUOOT0BWYB/2a9iARRVHPtL2/oFdEM2jjuMh+UKqBK
noehfoyyRf+k72yTd+gljlJ/HsKUTdyucC+dbXukps2zN3Uqbkawe6zeDw+fu2TP
yNZbeocU08h4rymRPXJjlv1SxfgTU/hTmEm/zrkYXLym3kmS/nW1fkfsz+qH/DG9
wuDT8MA+gbSNwhBqeaw2Ic0O+WFkvps2/MyefIpgjWMS4DbhEMouo697Urr+lHAf
jvUdMDKIX5Dm7flhBOUrtXVfaielROedSh0edpIrAe2pCJYl5OKhksG2AorKdWdZ
utbJTBVcKuxgQnNhxyVswPzAXZHO5RibLQhKlJUx7IQcWNT77Otxiur5LjiNSpyQ
UDntAHYQL0SDTsqFMld2XObH0AwgpULrrdMqiRQk1l4MAK9abqL4jYlNV44fW+Zt
HABIueoZeGWgfvv8+nKKYfzzI7HOes6L8azBYlelZ2qA6h/tM7OJ7IYYTbugVhlu
PJ2hWB54XrTZDnFPb/TVZ7aOetjjKom5i4f2xqqH9jPAOf26YyWyJDcI92phOvZi
xmgwNKGTpasX4dNL2RBXouPMv+j1A5Cqm/cvtOylu2ao9CmFRSlEL51hYFTdx6aa
eIBgA1XaEQnK4kZPuB1/uH8+mCmrJy65cmYcsDHDkK8y1yEdnHrTtAEMVapofOrA
MDKGxbo/NFvcC/AMvb+vmzA7Ml2UAWER+BjXUHVrnKoJMgaNM0xrVOcLeSMHq/sF
+/6Ro79bFI66ECi8BUhcAT7AmDWBRYQJVFXcd4uEJ3iVgRfQ7LzHzqeQfdfz+clY
NjMWPVLJw2JIQCUtpgP08rReYulVXSvDQ7RDrOXdBwx12VmcimWDNgFNweyH0oSE
EOEHTjjLPHWgKW21Hd5lkQGUwb4rPVlu+A8Cuhf/7vrWyjwSKksYmKTMR2LXPqIO
fLe/U5vvj+nesxVWqKAOzViqFDCKXo0S7F86V4TyFEKnDDQNp7Ysbu1peB4/Z2yh
fTEUdWV84g4W+RWxQEEVKwCbrd+crlFi/AWWV6QmgRjJ6+FWSno+xpkPhG8Ri0Od
3wJU3uutfC23QBleVgEjuxdzJI7XIMoX/Cv21EB18fHzhNqYKh5dN+c7zu25ixIw
22bXV8tNmQE7FQEEkIsbB5/m/HEBqi8muJV7tb1F3tCS8EcymHl9mVboScIzgiBz
gEglLTdZv8Xo/PEQW4OguFHkznwTvYwRtiIEmK4Z4BQhi1zZovXqD9yXQZF1T7jb
5OgMCfTu2GYL4J2aLguKjzqLWlmWyfOsrsRd/0vdhpcksaNXP/JDKE+37PcxnOjJ
DAflh4vy7KRAQFLIPFYCXb94c8l0+8A4N3kFgJyXaUO3GZD78O/pfyYR863xcfrh
RdYZY9g94PxbQMydh7Hoe9JqV8jKu4Z4wacTOAPK+KYkeQTqFizczT4ipjDT3luX
SFdk7Y2E6nWj5isAcHbU3cIAfC7UsC+OB+VSK/YCnLoO1HANM6eFzZyVEYebUZqM
mfKZ/Rtc19tWB+SsSu4VUFIu0G6jamoXjOcDh5gPO8qbhLIQlf6Uj3YEBQpWgDKv
+BHTDDehC7FxjADGcztfc/NdW2gzZR1W30tmz8dpn1p09605hVB+Qo5XQ3eol7+t
HaMru0yuc1hLvmo2TWEHiyOG4MKR4mqFNB6Cb6XYAbXI6hb8g6ak0JeCSAu9Xt7R
4fKS5qYHBbm8GlcK4gPIXtAgEBSfaiCwX90AJZNK0XCU56qc8sXoT0iCE9ShtA5G
uTYZEjf7shvH3EjmWX/omAr/DCrLWkkiUAHalP8vABnHwGsQAi3N/CdOmCSjF6EY
MGbLPps35MffEkKBjZlgf855++A2+nb4Alo3ZjQokdq7Y+msLxAKMmEQvDX7d9mB
o2mmK0/icqgOwJxBh0Gdbj8P7/975ZO3txOHjew3qlD276ZEN9pRekkkXoePZ95X
XcJgElpitzEjvDPP1etndLsxVavxMVppWsGvF1XAqln0joRWdlczikx6BlURngrw
8lX7sR7IZbvFn2Io2Se9o2P1NmZo7YiSK/SdswBj2tKnyka8PSRIwnRJ0sh/1LIa
QbKB8ih1cD3vgVNE4/IPqWbaXwc1aLTI3WcP+rfLwtqJtKxPS17EbV7mFLzt6cS7
3ejdjL3LvboBtboVGe3FQnWpKltNDKB+/y308anqIl4IXHBMxmKzEj2Ht1gVyrlz
24lG6flMjqhdH0Qnca33a60JMYv7UdciUYVBV7LchrY0RHOjbJX2tXT4PqD/xAt1
h1ri3U8tM95XQG6MsIHBD6URFhkwIJFSIDifgpXXC/oUoeyGFOoi3eODAHdexCDd
smYdP5qQWaSOPelQhERIO7mtRrsplMBxMWHoGZEP6jBTazULrLTUsiFQVjVTO+LU
2izIvLTUwT8Qxv5NyzXPB7G4AuCZejP7RdqFtdVlVK9+PvXxqc/cHUi1Rm+EXJr/
BySOAV5oM06Qxjcma3nw3zkGNtnzn+hiAr63IRocg0xnrlCDVTBGBWzHFiAlxguw
0P6AxrX4rpj+KlqTnVD8WY3YjWE2Of1om+wrMbMyr2WBvN9jElqsk7/dfOS/Z86P
IQ3pvpbT4drrPtG7PntPVIvuRBXa7+bFxLnRfjlA/ddIPJcy/vM8g0S77ePcVqFc
B3gDNco+kuvZP8nQMu2yufwBEg+YxWpO6bEktLcKynHUBh2GvmdMMWrMxySo+x2o
j4OdXLFSN7TGuN6cjyMMRx4GfM0mjTia5Y9aXtAzx/aX6lmIHXfEqgDquhBGUvoR
/Mw8vaGtMvvhErxHE0SGB7R5Vl1AGUA8BCjmSKvHUntkC4gi6dpn9uybOtEynpWI
+8veqxpSJELaPSzSV3icNi5rVdvJGDp6n0Qj6nzP/mFW22J/bIRUnFeMfKfj1xmn
CVU1Jrp2GByyFkUQ5UPLXItipwPDA+qpp2Nks3cERQNKKUBYIg3Njfp5jRLkPHb6
n0rAXoYyxVLZzqD9pPcPKqGfCts/SZoO1g1PM7bTxPNY0O/sP0cRwEwAjHkrdIFk
dPFzmSuNksIIDzU98gugYCxwidZSMnJ9K5roKXTHJ9ga5WlpHrF/sWbYLdw2KGIv
e5G2uckPbvfrXN3NxbPBCp/9hO9k6VbJvgmyj6LdwupaAr+b2snd7VKdq/aZIk+8
fPRhD+MWx5nDpLjCke1u2vVCPK+6tX9TRP+qVKJ/+kaUADWw1tIj1oj3zBSZux6T
Bly3P+Rq1pKRV2f3a0f7jsy8Z5+F8gJOk/IYQ03kCkHMpin6EBqrN2/mnDqmxaSn
nXLRa6UhqUujzv9PIn9exbxtTv/bu13Qs+Vggg78FqPPrkSEMz6/jVP7XS4tfrFk
wIK4IoTyYv7sqoDxCtsQ3TTJdR4XATkaVnGKPPboI+zgZDgMzgilwYcJulMpk+sA
rqgONW8o6IbOo4KkIS+Ag6HC5SKpCuFAPqKZASboYNGXhBuDPmcBpPg4lKoknRwO
Gv021TXa2OuYD067nCMPZOUHZapWvG36PWYIrUjOWm5SUJHlnkL5zdkKgiyY/Mjq
4FUsESFRb0bS32EH7jVITrVFrjH0EZ8NGZMWEI0HuX5+EwEnerGrDZ+9saKUPCKL
q7OExXZQRLwvUskoSXeBP5cS+SFBEnQmgVjCWPYTZ1oZiPxgFp5l7AeZeT2FamAZ
Ji1/awZ9cNmUjgfwNlJV2BOE88vl3VQOFOy43r//CANRKyZbpDSvS55JBbIj7mjI
fnQb3B15WFW2lT92IuObdDE2fOOFNeZcu+slOWZ9czCLu/02lxbbxLn9ff3N1T+h
yFJoBQLYWFx4GpFSI5QQBeptq3zFTR/9BTGGq4+G8pXVe4/npVkQOchzFqqXDsHy
a4hgP4FQZ4E8wZF2gO+VE2bpF+BPovwbWB0ICgV9VXR707w+M2FbSAGRA/PFuriX
sCua38Lt2N9RTbB9IWj1AA1YD8K7dhyOX1JQhqh+XDBDc81Hd9CQ4qa5jkLCYbz8
uTxWZnFscYARoh2W1fur/OsKuCgK8VcQ8ZPJlKqApyKMRG2ZN0Y1CG1PufGTkQO/
EAuEy9mtYdbxSwjNmZAYfEjjctMdFoqs/7DKE5AUiTj8SHCqSInNqTE/gt+fnyBs
HNFkKMGrPNFSLT0+w9z5Fc9ASGQss889A48Cf41RUvXfJXWnIm7Jt1eekVvfaXqU
PssVgezNwOyTvr2XJ55iDSRiZnG9jLYxYf7kyvMK6N13BqfeApvIG6lv2uI5Dz4/
HN9J0EL1I9kX2nV3vZdZAjnjh+YFkDXCCqBIDp/hn+h9qAu92NOLAzhTqYwC/iof
R4BNuQaFY6GcFS6VRFpB28cVuNHvdTu3XJ2SwK2lUNzPKVSXtCZTBQWytmAlvoBM
DofloiQKZ1BjIVd/9QVAbRoDYvXqt4UUOcHJiy6bQ9aqP+jIcPhGBQvZAQnmMKAK
vrkOU/CaoGi4+uZHZL1x0ZJpHpLvpYbnf+u/n0gKm9zPLvLzrtn+xdPZm69CuFzb
lii2klxWgHmsRq+KZkQnCRUzG2DoijvthYpH1GjHqrG1b1SBGRZO4UxwroyTjXDO
sd3O4eqfQo0KgtbxGSYslts3wWpZl8+U2MjyhDUuAOJd+EV/QD8Z3mq9J7uccogq
lMn26Xy/vHh3/wcMDHMoFEp812qrCyfSJrmB5MSjmI9Rl35u1x50ZLuLxUtfmjqw
SISKdWiAbyWmWj/lMUac+qlA/55XwKRwsXC7QvoGMGn/n9aarU1UmisQDEbm+GQb
+uwIif7A9xKhYe3+0gzxltbc5Sb3E2MjlruQ0FmkvwGqsPPDRWtPeGizJJcGurAe
4+AB7SK8fxr0KFDsaYRkpHbu6n3MplOo3U/uN+jU7yebEj5Z9MrsaB/ODpnr7Ucg
8CyZtHFg2o/BWCM4qlr7lPJVYKVK9UT9i2jfJYzyqBXvf4FNaWgneRs8cqdhE75a
9VJOL3BU6LwBHbvcZ2F5XDzeCh4II1sVtXqh05Lmp+DiggW0huryqVl5oXdHRufI
cMzkV1gF5fW7gA4/7oPfMiBgg4VxLl3MsXCwiejAKfRw72nh4qTyt1w++9KdIQEC
e7vsfUNAckj0Sk6JNtfxMSq7bbvqrUySAwgVbIjXlJ67y4m9aino8HtRDAKM4K5N
YKCxoYvvvKA6DRi4UPvn6H68g0jxIAnch5vHfboGX6qaRzCzsRdiEJ5ioIOWnVjP
vDc+yhKc6pclJYvOmr0XGT07F2SKWrjz/qQGdkA+zX+b0E9l4dgrSnLi1q6QRV8U
ih2vIpgHyuYa04WC7Rs32vfjTQlYZmNSqTSTK3Gm6UgoEHZV3vBHBPi3OvZw9UYZ
fzcbuMTQms9gwQ2kJWMurYklHpTfgwzzzEHhKqid+DiUBPW26c8mQG4y25so/uHv
/iri4qvVpZ6OodWWq4IEmkBSGJiO7TkrQFzUb8YYwEcYwvY7xBU9CH8kO2npmlB5
07o4Ydz8xFQyjHF1Qechq3A6ayl1egcjA31nfFHHWA3jS0g6gs1iHEhTM48hOC+7
3r4lMoDTG7aFqZ3h+1N8ZJCuqteD7uE4Xu5qvwTfaojAdgX6PfagZXTv/DhHScaz
kCTwdigsFXhvqruYaxnGM7HUulsnpahfa6SG7U4qzWaKvD5zEoIYEPz4MUTuFb/5
MkkZKQmkd2BN5aj845N6Lbi0dihtZnGW5R7lLEqqQ5/w3zn8ce7I82tXx9FW9e8T
XN0Z0JP5W+ZSlgvLGQfCt7ePc6ZGb0UzgcI5Wpow/qw8MbfgNy+GdLUC1W0hOTpc
Y8TihTFHda8iwbCKaH5B9tW2WgOPZ5u+ACAS9mvr8Hf+j49BMdNe+nw4k6OOVDBE
jVBmRh0LiOSVP6fIMNhIF01UGIe027j/SNy+3dLYKTNgNZ9lq/WzrKnOzGzQ59ZB
Dg4x4Xx/3CYe6c/doxQZUcjLn/fNTAOY737Lw+dzMPKuweuweCDLtfOWDptKkkBs
+9nIREuBy0czxZLOMr8RBG6OO6k3y3ZU5Hrm2Kny8aNFIPNoCdZzW+MvR5xPHpPf
H9hQUCixpW0pZp6FtNJmIv5dy+0QXskWHInGMasFEWK5NTVrqPcKM0PPSTrbKoXd
ToUkY/bxM0HxEOr3N6fALKBra37Jyvi010aAdh/i/pHbxbOiQnEo97ezuYN+uQQs
SlR/SD7q/FfJIRfQlo1OaWsqyJxAh1rR9ht2xFRzrFCq3tTWZS7ll9wzPQuG/QKX
G6ergl1EUrte5cjvr7Eoaj5bVffIS/y1WGBTep49bYCgvicywpzmLPzSSOeXD7LU
5CBxmaYzBjA56vLZZgB3ZWWI/oSJbCv6k4QkiOS2Y6Y49tZaX8fwCo6P2HZ0fqnE
fGlyIemsjD/mvK5mViBYAAyV7/NyvOMv25FXmj70GWVDPZ+ywE7Jlp4VqaS9Cpv0
2nxY7Ws5XG5GRKAOUKD12odxQxqzvx8mjVFIw70M+uHHVDIK91DRnsOGgX+9jsYk
3g5352eQrWQFgRy4Wv2Kf/p2u/KaqQ0+fM/I1r8ctB1cfYQd8X5HkjG1OfW05khK
7mQpVdneYWPFSaXmpLihM93rpjxSkzl0EswnT3/6UGZ5bTCUjSYHaUuE7fk4EhVi
0UmSWQGu5bNM4rwQKthW3tfckjIIW5VM5F3ngODG0o0xw3qtvYKJUp41HTh0bP5L
KAPdn/6CrIo86yY8CZDI57jrpxVDg7Lb6KuNGH95C4wQYdl8cD5V16crQzHEwAL8
YXKZrhBtu9dD6V8b4R0mr9gWlziuzSJNeBVv1bocaR5o42GrW+sjO3GtmoH8pwLb
+DPuZ8zeo1Jcuu6RkPe7PK+xp3m+8y6zBDt5sy4d/kxW22X6Gk221yJw4ILBchOj
SiTFS/m6gHtDnS2SSSbG3mYc+/qfxYAsFwO9Uri+DcWSj5f7FnpXf3KUAbwUZiGy
s9xCB88UUBbxupx73DGHpenT8qHMTkhs6TMxXQmAP2e1458Vkw1vfLPpOOAqY/Mh
KZ8hyvTyuXWinM5X4AYA2YGMD5Wl8bjpd80epnXjDqqtnkRQYgBj0zXz+SiQdICq
3k4dkK4ThS4cps2oZvB+K0uBs1HG+0XDaAsnc9JBWirXj/cQa0jexmX3nqROINLA
k+vgOivw4nwnT4lJo1SCunW0XscnFOxIYwCDKQ+821CjxnPDthdaqgcfu5w3sPde
mfKwlFpMveo8MvNbJKdf6DCzDfUh6EYPXBdGBO+kRjGilwGUgDkWODzm62ilHIfg
iPRIBO297TeIVXp0FAXP1uCng2c8f/mtQwsCtPurvNBJrbq3uiXiika2efgNlTJI
KlKVS1eCNVxt3hw1W5OhM/tpADTalkmPvLfd5sA4U2Noqf7JTZoqLxWegZ2Jyu0G
gY1lnHs6lQU3leJ3FpMePDr1F2XYpxFXev31sf3a/Nr2HEP/zEr2sTnY6h0NPAzJ
ci8PKvU3XZn4lF/i0VKT0sEmylZ3gWv3wvQ0N9RePD6z9lRKM6la3LWBzVXSLz48
S1egWFTWaTvw8P4+om8h/bbIMj7gUrOkSfmTjvX5AZ4LkUt5AABtQqYvhZ/WjZ7x
pkFDTYdHECUVt9Z8rc6/V4KPAL5xw20o7fRBdNvY+O4uXvZNyAIS6M8pa+UsuiN7
GMMfGkz2fJEemBMlriDvHcBXS1zv+oMBcxyFTKh2B+fmzEd0tXZrYtww0YEsWq6N
W/BqlHU9aajqY1RSpcqsYZc5Rz/zlmgYOqjOMJOiTz6oHyoOo5+Qmq7h6iNlEghe
UJQ+DqFbmL2JfmOMFQXzq20M0fB546sLWiXijEFafDaQajEv9bZe4s+gHWOCpWfI
vEliXIUsGocRhdmf4wYcIxzSzlujihLdA+Woslx/hQQYxm6l+XUuG0kFHPHvs5nu
zNLzop+ur3C3jzBY2tbCESrjaQ27Q8p3H7DEfL8ku99/oWRiHqA3tHxvH057/vpQ
I1efxLebz365TIQJCZQcR4i6nSTAGr/yR/6+voWuk/T5PWvqVQfe/Iz2jSiJHww2
0Upf/KxKP28iUcQvogcRACgVk8ajlMWE9r917Lb5UVqWjjhXE7J9JDoHbMNAlZrt
65budtL2farsrqPMZSI5w2slYYYpU2pQRfy0fSY+kx9AbTa52/Qn04AL2ycOhOQn
qMvQ/BMfRKvhhB/qqH2fv34ELUYF3ZCY81eS4WBsjUSZ7KRldigIWZE5tNP/euDH
lvSK3Uqgayo6oiaHpDixlDGDVEmuBBaNHCZ7d/rbKyBV4gLcjBtTbhjYWVcffGX+
sIlzl5Nu7vhR3MKjWU74lX+xol+44jCQGGg8wLjPyIvdQ0T03MDjcFTfZusb+oZP
CcrxhxI4A7qBeaI1W2OBe7zWcHc+GLKjZjbi0TPWEWJrlX5LvbB3lXEL5ILrEd1j
hTKzLqPgHyP+cN/thHZKfEzf3FKA/neJGWQoOY2VtD+bThkTtA8m2wXRl6fA6eED
tmOtOrBLeXx8g1q/GHaj9Wbtp3+M9wN5mQ4hVI1SvBItryv8/EMuWoPH0jbtpsC2
2+272ptjadhC6W61Sj8XK+/JNWOQHH9x6bYlo030uJ50YVL5qDzRxQekLk6vGTIc
BZzNQy9zq5tThtfufcvRvg7AtrgpmUH2/ytJ5ZxsMiGFxlqUpJqkzaovTWAGmy1A
fiSCh4pg4vAaaOLcATwPfAx2GGpS79oz6RP2cFlgvdZTH1bnlBQdDKqeItVj9w/Q
NygIxutNPi2tE4M/PVv/M2Xja3CdKfH17Fcp3/ewhUoEUIrQeih7f5sFuPbnxQzb
IJfxvez+4tiro7K8+a1O17I+nKnPYCKqDGJzkSzQBqkLRO/gNwcjX0sg//vtz3S0
0eoWRCUclYWLNshFEfM+hLA0zGh9aIRlDew3C/egzKzbZVeOW/kjNQx7xGOl9+kx
eL2O2Z42cx/ygbGD+ynqsjHYULpQX6x3+HLKOUj7w+yyltE4n4PChDnZ32ivJmK7
aMOKUXjnjmh5ugDv9U8nOnloEe6eATFRCWo8US3aLB18VkTta07bTJHCdSDNNGPq
ST3019rxZ+SwnCG4x5Cvj9ejyC9CaN3HuRFb8Ox9x7OrQhmVTrsxf67nX43Ukfb+
aM+P6P1bfh/iYgAHhJr4Qxt5f+ghP7UhAhd66XulHE1sqL3ukakO507tmqiXKJ6G
c/8cWndTODVTolrrV73QHsha4xTeZv8kRFMdNIB0eC1gPe8Q65Z5xx+eLmg7koJA
bjWMnkpgKSCEL4y/TVRJdhJT2bt9U5s615lfOqrHpn3dhXktHWpnuoIeqYmTIhqm
0hOP0JBk7ZnrPO3WJOL4Te+krLc+diiMrf81kHzR/bkJ8bWUQ2fz2eN8F8czQhIs
R2WBvf2vohoOJh4IMrEOrE0cUqlvVh7dYk/cgS1c6guAOYCi3Iru7eJB50fW9puu
pok/GWb+a/fMBUpXUX7peqrB05A+tB3Gd81zboKl1WvRY3k+s2TZFyTJTQ0LdY8z
0WUZxJNEf/GCbnB4rnTOr2D75RRcc6GhGkJMPk0Tt2FgqYGD6qBvrPqvRUzDhnRJ
S//virZJeg3nSI+HY2hN3Sg8Ai63LcbxaH2UajppfcLJbx6VCHCiK3bgWshV+/qD
QNNWtWfdUej428h/yAHN0ydDj+n+F6DpaTU+4eM5AYnzVMEqkFBpztj7bwYUUCPS
HYUiyAkYck/yO1J1OK4LVONQXPNgRhK8+EJ2oOLvHueIZ2e6/cgq+9m/ymU7RPSY
o8WV60UOtpXq9o2Q1MAhC9DWDnu//uwLshyqW4c2ipph07wnCw0/lsSuEOiuRwCU
Iu6/lbfJGiZS7OF81WsX7OYb8xGLBb17iQ06eTZ/1mFFhZPL0rx2bLZr35dN9HmI
CWlFT/dSY2y86WodlZunIbrdsS2EODXLyx8+4bmUHKHLUiTiTQ1uhnG9VQAV27Im
s9eF4oDEHq9FTjXMslS1T41ecsANApreD/qA6u3MLMqeMT5Q8WBUaCQhM9C+4aAY
dwRN3XeQr1Zcww2Zt4qADwyxzXt0pCyRx6jOIuATz0GPnre1XgehRHuz76oFe7mY
aPHdkVcnuqTPtbqjapH1O+bYIrCKAuP0g0ApR+F3khqKY7dQEu9ZylvUOzqLmYRg
yerKMifx5UZ1R+w5wi00GiVOZIAR3j+edZu0RKybUEBvw5yRcMZ7S6sFzZ/CrfTI
YjBfqw02bwUlCBkByskeHjVgQngUeSbO69Tc57x7cypF+I5R35MLhrHnra7teiAn
G1IsdEMd2HwBnKJpxyy2Kg7lNx4A6Y1PmR7F5FlePB3QxCIyerLMizzidrMkKIg0
7us+TtVfwK5r4URiRdGc8+NwKe4Kp1CaHxkYllC4Rk9xRWQeEGbweKHeLAr6Irbk
cjsnTEzuKBl4fCe5hUpyblij0luWjHdCtHUa/egEtw+hRdk2fsMT+mrX98ICbYhK
8cpIvw+husudCLQqaEUW9Uv56FxM1Mg/aC5B9NCuzBAzKKyU0P+6f/FeiwBQx5Sv
Uz+i8aDDfiK8IHRzrJj465CU9/XcKwiQ1TYRqPnO661rxydj6joQ4OiU6RzrJ9r5
OtFQVNL49OG7Ssw/woCB30Lvc3QvCoXLbKaHkGSjVT+LRfvseZrQNZszEwbC7iWJ
8gO6vG/j51oyrBnkh7MaJMwAJKVkihQWjUJDusIkdnyv81URmGtTb+0fwszHJAK+
oTDGAuF+TSWWgKd56O9OfyKABCP9m6vCRNQB6acMD4fEeFYGu92fNKFrPbhetILz
v6nqwVo1oX0krbh5TPPI5zqWlQHm3JfWbdztvVXDg7RfNRwFe3ECmk3Wb0Fj9WGC
yUeEeAWxERK0rBhqt7jXEwK0hxc7cE0i7TwEioBvm+ZPS2kVS+sSHG5ptcCov0Zg
qI5P2dET22OTVcKgnsr6bsJSGHgoUC/nlP/4WtH9wPNkQAqQu4gNI31imIVYhzje
KAX858FrOg/7bZ6W/gSOST30blsVzHGQNhFuMjVvg3Y9TLSZgGYqkw1vr9Resjin
HiHgfOBJUblRBjXGv28XF2SuzsNEQ63Mc2UrrMSpRDI9L9NhzSW32Iv2xKBT0JWR
0RWNQqsrjSnEFPtJz6ym+xePkYOvylKXUy5dQArBhq85fD8W4h21/bUacK2j8IIC
LrSqFqKnHHcUPYh2bB52KvQWLCEbkMQ89H8h9DG/UY5sHAiPBZgo3vaZ07JKjKmA
LlbZOL3VN2rTuHgmEEBwA/beaUqZLl6wRSnVy1jD5CKPnaDkMY13BUBZWa50aDT6
ku/Qut1ZIkyKvQcjRiU5uU7KXB+W7ocrHT8dIc8bGe1YnzU1ByhuBzacBpDdWheX
iGfwKbfXh62mmOonfPdomOECtmIWNLhmIPU7l+GOqwxGOowenAM2rh+HbEr8obvZ
CobQBbBX//kRg5TKO992JE5x1A4OWXbdTRecka11UXcl/r+1tqnX1drPJangB96O
u1fXxNJnh56I4xErWsYgS4bHRQPXpRtKTdTDPzkPRywZgY88GX1lXmy7EB2vP9R1
iuM1M1YDU4GVChFTEbVghRP8Etrct4WcfY8Mnai+VJLLlRKVWFgBGvXgCTIcZ+jd
5pzcLnSsqUGY4LfSGmalRUQg8XuLp9fxAx62gOlBjXYJx+dGKD+LftL2tiWZXhXs
Ual5cNx6N5O1WQqbp98A0DyrLo8yRtjh7/bRM2aOlrf4P2DEnS81v+iAIZ7ai4kg
jkisGvlJK4i/eXQiFpo1kIx6hpURzGHv3cYomAEZ+zb67er4SMzaMbYPAUXLS3kd
c6FVtIcbCn8KaeUuni6eCH5ZBoNGioHE9xwYGhggS2NGkUzsxq0ugGKUQPs97U4Z
EyaPlUWlxq4bZlrNLaLp26lMn3nRXL9YBIDaS8GNbfQdqVAOinhqKoBvwV7oDxjQ
QAoSkOTn9nHLL/XzbTkyweT5zaSXNoaXZFSs0u0aqoUqcBuLDbyerqKTLnYskg4W
f7C2S1MF3+MQ15AFkf04l6vnuAIwjI9eKzcuDCpUDlQ+LYeHxAtCn1fLQcENY9oM
tPCShobnHEBsLfYt3eCdU7KUL/3Wz3+yLnchBpM9ok1maTokkO2rHxDfIItsbScU
GgkHtNvqbU+2SsjY33fdmj3GBmXyyPKTAinuvOlovC3bIhatIu9S16lYEJsgPQrI
Eod0u1PYvt2MFMN51z4iAyVrUsy88Fkdhom3mghmbxMS2U2X29oq5vervYlfGy1H
z4xlSQQ4eHsfoDe11BYB/bABoxZHtXvMMChPCp4okWLcyVkQupCWoz8Y0rb0WY+5
SJX390Q9oaMyI3lm2L/N13GMRQ0oK8eCJ8jL0+B78AqoSJjpFun8a77XpYadh+YE
uy7fmiYznGL7fL+i32w1kQUxE0sXhfQxfI/yQUM2NRDDFIOSn31Yf6Rw0tJ14BSo
lQ6JMqaXvCMLJEFEgcRsHANs8vHlvpW8ybx7sWXIk1rHVOleCwDR3A+Ovlnoa04T
ehEk9Algg96Ha6ZZCVLhmyPopT1sCXzimnh1h5fm51FP9SbsyyCAfiXMwuihqybM
d14zxzaPkCztHpu+1GMMW+UH/bG9PNn0p9w2nAvp5gQDgWZamql0vCwwse0aIaFV
yrtADrqiaW8JhrXvK0LCYYozKaSWAp6NCt8gcBQmh/WIpO136sVtHK7tu3/Q9T0M
RuZAFysRcS6CqR/TctINghNFHll2UDtXNpzxaWt6cDSG+S+d2FzYfB2XUKYqqKVO
prTIaO/0tei8Ri1DKEuWXTIR5Ys4OIExYbNoP63xT79Hq8xq8xolA+DPN6NpY6+Q
5CkVhoM8CBvn0EDWBPXnsQ64zC/pWlNqPDrKHdsjdSDwXIqt3VDmCsrv8w6ClxN4
Ty57c2llPuwMNXv1YhQ9e8iGYdRFxM+gIA+ZPiOxUUwLbMEM9cqv9jDA34nAOhru
om4ljZI+1Yvv4A4rwKt9DLT4MtXaT6cL9/a9GMYdT71+XD0U2ggA81CCqfFtDx18
av8exaOk15rqO4yePfyIJCgC8xyW4GRdajH9RHjSACB37keUcUACuRmEU/dwqlXD
2B2PYZJdPIutk9+0eHqWwhPJ7NwGrwI7Aie/Ura+z9+xZwCOvjvAqHT0F2qdrcIc
66+KAGsz/HMFWOTHBNYL1PbEM1jecDYHA9hrQTQlId1i9JjzCmx0Byx3ihEUmihh
SU8YorIUjfRhe5u8Cnp6cvLhoqVNpsd7Jh6c9CdEsgJ5TJWkauurDYcv5bsmY9cI
iKGmqMhAdXY6pRhZ+xvI8P9LbFBGruqbd0PJiNKe5tGwzxFStuhIiFSEUOo1pp6A
rL9uwPOdg6uTNNhnEzXXlXG+NiLB2KEh0sNkb4J+k1Bi6fzBJUc4NYVkzZ2ho++R
rD85OBSc4r244MwDY8Y2+xI1257DJPsBgHAaBvcfF0EFxS06Nr1L84iCsDKsUxhP
3l+VRaHZOq+WhJKRy2T8cZPcgZ9rRZ801PPV243XOJMfdZO3NDh5nuW5soxzWe1/
9+zoCuohWpf72OAQYHVlQTc37+86J90gbFh+Z+ZZxdfYW8lonmAbMYBi2LC3mA/r
UhlARMHt7OLs3AEcFMGVsiW2Y59Em7JJce5Vb2MNG4m6friGiU8Y9b3TL+UWwssM
R9tLF2zP5XlKF9RoGWjq7h1rxVlpidoZxu1Bri3fOHL5dkvE/qV/I7lR5DxveGcf
QUEvGb6bCH2XNrsItgrpNbktYwnNDdTNDda7Dt7cAIpmiyti7koAhcbIc1g+UQeA
VGHsozVJXpRW0tJLveLLf/5/Qj6k8uo9NvikFH/4/hEoVGSJ80afrhQh/hk0AZ5a
16nkMLd26Pszh72bmd+6lVnFc9YWYyyMvDb0ncpSJQ4O+mh17N5sEEbH5ZcCJK2Y
ysj52WexJyDiOn8lIx3kxqlCxEE0V3zsf9/h4mBnhmXZWsjvb9lWRqPWT3pSuonX
m1MfiT+0YOXXInE6sD/sCPWkAXd61cWMAGfUgNrvwQ6VSFao4NGjKp5WZ6hL0iOa
C52JYaLIeg2glzKuC4/0RYYwkYgB8vv2rEwv3SUpeIId3Osj7U/J5MBH4gGfon0x
tC36sotnJivPacGgFGhoDhnpF3LbaaR7XgXcUn7Ojgaz5fh5qU/dHvRtF1rC/124
mwfAC/4DujOyivlkg13L41ob4K+a5Y0Cb18AfjoiJQuXdcJHPCIrI6j1kK7AKqQ+
EuoS7VglFbT2P+/eAqlKXfj27le2Gd8bdvxa5PyFDNqrA8xrlF8o/6Y4oRuIM+S9
1BtUlcEseB4iQBGVxUFHN+c6qvvm3qNmyKyoxH3330iUP+zeQJlfOIhqnOkZsrjE
OZgxAlhgu3/2Rur8TNa/KJo9RQQ1Ob5IZD51P5x7QmgSKcDYE6rAg9a436e+N8fP
vu1nYDtk8c41Jf55NYh4tOgJdoncgEjqVnPZtNGmT/r5ASD81bolrqzdspWWe9nC
S4z3XtBAUT5l+6WslS2pH9S/kU25w83stj80IUpUf6PzMJiNMeof3pJH2Q/1qaZd
03v/lHeBIOKI8n/3dwwaaHTQb7niLscswpb5ySfNwSmKqfSOKUMNXr05V/AKHxKg
L5vhLmkYn1CWwUXYUDEIRIdxCMBEDalhPbFeGbdJgH8K8Jx8D9SFu2MuGQMz3+tz
+yeuVQT7cuSuz61Yb2FTWeeXODPNBic+EwlMrPfTwytTv1oV/AR1ISRQHMS/m2+Z
C8zB+YBnkc5qA4/4T3XvS5f4N7RJQ7g9zhDCY5YEowVRrOaQa4EztHXdEyLjWO+t
IGnFoFGY5ZII+HMkm/IAKFZzKuee4l9PbQhV3JQtVwYS851xdMOHC9kH/tM/lNk0
ZuKEEHCFlZEIObrv//vj1igLzlPOPdhZOOwMrgzF/XqF+wA5zF4LzkVlR8iNvVVM
VumuTD9PM+VJnuWpPTTj/Ih8dwfg0IOykAy81xEWW+wNdC8fubvFjiokREyDvMdj
1nCP2tVBirXIZN1X6j6ThTfpi1oVoaC4VfwSZ6mkZsXZJU5kl4hL5heG66TnUBwO
OhSZcTZKN1tq4Xng0+XfmKk81kvuMRU4hG/MwgrZytSLWbeXPsqYITvY4+F2lN4l
A8lwQ//7xiqnU4yHoEor2cuUQ5/c8Hq2bxgrkDOwVda/QpbpXA3/e16p17PBvoSq
Qe4hJwot+19KELxcXIx7gNfRB4HDIdCwdY604MjoazW0SyjEcbuCji/EwNsT+y+5
USTkEYY2bkj0XUB0wp6tG+hvGQ+snF9pjXlSo6+8IO39Tuz+lTegX5qqL+cUAbcI
zSybPzkleFc+QmM7vkQdOjmyJXfNqa3d/niN4Ss6klklxzMMhcE4Mr0dcl644A15
Matnp0CqiBzUSjuRTczOpK3XFPD7wPj0zMY0Rplg2gRjE65BRpBNEWQe7+gYK2k2
TxQx/PKwzCrkgXV/4ec30DJNE2LjXmdZ1tFkunZPDn2baRVCJusWG4y1/UE8iE6j
qOUiw582gx4g6Rud0cTp3jzpWtYinjzRoROhQ66BoC4LTgY4+zte/qCx70iUqyQS
hp24HlesO01vVGrfCjgMGIob5hpoPyhOClnhndlhC6rodjzI6AMQ8Kj9oZyyoI0f
1DnGtfAnuQrzNdcjzfkAraF3vsxEeVroCqJvB0qhTZgD74SZVE7+gseiw9XZd2ij
xAGwMQnYtyaw5GuAiHBa7nJc1gXqqU5kRYEgjIRY+6P+c33w8Ei9u2kcZhj0vPFM
WfUrnnBEWWFXmVUtBqJzGvC90YsMW7mmP4k3sT7b9m2qin1uenuyt8LZFp220mw5
Sc6pRealHszn7kBmoO5M7eJlqLZzNhe21J9E/LsZczVtOiWVyUBruYNa0gvdL2aT
uOpgVl2bz/VnIFxKWVv57uR83restMtLkt1i6O10sdsNrNDTMrgq8zvIchfHCl7C
dILCoEaRZX1o0XpxLknEzGBeZ1woRpRf1O3FzZAsM77MN/jiODbOdXzyBprd4WLh
bM9bZk6O61jy1T1nzDmGJ3uSuv95V2mF0xCkm/32tRXQLJ+ALT4aRZZb0btYVuAk
eoMT/ciGFyX6O4rJszacr5nkhA8lHm3KD6hpVXL2cdwHyeK1miZT98uWVTDVe+nD
BWyWzfSQh1gg2Gpz/J7AvZqsEFf1zggPccyyCGpSHZSgsH1BkS4whhb86FHucs/M
LJiubKBNlHfA3qdqWBC/BiSw3FOcBlhXEc+sRTPCA9JMpR0puqBfjrA3HWPNY0ZK
Zn12/9XBN2C3dzIMG7FALFNpMQBuGSHDd1Qq9UWGmXxx9JEEtorQsLkVxCrdapyP
0BjyNgoU+R4CW+Ut5WYmJA3U3S189p7S2o6a/qMP4VrsJFaP2jufoz7uRsVzRB9C
fYgrb59FVnjJtDpv0wgyKXD/o/xWICkZAbpfhp81hiTBgKsbyUx1stTpMkyyGQW9
VNxl1nSED+fsBWQ5vw2smA5qC/FuaLaRNdjAHBkddUnKHaB4MLDSBgZeejd0GbNv
rsks1BheZWFSJwVrMVn/DxGoGTZlAqquFOY2fophl+my5D+9aJi+vOyOTy29R+aG
0JyWX8fVeLBBeqBd5ps6IMFpTi/mShAprBSFaN//vBFUiDepg6AztxYJJb2JA2SV
m94e5AsQgHI09m1GwnLS5WyAETi/npLTWEGchs0NpVHGayMGgzRir4OtF5uJXS7m
Vjihzbl98EB6TSUQShEkWwtssxKu5DCPUoKOTMrpZGj1YKxf9YH72B2bNf+/qm+t
o2Ut2rqDQEanggEcLdK+Rd28dfoqyeCMRD9U8RG9/4T/P6Q/XJPV79XQyVSIeEBi
Th74khSs6lnN78SrQhWhDtlpJwe7sXvRvldJtDd/Mt6dtOau9AYG1ysmB3Mhwhyo
phlIq1q+cmV9zm6jInGILIzZFT/skBEmYCn8/l8kzDAvmIOjZ+PEuZPYv3aiPSfi
SuWb7R+ur09DORWnz0JjxOucvbGxYqiw2HUi5tY9Ojso//J1R5CBaRxJPaSwZAII
YJ/yiOPxvC6tHI43VyMOalcKPEMro/5yHtAcErlT0Uc7T9ImVCEjnD8iVmqmSpuw
dnW2u46cAmEzVvQs/I+qZnM5zfmVj0Ql2gTSYpJpNgTu90SeMGHXFOZTWs2Al3sP
yzH/P670jv5+1TS/WaEHeSqNDRi9k/45pm6yGGt6wc/Sm4n7wJ5nE11ljVMNnSI1
fsZH1RKnamKRI3athZdyI+S2LC9AWqpLAm4iVYiKan15E92GlS4vwgL/LDwdieNz
i4+lYqlNTmd4C0SXfKWTLSWafJ4Boc+kTf+22LgpjQIXf/DEaP7GJLSiiwu18nYD
p3cixqAeqb9KtmaiJw1EKMBkCK315ecJAraMKlPzkZgiHko2H653zKj6qCkh13xZ
1wn9yKSVkqfq/WqwxkQqn2+BHE/OAnCcblgEc19rfJQFGRpH42XgaNO1DpEcOmUv
kvrdQF8O6dyJp3dw/BMsvby3A+a5BZjnLwr5zfvVnmAEDnK/Q12hk+auQskn9SqA
qDEz6qa7iijcUkETys5Tq7LpY7gKAHEWZkQhoKZuay+zcUZd+j/bt2FFbbJFfkvV
13Aj7WAqa4survkXwIjZN3FHZV6utQYVzJp+Hj5EJMlQjRu9YRmlJdYz80OcKG+j
MK/1Gj62x4Vw4eAdF+5hJ76tguWmEImJ3DnauR4gYL5Vc5PSFHGxo5W90b3QZHyj
a6t6BpjgCy4khVoNEmK0uytDOpyXGF+BpiDecTq21Z7Yh9GFJM2ix9Pma1agdap5
cvMAf7Wkgsak6Sdag0veuzQLtYf1/dALWNHT/bRpOYL5jg8kuKZV/+GVrh3XV14k
fvREZyq5QjeCL1LatzJsoSCVrtmkxj4FqknUGtkQplXAjapFI0d57lARybkxXYXT
6gvnN/xydW8qCzXuA1tm6SQk5Z9HaTZ1smi8da1q4Znuua1V5+c8f8zxyaQupYkX
BpYmkxQ1oNsiZd0LoQcp24RUUyKbWQm++lsP7Sh0svT5rC+b4asc0kYsZRDhMY3Q
3g6rTC9y0K8/ZaTSDITikWoUXOXew3E9cBMKsigKPQ/lME1dRNKzEXqTPEgskKX+
QlF9of7CQx9fhlbxYcB4MYWY2EitRA45GTIRLNA5bmiRHGCTAiBLazRhfl9WZXz8
Pge4Lo2/SrWzuKGnERF8UR8XvQGHpiP1nm8Cswmnfu20aejXczHnlQuc7DylkeRF
AaYQmqwsWJNX6Wad2RY1sBzAZVsdMQkx4rFaX3x9YbJnWVXNVUrKvNdaJYrtuGOu
Y3Ko83cIf7QXdS75m8fKhWuGMbpj0fmNG4E5sh4YThGSE7KueZ2N7zuniT8tj8Lw
5966tkq+He6K23gaaCS5IvvXXZc8Lxo7AeSVeqFRCzRFKI9NvGvzv3VWSWqYSzby
hIc9UzYNArBcPsVFG5X5E/2Tm+di6GFrXnf0swMd14y1C82dQspFIxBw0hMufmDN
NZjc8hIlN5Az+t0SaY9Zwn0EFElViolGOfqyyaIbLcl+e/1kCUTOLS007cgMpTZZ
qy+WRLRFMgmMiYJk+8LCgfwHDLfjsPsFGZfHiK8Yg/80SRB7oyqM9kuM4NdA0Cju
d0KSbm1ZwkUgdH1iaMill43//NDP3J0bY6sVVAN1jW4Tno4/7udt5jgzsYo4Yd/c
7W0d/SH6pEf0d2F+7kE8ASiVyMPfzlbZcff2SEUWUJMoCwTj+9GTJ2Pw0N2nKDaM
shJp6JgD89Yd76mmDgNqxR1cwaaqKNpJOci9rwgV/topjyoZJTq1r49//0baA9QQ
ckY6GcnN3e6dRRJQKwAjPHAwwkby55GlSPilCa2sTShtoqTxmik2PWmgrw2AbDF9
vM6C8D2SDwZq68ZuMG3YQe9Af6cuq6SyYM/6U7ioVGxLqpZrD50zQ0jHfPciB5+W
Ea3LYTVRqiBOgoDMbPZ42UNHbl+nN5+7FvsDIswsaRdrEW3XYmMoxFJliI3+6lbf
h/vPW498HfQxbPNcPlqR5UPera0NbTQaLFLtP+Wpa3JBw3RDhZ2zRBmNDAcD1E+x
WV/qF5wyV548whxKvn7X4z18PUOe+eERGoebcJlBkfEL+w3+caXObfVQCm+JK1fQ
VVH+q9vlZxJXNDf1XP9WZbc7u7HiQtSYwugw4f+FjtS8LXaDU/foBHs6jlUTbYwQ
6Jdoxb5WyIZrbXAK/ilrJhCETmODIzSLe2GAS7KdGnnPEvobke1H0+9vpGUE7gZ4
KHGVk9NLedi/wlIcaxYvm2QN1Tvta693YVIrdfXYG7szToCKyfd1FjxaWr8/+7j9
3rLekwcu/HAmDvL9tIuRhuYn1qYFhIffqxq+qT1+YMuehX9QAmPAT6p+F7Lj20Pe
JHJGVon8XGBRjmtHQ78TG8qRCYFFCnSrMKZCDiazWV1jP33PTBc/A/bYUbebNJ5b
TMzwDEILeyeozQ0TTJC5S+X8k7o9qE6uYINXzCSvhh/Zn72HUWg1RgOf+AtXRodW
nN7HpqOm0nYwL1u1qAVzNsnprl/u4XXq2/ErRMmdSqKqy80v68J4oXaRwuZXX9YG
O+G5YTYUPHvZV0/BcqmL+7w3qOjsSd8dy5h9CS9b9uz8QAAn5soM2/cUR3kyUkbh
XblNgWD4L4zllT6owy788vHJ1CsqOj+3tAfb46URwblAsPoLY9h1gIbbGH7opGFX
RrmhF7LSkrbZikL2U4Oyeml6nagcnWGUbX1hD4NEUqHss/IgPqQmjJlp/4iFLBEN
MgIU2GG7DjmkDO5Hoow9RnSN7PoDyhf6XkM0VfaU4zw2uZApeRIhRdkIB/Oiui6b
T5eEzPJUSwqFaDGdSlXKGf2tz3YHB0WNwYTbNe6KvLpleRMZ+9QTYoMK5IHKdBHx
0dqiekiIXb1OxRMLy21QvYLWIv081e6Uq/vlrw1OQLi66ysGtkfQM2HRqDKegvtB
yqoNLSd+IAqNbnWd753iLip1oaldz/2mRO8T0ahy2DmEhUCcP4Ozq67e+O4hP7Zk
4u7HsToTv4tjsqU2YTgxMpYl12Yk4Dtg27ZYbqqqlNhTH6z0Wa1iCuFY0DQ7UWbM
tb3J6Xj73kFWReUEWO8Zhrs5Inj//FE4Pf8CPNkLnRk4UnuJPrx+DJjVuq+zlUWp
tlLakhTWOawsaxNpEmsrZ/3a7/DyFRtEkDGEtxPgVr2qzObcT3aOHjtkzWJ2Suyw
YMHv4xAKZ6DNE2QHUoyZekVjDkrvU6E6tuzEGYQhr/k5IV5heeZ04FYEfeq3N8xV
aVqOZLezWxuqDuDk/aMY99fLKOPBSzp4Qd/PEoPNuOmaKxU52ji/cOisOhu4/vjV
sGxx17oEC5PMPjkRJbB50Kv9Vr68DHXojNbybH3hFa0cld4nwgzui9wAITm/PlkY
PN/CyRgv0QsueUOta96Tcv14xo6mhthk0PCEPgPXZ+o8EPm1mT7pLJ0nWsjJiwF1
xdTA69PHQmF+ON5fHEP4dSA0Z49N0QAzfLwsmrnsjPDSHB7kydGVn8OuCI26FVnm
8YElF4hPokFH/ydBhmLfYryW7J2oMnNBBmlQPX+DRaIMWZe6FsmW4JlI7S7hE8Tp
vjYb0l5f97Qcd6BAfPwSraC3lbR3WluY/euPVnHbGFMdQe5tM98KRNd2030990/K
1e2jxL+/TQ3VtDCuEIJuwGHUO6y6oi/UGDpQ4bu2uVX+Ms59JuIJbbEGgFnQFCa9
P5R764iv3L/4NlAYNHw0fu3hRH9+pCu5USq2ky2NlUV7vHqJRyCb5A5SfWveT+49
DVeifQwOgAm6xv99/aaawzhOsbCBcGwZmKlai09Eczf94/yvgY1wTOVK9Wo8J3an
YaPcoBIjlxbiIvVN5/RDuF7fyDBYqDXagqa9U0n01LO2sqUlZRi4k2ljJng8LpCF
z/xPM6ZvnNPAzSnsXxdED6UdB3DJFDZ7luyGwftZqxR92nrsAc+whvFYIJIj1OYj
X+ZmxWZePKkChjrezFkZ2hzEZA3QgIMTpmUDjGoTFqHQCMOBaa5+tidMaVOSbI3s
0rn1SvUg7scDH1vP1E0XJbwjb/cEZ6pSLkZpchJSHEwyBGNOH2J+FrtZ2BGw8udH
mbihxVvtAHi2gysdPlXE47MEKdt0eo9J6nJHa9YzIHmx35yTqS+bR3mgmK480sgc
MRqi4Q1uTol0tlncXahGZsB4MyzwezFUSteoAIKhvQNkygvfNHU9k7F7JMZ5Zyfb
18r5EmTu4K6jMGTBJaBnaXtaVwmgPNhtidkS9Tk+1yBxVtdUPYlz438ML0luQZtL
32Y+LYY6BmsGxZJLeYCMthD4UHi6ALGEdi77mcQLhB5xtpLNOu//3MLmVA/Cxb5K
UQ+LwcF/P16HV3/QbfybG46Rz0Pvn/TSP/dnRyMC3YgMAoR1x11u9TiVXz91/l2M
KG2c++AAcKmESd86ZI471lB0uMprEi7dgu/dPKCa0j3cXkVhE1SiCkOyb2crelqL
Qm6xM9HeNV43+MqGn14TK7+EBHKzehenhAlTt4cV8w0BJuI+V3UxgoKCbqJzJD7a
muRdPZHXQ47npMr+IwNODKbiB5rYWKGiAjzgCpRexig9WoAi6vJv5L7K+rlamsiA
O/QX8vkG+d2beDdFZE3DrhHxv5d5weEPzc3xAaI6S3IGRGbFNBJc1b0ABfnVEoAl
jxfgXdXjcL52Z0zKUJZQO021tJ9N4168aEno/7jFc9cdaTUZXfal+9UaNH1oHg6F
1ykNX/9JSZxthxNsgWsM6iIHkgMPCIDMajPDzLFzDH3JC3EJ5LKfIRdT1s/MDYse
SfmDFvzeTrcHFEWWo7TDdyYEZkjdDquFeOTQ7eSy2hNxjYWj7gAM6R9WjqfVa3V+
NTAbN425+aNsq8e332MFnUfkB9vUW2+CG5x9r0L+x6lcntujnMsFUT2Oku9HNhwL
AQWqveizmzeqzv910nK/5F6SZBktc78xMYtzDGqAESWCZ06KHJZ8h+82G+gwWPze
p+QPhm+54s9MCp14iYcgnDlXiMgYIFgHU18g5iOVnOH6Kh/wsyrfZFkGfkG63QDP
0kSrSJIoxUNfhg/DdV1HsN2pv55h/YaIdxOgCAL/qq6UqPeikY3O1l6/EQXCOyWu
QFfVKQ8G0MpTq6ouzxi+XUmTdo552FpxjiqGKTun6/KgOmd4SquqeDVCfL8ERP8p
IDqrnoXcABLBq/eYorn4vfhLPApIveru/w05k0HeeltJhFAgv+hiqVYZrtnTPO+E
bxxsHPCC4B95mZJTUFcHlo2D1pEwVVt4lvEJrFCyAVisMpWTdbwz8GxPGROSHew4
fKFQiOZ06hC7xgcAPpVGAG3LfIm4WUwkryQA4opcpbU46beIrsOGw5LAZ3LM6aAa
2fla0AP3zOxn7nSh24MGQKk1FzwCHYVdKIhzJE/0K5TYLdXO+WFvkLcisqLWlN28
Z4N1+PDL0RuhXJeh0gqCs51tjEG7z5veRk1SJbCrW9B3p0wFeSYW4QUylKdOlQpl
8gHARbWTt/wTOyS2nwXVrrAax+u7OPJzmrFjMfYW08aND0byfX4HXDHNXWVxPVhP
i5E4KfYi0pIAhtXW17DbpNWzALEA0EmVJDOsqc8A5Ga7TTmAOpgeoJFkPZAc+ZGK
XxZ0Xjzxh6VHGc2MZU08UXWFWbl3Ah7yONAG4qo43WRyIg364KCgSAR/8B4P1z3D
RiAMvdzya9wqjlXmLQ4LIGt+j5q6m80CXwxN+R059K+IBbYFWZIvcdHEgZbuP+MS
GyTzHSX8aPFL2qvSR/0P7DZrwUFFfScDVfHH6O5pR1jrSvVabNFn8fZHSsswUidn
iltE7vWQbiQk7Rltc632VPzxkqkIImOQp3A/Gsk/TCKfrJDNjHsdxdIWvNLVka/z
hKrzrShxf5aiQqUnRWagLS2bD28IHtmd9lO7OkWZ7u8bJIMDD4fsOAM/N/83saoL
2n4veJ+JfVLA6XA6Un7axMjIUIGS0vvEtRH5F9w7Cgg8O0zhuDfrjeLE96Q82JGt
whecbCTfaXyd1rCJkJc2cxLBGA1FBTE9bLKbTj3Ui78t99tyMf6ss2QnDfMypCaV
sRiZGcIlHAUfFBK3ODalVAHIK+TQRFJeMj+8G3xDP9eQTrXzVSKEb7tdJqKr2M85
j12crWoDQl/bcq6WPa5qU0NDIunR3nZxMUfjgM2mrmpih9fUu1OyxIk3h8kKUxIE
xxbKswsofJZDwpDNiBxV6lNcs6PzT5GohDCU/8zzSh2FhChOfwIgvUeip2GC248u
C9saWYtqwe/OwvCt5tyZpEayksk3VLbBybZ5NA8sbJVGBpgxnlomQdd7xSGcEqvs
SDWxxmQkTCaU6KLNegNblvKoMfbbRRIeuvoSaTUdmfsTNjoDvgCtjg6TYvU6HoXe
B1LxQiyw64RyT25iEjmkx9FNgw9O+Sv8eVhABBQeA70SuoWdWAPJAargK5n/ui6t
tp5Hp4g0wRDvSMTc/camCmLV8odY9eUWHhXXe8HP9DXtit5yW86YH3L9W9242xTz
/mGnsD2+ZUzqPTli+ExFAZx/fp1MBRw7cg+wbj3oAEah8EILAQkUfw28dycT0NX2
PjVQUunX9jN3cE+aZYit0lBLzelZU2BJ/2ItO/ro2DqUSvc7eRaiCVeZhNmuzYXY
7xe98qxNZ17ZmpGdaCSegv+xPgZqyjllkRIphTjWwWKw+pljN0ryiWJZTyIv6oSN
sZG6rh71w6MI0mWRbKwtcbzPw77kmqaulBugptP95yqL3bTi9T4U1DR38ceFsKrI
GzSEodtj4AGOnXdE1wsTfl4denhdqQyqMuFhrTqvp1BiYYNi7dDXBHJ4Lx0dH1wi
7SgsIzL5tDf/a1AViuaYf1fZYho9C0ED0Y9cgzEfkpN6urcSU1RDncqDJtU0a6Gu
JxKnOheL2uhB60gNIqcmXLpGVRkXD1qVwaDn8Kp5bxrcGCljdiHIkL5AhsH0DvlW
+oO6bRP+rkeUrDHvmx5OgiR6hipw/4kBTQX2T8tFN6LlyXQtvCsqaZ6V9271Z59K
+7bV88pI0ap8r4qQhcOzEjgTASXr3bgelYXc5k/Cwp7kBibz/dddAlke1chGugRP
n6om5DFmKmOh9h8Q7w98ABhm+Ih8a3HaZviGUjllsWyDSEPbwEtOAl+Wv1hmE45J
XHOQCZdhNYjW3mb0fPf52zQjm3fcjyLfvNLH0joCYIQfMPIQvCmtsJn2pytHZIRw
F/AwA2x80tMe5U9vsbZVmccPc2pmfREZMLQkZP1zXc8/yl+47uXhgSeXygCu5yi1
ThXyF4k4Rq7oWyfUvmSqAlpKU+M6jR0xYvUQ6ELtDgCp+8xr5UPRr3ai+0uJqVmT
viq+FioRL9Uvi1UNWy8A5/46OjS+zVUa9IFq7lyjT5AQazdDPqqhahbohVXst/6e
rPgpTFUVI5XVZEHea8M03UHFY20fhSJomtWhWw3G0peIO51Wug6axdixT1znZ1K9
jVL4HqRJ+u1Xxd7+rOS7YcRIcie19as2LwGHAxjNnxIP0WWMzszZ1NOGVlDc/vrD
WIRANIItgP9OUYWWY7Z9AhNy4f31PRXalcYPVy1FeE9rHLqP4DV7GqpZmCrkQC/r
QpnyQRa1L0NwXpAzJUjN8g4/So51dnJhpwV+vtWctGDw3zXBM7QjIRhWE9AR9SN8
hGadXFU3Av4qvuJrFmYgIy4sKQBFM20TKpmIuB3DhmkHaUpoA8Pf3r0tTqfAaaow
w9gv9m7lOrGeCEZBG3lukl0wQq73MPenjYLtUauImg0oR4bUWd0I9WfVvpZfd4hX
oW6cZ0D++EK9ArZFL+4bsysOZJm2T25QslEvnd0uhlSLIcYSoHDbBc4yXkLJKVwh
I9NCIWKDGWlxbZWBNHyNNNJsccJ2WnKcgu7+woZtE+CWjZFClWDBZVlUwVBdy76T
MaIKMOCbtOicDMousybN2WCuNC+UX5t0k9fl6h6JRxBGEn1gsPXPobibwQM/shnm
uj9OGyE+SFkqDv5Kvucv8L9h5zO0tuYpEzSZLLHtF4b4pAK/OA+4MSMILXv7KNSI
s0M7s9DKadkD+UCogt/zJws6LVyZnb74KbFICFaCkOziRtwTsxzfsz5DH75jrT1g
Q2N57Kl+HY1LeQCBcdmovVUxKHiJ0Jhbo6TKkiw5Lm8CFPxPgpaVppV83qD7kH/5
5BYi8gwzwtWF8k56gtpFAajlZtqdTi2Kl5xpAPGw2ABnyrLfz7ttUBK007wZofY7
qUnh2/IMMU3spaqhQL2AAKH0r154X020Lrhmu1uTr6reGz0JHcoPGebAMY/wHJdK
J1MDNpNOtZ994MFRvandRU3GKRSZIV38K8zPq9FlW3WP+dXdocsr2YBWudvNzkQV
oETWx1c+vYqmEWH5y2y5WmRivlmQQ1kepm/KoHzhNWO/OQYQWUQG1cmcVHH1Ti0j
dr8YQCowTwaaiIKaK/hdpuSZd0ciXL0Xz/7HLcguBxbEujkWQ/9BXfeYOHTXeUQi
bgNzoYL/IjcIPd1Zha4v1TsucVUgv/MdAq4C7x4dOZ43D5YCYYnPuIoO/8ztGZEy
ftDIU7O85LKiRZ9VWqUuVOsCdOcjSHivK5mT1U2r7QFZ4saR52cv5Z0sGeiZw/EC
OChSPUwpmEhMjIwc+vvaRRmECs5GVWFB6v0DHPtF4fUPKgWwSTNx6DlDTMSH5TUk
qpD0rpVik2fPC7lRCvGvkBTcNSmRDKBep1L2kA24ja+2WuXkvBpLpxQKYLHnOP+I
MYxRQk5czH1H3tzP3JtSnCF9lFJNqy9iAjSo5+CeVbab03PoKvFVpGGBqrXUTnDO
wU5X2aGA2SmQOFbI87Q/pTgFRFetX9z6WYD4y8Ki4BObjW0BCr+2YgxuRm1ggGLp
yPoF+Ah9xYhbXo3wCUYwHolggmG8O6gowJnMyOn3JvnJmmLJokUd0u26O0tdXbyA
7BKMX+nov82yPzVRC29UpkSmvfqqXQ8U2FOy0e0fUzju0SM6goehvtNNVc9ikIOR
oP9DCUdfJzlBh3k0xo2EI7AYKuXZBZGcQERwB7o4M9LVOI+6pIHbllr2iLD0GT4u
b5WbRqA8Lq3BPjUlcsaCGxLHCLyjr2LZ/OeSRlIRd6IB9XS9iEcQgmTAnsmfRgLA
73wTiOgFdqMFqLrZqqmcBNJ26g6d1T7D0Rue4jmpZCLwHGGa5KUowXnr15G+QaM9
QFQfWclw/M88UwuqYnwuZczOrjn3VtaL7pJFMBGjrcclE8ya8gCRwlrTFNJBUZYQ
5/yPYF3SX4Kzx/JljAD2Yvuz48pUmUL+n3f9XDs/ndcoztF+LzyqDFm7ql4X8YTe
j78xw2mnY3tI/FHjLHephFTLR6HD4LbjRJbeClLBTb++xaIwzCKjWiVWYeVXZkt8
oyRdKqzE4HSbylHA+gY14xH4nEwdSsFisLiC/W4Q2Z0ecVGlU2uRWCUwWsTD9Qba
L5KQdtq3BpiSvSMrH2w7IcPgSzjDHvhkl7c+wXqzWPoGPPnQ8i7KxMidaiglnaug
DiYGLtuVQOLLrOuR13E2LafCOsXu7nO3GyaAB80Jbb0M0saGaUBISUX5SlHtGHbU
GEjdgup8QOXv3ho17jELodcMDNuloAi2bDryxQLUM5osfdWAihe8uO2XcoHFqneP
kBLlVxv5zJ2u/V0EwlwV5JSOW9da1oCjcByLFbcRa1s1G19FYUylgKWeiLj7aP07
kAlBuVPRuklkzTFAQe9SsHdH/EtQ8ljeFtRcrHHPfiXxmGlivInHYO1Ec0cEMOEk
1AWOAhVAxaWwtPT4JbXS7Hkpysvzu9Kkxgxw/SAgjQFc1WsnN9pOGuAeF2wsZhtV
g0/y+MrWXudfbte7I40KHGCrYIejnmhjR4Bjs2RCQnRiRWyu9kXupVrKt6CWHtYK
DPaJCM1VMg6NJ/A7ofBn7L+72Fl7XNXK+A5Soblssh4IbKFTWU17J6JdU7DAqk0J
bEzMrv3YeGHDSc/aY2Ro9sMVxXYhK806YJBei8EjAMLd+PLBx6jy1chyV28RUtsO
kwGPe411C2s/4dwKTH1AkNAwA3pj3AzEctW/oNGgpwtoaxYmjruwg+QqDwVEIEbP
QMIRxKlb9bM3jg2JIrjM6tgKTjyYZl8dhqkQdjMiOox/tPV+pkJinHDDKvuSOp+m
vAGhpKF5sl/kvQvcaI6Zk996nsQR9t/za6UILXEHlrC5XTdvkLYMNAx0e2eIqfIW
WM4/5fNIa4C9Ssf4mdnNjWwpZxK5x4MJPkT+2HDmWNaHy2+FNpN9h67O3rx2SBjG
P3MyCF+3a2mwp6ulio4s9dRwYem+1JOuruIpoFGaMCrWo3M7AMs3e5k3L0Y/ghFu
r+lZsLZUDdeHOGYVvzGptp6CuvJSBvSnSddR7SbIq/r3aJVu74cKMl2KtOx73KFU
hZEvQVEn3URaQEx11zWm8QX3ZdUACSxmxREO2rvxe+aMEGucuPBs2J88iw9B3msE
/tmMpmjvZXrftqeUirndoIOvkcMiQk6xvl1MYkQOBrRgOZbgJeo5XLexnEkb6AYh
lo8qbq/NSlplxHdQHnilBUGrIy14qq+wkGkoU7iXD2p3RMNOwr32F4VdhdC3sUh0
kKpPxIuEVvoinjp62R4/guvPegFimeUQdhJ0gD+wStHQ6EE/4Ou+Pg7xakgdGnsQ
NqMz91S+hXxd6HdeFO1mZvGvBpvFtHVMivj9Q0szZ5IHMEh3EHZv8lu0AeWVGtHz
HPPvD5mlsgBjqqXpbtD5tBD9g/e5lhEOe7SQu666mQZBzGAZ6FF3bdosxgyx3kaJ
viKIXqp+u5AUeLAPZRNO/rIjsIN1HSMR+OjvS0g6eucxQqZn7G+eZYWcOPegf8FE
Mf9LtD6YwZtk4kDarH1WNmvP72GSe1BiNAQOGSNzWiAKuiDoTXQjZMyl68lruPS8
o17ZdON9YWM7XeeedPnG+xKBbMiS1r1injnRFVCblRxSn4iOk9gZx9wyhjS8shvp
oWZqmFSK28aFU4W8eCDDkvZOBijxD/mkREKerr90gDyGoJv9FWaJqZVS+QQPZnRF
atvylM5hyg3XnMb6mvVxis687evoaOjAZPWYs0yD3ZsZUMW/JbvIyzgyC2ncaRmV
mouCTLVP6TfBWQmc3HheSZzEcOYLbzfUdU76dwGk6xlSCaGRktLawJeAcv9Qq3xD
Gwx5cWfenVo8ZIIB516N60X4YOnf7pjjx0+ZEDERl6rSfgqk6iKNTqt6g/ryAnqw
1MvP4cRCYfYaWxySrC2U2EYJKyXr/LXobjlRMYWsKmE+IGJv7Gfx3nSYi45lvGqh
yPxcGdCDh78KWCb87IxAYhM3qn6ekIukYjO+glwef8TWd+78yg2Pamn72EqarbaI
BBZffZPxIyjEp0NP6HYjMVRyRjw4YcWMukTzeA3h05wAmAA1vYvJHtpjGhmXBv72
Yo8KT4KquaZrbCxfvkCQO4rpp8j1F8leBk+jWNPG87YFQf87TUS4SG1ojqp+PekU
gAIakEjy++CiDpfVvbdzjXGqjVYiaF8dFIDpQwRsaKvZrjCFi5F8kuJKcFk/UVWf
rnOF2p4UYPyyykEP1hfj8NaoNYu/uqHMNMER5GK8MRLo/M6b5cm/Lmr9xaVMmKeW
BAWMTiH385gDjjbe8SWuF4BaxUmFm1FzQILtLQOGGLzVKfe/jxLLj1vLnsVKnL5A
WuDaXizWjiEmGQ+N4xzX8RLww9uLI0lzIPxzccHq6catho/p48hsA+wANgmp6BaY
5rDmLOIBeZDsBS9rwtnKjpbGg1nWMXStYIXoSIgIalLb6VxVQ9yUG/6n4DOgK0FT
/Eze1RlKdpvX999XjVAcHnHfUGFCGq1Y269TMcsGQKsYt+7G+z+qop/AFGJIoUZt
Il3K9njJKkbwt/cBtU2DRvt69xAcTtHxZF+oAIbyQLXbk2pv/C9fYVef07efNNSj
AQQPszrEs1nCjdpufzsFn7nfWvtACK1b+bv0O8srK21V4NPT5aKUM2WhQBk4BrqY
uVY6oSNcIvwsH1lTEeaTl1kf+Ijencbq0PWYcdD84GfAOdDS7jlx8sokPPB7Swu4
WIOCcMP1FDJneTztHER0I4im/4a6ZIFaw+VJBlorvf8TcxsWeytTXblRoE2BWSk2
gqpL7WmVeLTLPu6PW1oNfwi2HzhQ1OYt/WXsArKWu8vKEMSoYOFW33WyuOcMWkGL
xFKbGn6eHKKwwSbsfAJ8cdKGste+gjkmUrpX+QqJ0/VcC32Xb8dqWS+JBNbEOU7P
ayG/Q8jA1upEnIpDn76J1h4xFnQth4KLzIZaQJRrgHMigeRdxUjqF7nHymvopaT0
8QYYVaRoYSjQqJfpRwLgEq2a1KLp3WqY3CMVcbheTl+R1nTzvRKXJ3LxTkH/Y8kg
P8B0GiRfo337ZLniwyBR5Vs0DqBBXeoWIjXDOsjDWpM0hujcDmwewyh4rP7srFbG
URDsTFecpSC0IKceWvjps48uj8nIKKUY6jYqS+UHNdfrWE1K26NttX8fSQMqnNU2
DW4pzWZ3OYnnoLSq+m/sZNIIFIaWIIBmeZLuyJk+8AivCFa09nMFYqxCEcpG6/Yw
fq09u0Pn6nL1f8kN5XsnwvN8vj4L9cD1+Qb9btC2QGow7WbwNg59a0f0eincvlwV
/OmLhGjCg/jwc4KVSTB/quD5N92uEvhMSXpZAHaCqMn/WUj6jEZ7vSj1XjgF9nP3
ZzksM4PZ6uqasgWb64cFvBfpGQ0Ht2k+lB2womvZGJv/w8Vo+p+outcbq1oY0BeC
chvJcQgVztsEftBBc9y/GRiUE1q9FfXSg7q/68gnLIi6NAYWgWOD8VqjmrRWtzvV
PUyqAWDzsV8fvMMt/aiECc1p3LSFABUB37aCBNU8Kkp+tC8ti8d8jwS2FAgmk7j6
3zB/sxPNmjHX3wTDbYWtf27FO0k1BgLdFywLcWSVtq/O8+53AlH+ALEUvQxEdAc3
kcUYlsjdB+oshIBDSGIk6f2EqmJuVxswV2mqmpPW9VQgSs4KA+jbE6HEV00mXRJP
INbWYGnbwtxxBlaJZEtNsP93DzEDhjrnzL9vjA3kqrMryWajie6IC1v/ThgcYzg4
+mEunhZ9WHkP1WIpl3WJLQaV3IyF1qNOD6/sCYjRlAQhGjso3+hU42kfCqLcfSak
gWxvpUioktSB/wRdDAR6WVlUgDDw1jx0RN/FKhd5Jb2oJTTAait+F/+2n494huwm
13/sxqX3FtbTKfi5Z1NwxECCjZ80i8DRvL1bTWt1QOtgaGB52nWR5wUkll1N2dHv
MAxGfOmrujmEeHmJPokkm+oO6QwGsUlE4aJ4pO9+WrsbqvZ+Nqrx9J4oxMgeoMcb
MX3Tc78dq2n3I8XN3LXwnSHeQhbdVapm43CgyCw0uCQg1tuzTpBH+RaXXZi4qFYZ
gUgveAr+8e+WJ0KBshiIbwrqTIanYoLvtsa1GZZ+zaWTxROlsVNtmUirakDCA6uN
nK0MU7719L1FAb2QDNqFixKJ8O3+aBKTPdjEHuILtrZzsyCTtdRCo9kYA/9VkU8j
1mYNRBpwgT6XB4yq5XRKELKxXLs4DutvqAcms1NIwG04EMhUSQBic1aB+yDWwFDF
R9VLN8hMV9OobgK8mm/wool2qqrdtTHG8Dpd8CFNokV2pJE9h5mrViLIKuiURGNw
ExH7WNKpYOMkBsy5eD5v5dc6ZXn8kYofOWZ1n/cDWrbmIfrbBKPQtnVZ7KJdzEet
7oJwggbWDSSHWC++YEHIkrx3bqEdZgHCJvsUF0FLqbJA6NZ4nyoUDRbDvCaf5TKq
EUeVMNPaT96R2/vNMf5Mz4CqD5wIZElnW8vZfB27qvuWDyqYh7WYMrDpJaZlO9hi
qkEd4vnCB28+CVK8zUXOnsCMpA2KZujWi/dqTrsOg+9Zkotbzcv78vAn1uQAoV6E
wujuQjLwYbHTonrKI0DHhuQws8Gfb28vsW6jzTnz5XCvr8rKScjmFD+5EitMT38r
xW1+ORNSRkn/L3sRicKCY/DT8hK+XdLEikK6syEPRP2RsrXlA0nZQdLU6QlA4WNF
86mdEIkNKL2fsGKcrBEZgGSJ16gYGKCGZOWszqX40oNHIp5u8xchdfIaLX04usgT
FSoNHtXJyHC0oHta3CpghXrLOkq/wBGnjp3c5Ejh/esJHABYbq9K2rEz36FoLURj
Bh1kj2OsBOAPBlr876VlxxRqCx6T2f3X/yx5ro73nmTJg1Veo49pgPZML48a9yL/
QJcJoUKwAQ/nreH9q185PD9wAwyEB33JEPFptKcgHlFiS6jz9woymzaJUG7Kw3Uk
LwuYkFpNeTMU3BZgZB1dY1vK1U0g/tWS//SM7atm/qLx76YSAJO87AKahuc82kE3
iHovHDWGbVDmkXpaAmzAuUvX2YNGv9+CdziUqrX7DeZLli/zhn50yZMriy4rCG2O
JYi+q0N+jV9vqSA+p90Ss9khujTBoA/0DueJBqSPchihVVlwEdua1GAqNR0NhuX5
Wxk3bUvx3ajmh+WjBqRF54ULhVAi/ho3vWJJHy8xCnJMewwTGdmPOosId8mHDc82
hyc6QSATKglSlrnXekiJ3Lnmsy7YNxnnlKSAUtI722wX+8VcPLTHxOBF0pss0iiU
1IACrUuEjkJkmhVWbWSpU1b+5kH+IbFQfLstsdmBKbxUgABMgGZs+Dr37Q+BNCz2
i/o7Vw8N6ft+N1xjoEFRna7rhTyrZ6rTGDm6wTr1xbcbF8vkRCM6aEGswAtnVM5d
kTjUepE/F+s4Om5L/QNID8VGY2y0/+EF3+xLYdIRBRlRL8xd4WSwDO6j8LQPKykA
4FoUFH89NeBr9rFGqokRRB5KVaut5ene4JSPnybWfpcu+36N/6Y3C+jOxB1Mrcz/
U/lODsS1dI3lDx3SLQVaFITCAPqQN0wxikBrI/gGtjESNz1eLpjP9kXdhsehjsST
6PmNfi5AWbyJYqmMpyCBSX4RrJA8p7UlqgsPdgC/Ywpv8z/yiFu5DpihbNcoe/Mw
NkP6dBAL0fifCrMq2B9v6g+gezmy+3aYWE2Oqt/OLpgKYHj/KShFS+LKcUCvMtgJ
ncRU6FmrGVSOWGZa9SER8bhkZ6U5Ibq6X3RNtjEsX2cSugsiCtaJGiQJpdiDFJ6Y
YfJeNvh5r940lK62py9Jac9n9YUk2gl+PNKrm64vOcGVLhXB6l1MVTCHHxW/RCCz
iDmi9Jtf9Zp2f9dRhYnPLTQ7ouTdg6vDXDWBqWbfPxSgqBVR4JWlSQCouq/Jl5zL
k+t+COK0rOG4CU4KsqC+cLgIgd6rhlEls/9ZRlfBauTHA8I6nhaUnA2M4h1DE0cj
mlKcbzdMdFemNU7jwmHa0gJ1H61y9FRqUOoCyu/FEuSpzF+6xwy/SfpYXnbE/IAC
ekiqw4fIqX9weAO4qd6fsGUw0fTchwsZbE/MTDoxW25cmNaY3Xwu0YzUxmDRhXxv
QEzoRraE7qTYfHs+3/JZYP6cPCZxqtsEplfVXcAXDPJn+B8EK34qccIm/Qnu9LcZ
yu1oG6tr6IMNcAPg8hgTIiWYadIGzhNIC1xkJ74eiW73NkL+I+9+jYF+gkcPWLJf
3XVvzwHxwZkcdIkKbuxXjwuk6RTmOr9vj6yef68N4cWAwbvrxxsSNqFy8oL16QhX
k4mibWuToY47fTcT+KOgCK5QB9L2u7jtm5t0aNmvz/A5DbhjU8gl+85LX3i5IY0y
KhpuGs3kafNxCS8sF+9KjvPv1oanNKon4E1320YCU2erpafumn6T/WsYAEjqWd5R
W5P87UUJDXnDy5A/egbTrMv56klKL0Qleg10/LG7COt3Iso5oy1GofmbkBjJMrLb
uZpmG36t5i0x2/S3LtqfBHaNquntdXrHK1Wsi8j81WBbshRGpXpyskKEcP5i2EWe
mkW9snVMOnVgL/3jXqIbZSGlsddO8ceXm4cJo3mQ15Ecfn2Ve/6ddYhHMsUm+z+/
zNvoWCB398p0V6m1emcI3YfMj6aaTVMkmmt38D32IxLOGPOwmkNgP9s/UqHbmrQh
qy5/KoXRYtcp2d7ucDwiJq/pUxEz33J615FHLP4zQBAF1C7SaVf+r+COwlJi2Rx2
8kUJtf/Evwhrd8oXbWdsoQm+gtzwvLwfqoIXV8WUSMtCdecC0IEGspxkVm3mVYoF
JwBdnYYuHk8YYVxYfowIoqVPSOt5NnUbg8aSam5j9fjQeH3N88c4hWS4oo5WuPnk
yzGr2+H0qDTfFLBtE26lbpUzpnoaflqnUsVmwD4BV8JQP79ncOy1wcj7VNONqFdi
TN97nwbPri8zRikRzNA9a1o5hZaSH4+SEV2gyWODPM/UhWp1c73yesIUWVeiKgGY
TIk8Aek7eiSMS7d0ffs9Y8p/a9TKq7HxSpeV0mrR1s5ACp0pM3PEqOc2BsWrusDo
22XinY8GMpVhcRgqUnf9AEgeUPpVHcRu953iHEpi6UiN6XLgKQ+1w4WqceqejSfE
16SEjSaixwDcmcH/ZhFM052tEu4BcH5/TcNo2nQ7x04UqYsl9P8RutrKYWARf17L
fBBkercne+rqTmbDDzEsHHJB77im5FmFPhRdTtrbIKpIX8VyUcWILrblXZanGl/T
An8GAd1mRooyarn5XjpxfUxitv8atV0CjGQot3QX1kVcwAS+WVo3/4c7OqaAm46r
rS/lKMlmGnz3XF3QqbtinncsuGq5fnXDOmhy0x2LmqilriG2iRCa+1xsXNjJ+FN8
WUBk4dOzUwIiS32R8rpKQHibg9OP/drmDRvRbjic2GgrpGzwQNVCmfRggzCHhM3z
L92eSZwkRNpMHM8pNHjrSV8tw65SG+vK3LO+yv3d3ARs0rBh4Tb/mznq3gKUsK+z
tW+41aK67aDADJo2Yj1yPKH61vDK+vvm+ZIqUnPAbN0JHysdKzj9IId99O1D8/3+
68GthGDS0eCO4s4vvqYTMiakjrybeSbfSpA0SYg2cuC97EZsd/+qEWlOXKFf4z1B
+2jEW5Xjl2EhiYNIE86sgxHwgNDIN2NIzjfvinkEbWYUOAQ2ZGBMqB7mZlKJyFNM
liw9zxshp1Wd4uNqf1V1KFnIF6SjcnSSrVYI7kpYTalV1x5VGNSpoYHylXrmdFIZ
PgSAq13e/HYF/BGC1C9vjYY0pfSVZC7l+GLIj1N3xUcTnagcDFlYDKEJCRAV7QOw
k6Qq5bWEA1xX99AnlDgCUZNCOSbNOueNSrXnB7MbplDTKh/sKTND6j3mMrRCKTBn
4c1XfxR5IfwILkmbNFzgk2vvRaDLcCJ1O/fQNF4qfCRnaRBihfyDFv44W1LDzbli
1jfi1izh5FOZOhnppyJqQIS64lET85iWFydgg7Q70EENeEDhfMaQxxWdJH2bGVbN
NGTWN7Ed9qi1aZyvMPyvMoVLBv1JEUyMFUjJ3/UT+7nZ+h6P7CDQPAw2oKQqzrg9
quVK6GOGgXhpPVBIMcJHIo3wAkWetbVkqDhN4e0KhjibbZFK3djdn+JKt3lEjUiv
/bL+4btaeJkAB+QBelhE0ELQ5E6K0tzSbzvJNEVwi9l5J/iOmoiGEptPErAL/oNS
WvQDum8InlJa4MBPbrB1o9iR1X4NndWYIBadZROWIfsmIYid1/Vki3HXDL9B0lo5
fjev0Bb460s2L6jlPfk6oY5dYkLiaVrt2Ji1F26zpXVof23GLUnHf1EesdpNW+zO
7Fcxgrm8OA3A0fg9MCNKOlu54RmYy/jSnQxeoAoS0v0nf52eG+3cVINbLWFjhu2X
IaCLNAp03EV8xB9Z9sWXpRziMwqaPC31vgRNTPyxAkIJFS3z4q73S9oC8G3tXoYe
t4MqCNboc75Ne1KyVNkzaH22d7FjI907cmpSGVAh2mCsyPzIovR/NFC+NfK9+0zP
BZWizwCvMNYUrLCgYgUUbftLQAu27Fj6dtoEWS6WDGa9KRR5w53E8vVnEl0jEZm8
SbhxWwWNKF/TuMMJR8vz1fgLRN9SHjoU+kMwKGnhhFdRfdkOMSrboh5d4XrNYKlj
n0EJ59kBdw+Zuc5hPuuv8dD7CznVQLYf2aRObxwuqW260Bd1g/RBzUoAMTqng8WW
ETXGzMjTZYMHqQXaZlZZm86ML0+J1wo+2OYktGqv3kTBnNVmlXIMQhLeIDzlW6ds
HJd01Ha2UyCIHz8BuCu88HQgsadyZbO3E6pizvD5CZ596oGlsf0oAHLI46Fc0jol
Lx832AsaJ7iKaXCBJBwkwpQTYsA7VRq/U09KXQKH+dZ/xst6o+QsppyRQ8Vp3WQY
AkPJJLOCltxpyv+mi1q2hSttOvtVA3Zu9Vf5XBgZMnWJBFr7cZ3SYV/m/sHV5NNV
ndlDoRuDP0TcGRvDMmQvH9i6ZdtY4vJL0alyXyesHCF72Gl8cD2dKBjM3o4OpBxo
EKYOEOF5j3XOyT/LbmScOVZDh6gwy2o0jWQkpvPEq2mtZ1TqtG0Cg/tNNehOFtbm
Sn6WrGnfKsMu4OZvRJ8gcf5pPrmsFQ2nsyvBOQe7dI4RkvmIb/PD0hrmPYiOceu7
J7fPEjrVPj/ERIf/rILqRj2THt2o/MsaQqoBPthpGWKCkG9kK9+O5jFn00VkCP1J
w2ajXg9aXHcB7GjEGeiugggVurNFn+oDZWCDaDGiQ0nNfPwpsZbk9xmV6+q31e1j
Aog3sC9MXfjGS4C5Zpt7uhaDmdIqcqv5EHKIxBTLzCdmQ9+yfl0awaXEKPdvyTFm
1cQ0pn7UWWUrpOzynrAjy/fj1xeQ0C69qx44mSlxNKlGPIShaFFj17CD5F2XoAOQ
HLfl00NgLrEcsvVBwV5+b4XUi+1LJ+KwzYP7U8RwTJz9p06gNPr2+Nt5ZpjeVN7p
zsnpSqz8Marmj1paqFUpVr6C/U+u+hrSmFcA6SsUZS8EVe09QlZCq345GcDUHCrh
mtjCZXtqFdXEr5dICavk7vrQx6sug3MduIDSsEvBSjmHPj7Xtdq6AS0y65u9KqlX
CswMWp8DNawyMm6P2iu+FE873cnZ9MPEQC3NB5bZnsngKeQGEZHXcD1CxZaxM2fr
Rvaxc5/NjAIdm2H9AWIYo/QmUYFFI9MDV+D7qhEsFL5uoiH3vq9MwjPKJE+oImQr
XR7xmfUnhnWSw0d/mW2wJuDwi2dcK/P2H5LhFQlrFfHdomP0rIGrNQeFjwZ8sG0D
bzATEHggGxY65IymykGXkVIuUPL5aDmJRiGcq60gkX+6o/JfD5e3BlWY7DaL8ri2
w+rSXQZbwmHrBC9NkXAa9Ku8QkGtuU0NYzkrfGelYS0mrI9BvpFy4BWAwBH5Od68
lw6sN9YB0K8cTJWYOohWLGp5FHYsSHZmib/UjqmH1MexrPyd4qiRwa/3F/46HRYC
GV7LsLR7AmQpJvU8GzJll9T5OSwYzdHN+xIXY+cCtoWgrB7Jw1ok6h8fMXMc1psz
4nRE5ROosUEcUEB9gN29EQtXJJkwoGremSzx7SQ3EExSVgbIuq9Rh/vqiriewbBX
5p5Jsk/4cnjIQWf7if5TYsW3Oq5nC5Bvld3p61X5YIMqIdTQSB5bY2S/CbqhL+c6
j3HDXrg8Dt7yW181DcpvBfwoYFGAQoRWBvE77TP2ijpzq4j4Dm//VIZjfEUg75bI
iQHhavwVmlPOi9TW/kysJlsuhrmffuIG+x9wZMSdnBbMWHAPj6goJmwgquPQ+C8Y
eLeTgwSQYwlJICmvXUYpTktdoJwesgDLfToi8O6YS60f0xMklTaBHWIqHNHwaCck
d1cGf4PBWVFUI+fcF4QMZ4eckpgUwfZ71pLuBbLPxZAgQFdOppoXf4oKG2KOe8tk
nE8kpm/5oEg+VKdKvL6y6a0+Oj4cKdUx6OqOyzWjM4qtQ4IxTyefMr2Bt7GtLSMT
poI3U+J46djbuyZiKXy0dqno0yhwrBYFIdMfSRFIYqyien2ccVgly/1cyaB2u6MO
gbQMSGXpc+9EemPdaRDIP6toaMUz1OnkN18pzLrd+0YiigYqZNsWJcP5F9QLGM7u
QZxY98mu4cUKmqTPpD67n3gZF9/wFkpsvNlc5kfdhLYh7bkNbR7oXd9cEFSfYYpn
IEKKjv3kczK2TiVdKiKIvrxio84gNMMXjds8bbwVtw4+JNvZy6lr9rDpKhg+yUpo
GvlKEaOMgpJ+Vas23+8MsA7drdg8cd3j6ceuNZiFAm2tPBwrOm30Ru/thHtNDuCp
ZvvhhJWqoXHcKZtQG+Bc9OgQt2aMDl+lAD/7CRuZAUdfwJoBVW4ni6eYMG/LiPNj
HLzDfXGR+MtoR7acx6+94VwHlbEphT+gdLI+NaJOH2HcKKLtaEXUROE1D6Yj+1p5
7Aose2tfJldQQs0blUHaFXrXA2QQ7ZeF1gdzxXNmxPAnfGvEwStGLdcxdfA+W4n0
Qx0m08xI846f86+LDrH4Os6I4fAdoDqIWA4jd8EwRHG5vzWZh4cD/mNATjgg37UO
0YKQGppH2u0Ay1QCMipmXWJVr8HOmq4XIvnNDwELhkS8kC2dP6AyI5990tAaNDu3
MIkDFZPBSjqEAVZ2FnEDotyToDFANMR1hIfeWgbyG/VxQi/Pp55gecdjr+TAPxIl
LB4Vq+A4HBJPsgVPTpfd6V8QRFP4OXfFAd+WKs9Q6QbNRcJSfevzOWQEXIt2T2Rz
4HgBZao9GcUu6BtZZvcbGjdeRmjfaiKOh9pQGTVvHuzP2xXGedGLAT3DQgH0pNv2
E41Y06lI02ykua2pAgbBkQ6VvFUJ9D7DrYOKgqgY22wqhh5P+Qu+gAvdwnSQgBPp
gRZKZZHK2cW++jn8I8NMe9y3waikSLskn8ljvrVZLA+4fpidEeW2P08mleb3t4Qn
9K1u9muIJ8wBLVetZo9j1+FcXBtJG2FWkAigX9hrLuOSLcbEjpfikKgSgMPAMioq
sL85BiH4CdmZDfsJhCZpbG+q8wBq+v9KXCRHPUBzHElWsfoBLzo+Phn07KHJewng
i6TXKch4rqz7DLD1j1Z6Mt4R5Tx0rICZ1jyjDFMFA/qNmL3ZwtNgkB4avBAE9IIN
2kwf1IWqYPB6R8DCQ15lCsqMXu+V96xc+Jabs5pnoqoLiY62NjSc5vxvNpcV9Jbj
E2O/TLj8YdHEwohlNjQ5SNrClO1X+pZjy2f4BmBDS8zY/kJUpGl76E7n25LYI1dx
pDluO+sTw4lWi9buHHVRuND9ip/lhMZigQWV6gvSJn5pTTnVb8OOnkTdzDg8aFb2
bmMUdy00qbWo8lVXI30EzNeMIpAwPqEfNOC9LWY/5SVM0rvU2U+gnI8/7C4lAr/B
1XOpnCB+bQu+u3wOVpS57IaTQEDVobKtnGRY2vTqXkw/ncsBoRY/UhTYUbCSCpvT
y8uTkfihuj4q9xjypMJ+vJ1PfMAUHWgkOV4yWXn6JJXuwrshUwqz449y4GwqEaOP
5P9X/ChES6DI/jZfcb08DZ/zOU++r+kHMJ7nyilsAlJca1X8LF5ny/dIqpVy5oUI
Ysg9KpLwz+g+btJNV0htnWW0j92AV6f0tbB7fuh6qWldgXuCIaipWHaz93Ph7ylk
tb2kZCnvAhHq48JuhXB1BTz5htFs65Gx0mmvOyS90DtkJR3mcLxVS1RO+bErzvzy
PZzUNdMxjKzuUl6jQ7TDFdjQpflqOuG0WSXekSU2ruVmEkT8/4fXJ7o/PVVr4tmN
ZMOcWLqlYGoGDUuzX9w9O6BHF41iFZrKKiePCyoiNMc5Ufo11SOWuwGE/I2+9Jdu
qfDzxh3Z73yBJIlXV+Ngd5kvENJrkvaCrohnV0VdS/piZzI0q1bFZEVS2J67UQ+L
E+2dHpvOwpck/rkCwkdLOXaYq4LGpARQiuWN4RPuWB6YEqsy+bkvGzmpKmQywx5n
cKVCpcyZ8EF6Lzv9m+tdujQK6EqFStY2ZA4Y2UzS+xnDB3HQSnG1va1E1A0fx1rn
TX5DwYyVC1hRWh4Rywb0BSt82f4F/ohg95LXcw9VypfYBs9/vhZ1/NUEb8nznU8q
kyvnkoKggkSIKSUp87rP4Zu+AQ8UcRPYSqODp6QLTQ1oaCNhMdZQcvm4XpxUQubl
Jd8C/9QOg8MrLJIalE3JZduBZiy/qq63nMCsftX11MHg+sVooTAvbWHp9uRG7zgJ
8OEE2cYiiLniZYw5Wnpq8HsDcGOiCRPA4QsKVTRuDuxwHOjdsBZtjU4J/QP5lVU2
+c9XeTMDUuWq6XIAfjteWgJ9wPeyeyPECyokBpo10dBoXtS9h8FP4x6c7jr22gmt
QEEnBgd5M6fwiK0OSiKYoNdQhe2z/CbkGNrQ3xmx8iD8NY+7Lji+ikKPINnzHwHG
2Mel292iqX5OLN/LJ53xVZVuJz5kM3fwdbd3d7zVlxH+awKjImKYAdOrmLIBe/oE
+LgAI9z/RdjRALRb01Iw7goBm4mIkPRaSk2NH0M4qY+WpzW+FKvgK30QaZ+UFo2s
uQnDHWCa1RX8AXrwxxCHUsFnH+aCICCuhVXLsxJSXz7k7dO8P9ifQ2a+dF3l7jm+
XCljOOdZxfUlIZWGVQbEXpaXXRUesJTuu52MWGSEUsejz67FubB0fosMfB98E9FL
wBhfnKP59EQxPC772yfAvSo+IzbQsZd9j9JNazLncid6VXb4+HYq+4HWK0uz12r1
SWGOOwW+q1TVc0uD1eKizdXouoDmXnjO2ak08jAnNKEfPfKGtmgzWF3ilQSrnPn9
x36zKbAKtLJCbEW4D7IiDNW7q9VVzJuZpbURfeP1MgIt3Qs6PVIDBMJlAf/+RD/v
WvQhzpsBXvCOaNlFzWLJGIj3tsKh130lYGl/Du77GZYnLP3D2YkdeMEtaeS+cwbi
KhncLXfGGIT47E+OupNLc8PsC84rmxQ6K4/OZsZ8j/wYKxTMamhwcqDm//JQE8TZ
iBre45FqMyjgChguvJ16SI7P/Dv04yDe60w62P96ta/UPuNStB3C50oLtXZUSeXG
8+AxjzaQ1edx1eaDLE/kH4aUgrK0Udu3Js5epMdgmq3zEeDGbwp3zIm/ZNY9qW51
HdC0QKKJSBDAiiWl4MvVzq4yn9kEG/h7eIoIxPgWtKZt0NpJobyW9IKpq0EpHhB8
r9jlNcCyikhJVqApCY75KkeZiOXEaUdBzGBN4hUuOLZph2/kV4n3dbvAC7vnhbPu
KwF39FgvggDbxKVIpNRdJhvUtKp6jM5Jlktt0ivUiFmDxcvYMsjIyOai0Xbw6yMy
cr/stDNOk9N3asyVB1kHPu/EWwzTM2YClVvYXaVW1wvb2DJNjh75OGylrXWHYE+2
yHjFA20qlC+ptrV4khYoLZWWALU5byBPlKMw929/lDM19zA1ZCvM7lBp7cMesICH
9Cl2+R38EvuHGNXoASqevnXzyd81BbIEKa6TXZhiI4APD4SAgbpEgYfModu9lHnd
/LRw+5RKErUMRDErmUIV64i0tXgf/OFeNSdeTuWv0xh8ZWctUeUe3p9FO/Belc/7
dH2ECjoiLEHC9iITyCFFwznmFM1avHwHOH/DHyQMh+WOEle/ALukajO/QyKDiQ/2
AlXV8c8vQok7HPVMNSaTEnnxIExHPY8/2BJYZvWdUGqGY4CPOKZ8ijaCcU8u0HqG
EGUhFplUmQat1XNWESsQyEP7P/Cn1l0xnWpk/3PCveNZvPzZuBHem1vZU4Q2/XJc
4ImH+No44tEWZ7qob2RZDj38lXJgst054bTHCLOZ0LiOVbotVcSkcTQqS8OAaf63
mRaKKhl8ZS/RDDmiaWwLPSrldWeR01NVwI9m/H3DyPGSyxiY5YkTGZGARbID2sDO
i18ORWqbVcWl2DZXqzmPjaea5xYuD1UqMwd2QuFxUNTPAg2wYfopSrb0yD5OxUfR
tJrHhlxhBoAU+IJLeNoTnDilY8sEcelscyjwxBR/lljC1SASSZR/fUGbxnBnO8hV
Oo2Iqz4js5WqGOIjd0qPgpqR0VkRQ2vPnALERVAoQ1WqCiSd9brqxJMuX7f1LJ2w
lcMKMkA0Sf2H3wki8t1mfM9hh6sDP5NtGFRz9Tu8QFUHG40WMD+0+IOeD2gJ05hc
JGtrSg0MfSc7dZpIt1E6j6tiXw4xX2+aeu2XfRNHQGD5nXmnWtcsmDg/XUUoxMYA
QALDtj7ZcJfhwtAMJDX8W6x8pJfiOVN2NABClirxuqxlWPX69NTSKx15d/I9s0ns
yQimO0kdBA/XpDyU9i/8ECat4oMteKwpCI1x/of/pB4ia32jVzOnyN5swL2WxW5t
WxBNCTlpMUg1fCXZjkTeFUNleJVCS2xROKllyHSKnxVXKBPDbHwtFSPtn6qPU54n
GYR40ruJn2b2QVfVy7oCAqDKysNfGeKpHrQbbcDDBYOsPHPiFqTsWUszyQO+aE5W
QzN0OF+xxs789PWcOQB+mKDqWfSRcbUTuGyiNscoWLKLhxSwWYoQngeYGJbzsReP
u5NCQ+gqeVKxbmtlr3lNr6pzWZy9SHb+JlKolCxjXqPrG+OxufsS02gD+amcJZF7
y2x6UowwHsZp+QzMLaQoo1pjFcBtQioiG4cx93h4dBFzMBWjnHhmfGJ3uE32DglD
io8rzJP2ybvMbNXiO61gn5Plzg7D/NqMj5o0xoxZwlRRjxkHDYtRQqO7h51Bc5kU
HNG6r5XtQkBM7BUuQLRg0aiQaBgkhLR56QmB8mgj5plEPTPy1VX9U4ovEP5ln1+z
pT6cVaZDqWLboiX1vQiqhmb8zrDeOnrqIh8Z3DFRqKo0i2vZOZfoF0VYolBpSQkV
NkmbpmrL0/2XK+GDdL+zzq/KURuPjuVTCj91GdgpBqwF/CtBxwMHEXdB1LMbvUGX
fI4bCd6bF/sJN76Z03NKNa76P56L4L6DtPPuKVHHCTQRxbkPVn+klrrTSkq8y6bZ
34HRzR54i2x7WbSwc3vfdPy4cwdtMaAgQohmIgTPfCtvYsG75/XRVh6NqVOMt2pX
Gmgig5YyfHVUPyKkxrVT/9hAlVntvEvcuO2vQXeqscjAvYUx82wxxjbZXh1XUAC3
KwClS4+BUNB3BdrS3A8FbKTd71QYKh6k590krRtFaBOZAN1DihTH5XkNdOP9X/RH
NGk+iqaAzhSsi2OpVgWakZpAi86JtBPDOgb0R2H3nSnsyarGluECg1jpSxuzIwUj
paZmgrNOPj56+B7orZsqxFrBCazjcpV7MFdy3lKuKmwa/xA5QLngJ58Q38WbGnQr
EM44Ao6m1S/b0Jj6J3HZmgUjvaK426dXWiqTsQRHSbr9shhbFkDqG/gcqP//4Jut
2r16ZH5VPkiGUQQL0q7irY3EyPqbkn+g5gWDataInJLAgqHxdYayELOGGz452mcu
M954zjH9DI+JC+EvA8tdPUW5nntlaRXDNKlNrFTLWzW2Rv6pt54zQEAUXZB4oVzS
tankyCp4SPexwnweeP9eu5iGVCqZtA1s/c2YFdAUhRKqfq2pmF7X9xyGDndmAZA7
n1ClG4Nd6cWxSs479K3g5wsVLwemVh6pTsbg50Ww/mB7uw16hgk9Xieq1rB/aQgJ
X8keSOY3xd9tbYnOIlShm2KaP9oYzE46w5Oz/7Hwg1hyDev8lnChZjXXhtNN/rC5
+4VwDhATvIerscFUoGOv89QmtXbLBpu+MO3px536BwDKGQIG/pJ5NLt7kJaBO8ER
3tyDDm5V1jhhTjcAasAz7xqED4JuzEh31WERkpmS0vZkzA32EKrAi1tM4jYIGr71
os1U6zX7rTRYmH9ywMZznFCLzOSIgA1nYnlGLl8+HyC1wdXCz0hT0c5VUOnc7Y23
7hXa1L/d2tHSOgH2TLs3gtYOpN7qvyEpTvvmeqDSkj9oVh3CgmzUTAojtgSSO8AU
ov7wzyr1SpzvJjB7MmMuxGl7l/6lzLBOqvW7GMOpTfbI9SnF9u36aG5QfpE4uZlr
ORjvvLBMdI9IXJEeT5JVaDiY4GmH/+GSs+k2GZ2zURWJuMkZpb8NNYyonSIOa/iB
fzAFsFgem7ICJhQkA03SWlxKMoiBwXRV7nm5McnxlOzAurRuNZ91tCcvxdW/sPVf
XnDqS7oZPh6MCSA7iOcERA0F9UiAVV5yHsuBwZXYtDIJ6X5sM4V6kBqQ+ybEBsE3
zxKK++mPmW8ZT27NcIaHDmRJSz6NScLX47pi1Pymnwnlq+0HtmZuMTpm/4FZzC0S
9ROYcRqkUzCyPJpV9OvIokUepzz8Emtc00+ypy9BYnxMveYm3tJBgk11y1cU8oYy
4aFSANDi9g1w0eGQWJvxsR8gZMIqbqCGNhnd64ShT1joPpgXIxdkqcNXc5zdpjJ0
9Qc2d+hx/VOwFmLvar25VWnnOoKcSIHZUS9kBGxW8YVNVzOk2s9mwWZyvhBYoz8Y
zpVG/Au+cip9w0+GlWH1Bk8OQTWJbZmH7E0mF4SHGoDxJuSoeCZP4KccXlupIGu6
WWzoK2U1yZhKwq6se0K3NK2MXzcWaK2KeHWrItU7LRt8oHRkyCBt5iEuRSGqeFfd
NW97xBoj8muLErgoXw1nm2TaAcwxCTZfy496SX16KYJfWUJHSIypGS6Hr7/yQmwR
REEpZD7zOCHCq4ddH3kvEXgAexkDDj+mcZhPrpbI7xnddtO/xiSvMXJzvDLUb+2N
NgeErKGLAc29nF9NhqGygcLTAXnAbSHNThkBNUqZqJNoGUBZr3/sSrkeHnASs8Y2
lAdm8Y/CMkadryRI1AQjku5OJwxMvbJoK766NMBpTohBFA2kN77LrmPdVAUBtu+q
cNbAHH4Rp12R3yB+17whQ1pb01nJSQ2QkAGoECIHa5KgOnxCiMV3ZsfjjJwiRM7o
RvnUguPx/TytMltReW7P0FeZiKEq4mQ8vVsqVeVQDk0IW89bqyDjJh13rUCO38Gn
p8Mt04061pTEYmcg+kEthkecZeLelV4HxuEuNEsCFzx+1H64fXTZ7WU02Gn0MhV4
oIs0um1bvXh6PM+tjP7jj2XfecYxLJiVwWEiVVJu4s1Ebel8WnMotdLG56G2Wbr3
If+yZU2W4vDvj22DmkmSBorGbNJBnkU4wf+IGncW5UvEewLaaB6x/xgn/xDoxDso
WE83pC9hzHCKN5J/D3wP3dIMjVQ1HAAgmZjwC9iU2GFu9KZTvvOGZPE0pAQ9Tziv
qXtiW8z9I0Wy4eNYHmxjXEmJhdCCks01PVmyBzy6X5a09N2NKV1foA+mmdGiKXVo
i80Vwy4X0MCJ2CxEzqT2uRHZSnyevy3MVNF15haAA1aLp5oVIPjALbg3ewoC0LdF
KB77lU/MIO1UJ3MD3HUIL1I+7PGw5/tYlJJCp/zNvU8xpdp/depqpzceyaXCT7Iz
o/hqP0DZEs1R0kibZ9x4zLhZBL7pB+qeB6AoMd/LohY1L+YhueK25IrQyqCLi/Bc
M9at61N0R80xvUfDuHGEClNX4U6VNNP5f8/DEEOa4c2BPOSWiNm4YxbIDUtUDrGJ
ZiMZQW0ooHyzGsYED14vKh1K26Q+hgq+4Bs4j3twIJSCbVUoTYtPFLLga/ANdWDB
I62rhIcLz8kARpdYI2FwrIbYL/08Jm9wPY5+FZlfvTOFDcoDZM0zuS6jWJoPwfv0
oNHx5nwvD4hIbZeSSA3c9Qs+VaHVPzgmsyXVIO+WumIQWAzkIR5aXj+wsiXAUfqE
GsJAPhqqRw0Yf1tIpuGOCzM0lHz6dtrPT+hTZ9iF/kepmrGZjRlz181mTRbwhhFt
Ibe23ca9SEpefMKAyehDRWFumcJUREah9pe3QHGoFrp9PGTrLqLvoEMTqU03BTRF
66NNRe6A2XiyoRyRGMPDVic+hm/aRv9Sw+voW+2dMsBlp0lGUavx0yF6Y8L2+vUh
rv2ipa4HzeZV4h8yupl7Kifh44ekD91snMBG3ZP3c0MuadNvK6WB6LQSpv9t/AUQ
H8LGSiSWKZ9KWDaPP94r3mb53MhFeBxAXWR8W3tNv6ypyifVI6XpqYFSzJMLiOKa
I6CHi577KiPKtZkQlkdCkoId64y8zp7k/BtUJck++XtPa8BIOiX/n62XSn9J+d5I
UA00Ju25qHav5KFXbnbKHgl9KZMa34XgbJmkezW7LgHflJqJgqWpg0+wPZaEAfFB
bldMzt5TMleO/AO+TNOowKeEQsbR1J0pv7xkobD0mLAe6LZv47saCo2UGpZ+p0Jx
pvb+aSFeF4S+YtS5EJgfq3rFU33I83fmLPW4oE/IWyRpOqc+dDCyzukfv21vW+wM
A/UHPrJYya2uyg7dH1DrxxXrD4H1q3xmxCPg4/p0VqhQ4j+Q0yNkE2o/mBgYrWBu
sZyK0vqBMwJN4bk2jWJ16JBAPNwCPQJFB9usyg+vBzIAX/fFzUBlBZAtvl0InxdE
sbBl4X0vBMZUKRwKJeSS75UZ1ar810txXbsmFJWYv7t3xelXoQCNcTw7MsZnfEvy
EL897J+eFz1i2/6Sk7ApD/y1A+eB/ENoi3Y3pcSsoiEHGK/2YLZak+92NR7iVshb
VOu1XP/z2c2ycWAK4NfB5Dn8h5Kwey4D0eq7QBvSh1JI6KuTtpOoiPxAQuygbg0f
w73RMQ5UyjQKt9FdhnrOn7EN7kfpYaDVKAcvPZdnPZYvEL0jjGA3Rgzp1ty0m9aI
vyj+eIkv1Z+skv7s0aVHfr734EfZE2bE09svZR4lpBtr7eHVZx+/C/dbDKyyCdg4
ibbeusbyfoB6I578ysuuMTnD484mXaBxr2leJiDyPFb1aEA2Xu9V6T06MZ72dRAx
3oCvBJoC7lmKe3WJOdcRLKcERJ8fW+CNSotROn1/N8QbhspJ4KExTqFzrDCmYDV1
q0AQnsHoDEFc6GuAHPj/hDU1gyqc3sFmB3EdN/LIy7QZFa12kEwsoYAakQ0+TG+R
WoKfZTz5CeWNoVZYm6Oa11RtaQRFdfUT8/pBOa5P79GTpJL7oXDQtbMLFqN6YSDc
NeDgr+nrBCSDmF2Qfa2WhOuOSJVQyx8Z9zKP6U4qOSWlZb4IS5y/zn9uHpCFiM7+
0Nl0GVhau70Dk/YTCpJz5WHC1Djxzvj3vqdHXLMgRVXLtx1OmOp4vRNqUh7tCg/Y
TAonm9n2sCiHB99FhIA8G3P4AO8sjc9v10L9fOZ56Wx1YcjhvDFr7ZcD/Su+TN2U
syQUrLH3gH3JSLG71wysmj6lv+sLbRK+bRAbWHRXEnhek07tAYSOe6izvjye9NBD
/I/uelk7jR9bPhwX2XQ+rQeDkyIZuO/+c0aOfpInlJNKBRbnzEBS6gCk6Ua6J68X
vuZ8f9uDIq7/aqd/yWTHdghIeS0dxsaICw3WB2TsdRrOIHIH9A4Gf+2WFPg0dOGf
A3pHe3vm6pAfOy9Daa4dy4MdoL1l7wxLpQflizIUDyZVbdm6oGmkDEeo23Jq2wXK
jAkefz+cmfQ+mpAc0kcONCTiMqW/W7TPrc58YtmMPX0O22kCSXOs4pvK1Jo1iOEo
9Fu2nEBsztk5UVfV6LjJCej4fCMsX+n/mS4CI9qE2eohvdCxTiclv/LoPI/8KQd3
FN0nm8rqeF9nhOySnHLavTVI8D1RbGrOBh3KhakXxMKI5ozBXq4hrjYbVPdvUqA5
yRLHO968caePDelJUlc74Pb8KjpgWeTfwUI5Rrbq32zrFYvt67jCmMw4qB7232Mv
GEGej5YFrvcCib6olVn/243RjY7XRxllWmXZtz5VYX5wiRzZXn7XKKns6xg3HlE3
nejx4Ff+AK1w59jECTpPOXcP9NGB4f9GwjaxuyUj0q9D391RJyCzhcbc1rnWokkF
aaj4JisgPWu9MlStYEhu6XjnbYJqLSTlvecyO14nZssWCsjG4PFtTLeqONKIt6fe
AkvXj6iKnJWLnwKgyR8piJUWLQqqqeTUMPR/Hlg+/m3mdHh1M0GbNwjbHsBDQE34
ON+oHET+8joKvAc8YvNSLJ07iTwrwUg0aBNOrYBFUJ9tIaWEEe8Jlz07aQkz7hNs
MdSMPyjiarBzkCDFq7dfJn0nJZ7yXC1C1r4/sTxtmNsLa//OPoxIw+OFxfjOez2G
x8D2sXZz0Jl4TddL0LEviQGZ60yhbot/s0v9rq69KE1mgXhgervSG/ba+fAexwan
vYG2ioLNSLIyss7njYMmfMbfWZTwd/kowqpEe4ldfCxhzz+oy9/fG8pfS6YYpLJs
ptv04jzyh6h6tZOuQX4tm2X+aK+Zh+ut55/78eAW4gT0YErdevSMuZT5QRo0u3NS
IVSy8n+CEh+uPZMOYMnQKPBk7WOdjkEzejhszkROKXbGwBrN+OBrEf1rl+g/f2kZ
RTI7i69icKvyuNS7juUQxOgvH9c1itelDd1VDudKxBCasqrjBoHWfNsLpdZsZrhz
nI50/mBVyRibHBtTg4Pds8iUx2bTVJAMgML1Jjl3U+QELC8boJu2dZKjjbCcycnh
Wi25/10oOX08saOIWU2sYMBk3BzHnPuQpL+pYhEFCLLXIAGTU4Ld3UyeGiOnpXlk
q3vMjzKK3B0ZIca9K+WjtGSTwZVmbZOiV+kEnx1Nri34A5pvkReB+E712TN7sUlv
6fj7DBlPI26I1xFXAdG4THDzX2NmMjhILZ6XZ6mE1GXpKg6QNk6QXsLpl8QDBnnq
Ly5afRN8Ctj/q/mZuPgvGxSGETQ0ABf7RQpHDIBclbHsHEFzJCP2pSr1+6482oZ8
v/rwiNyQxWihrdcboGsOKFsAMIxluwQwTtp5OmkBf94Kvz+vvm1jEYpvCbsLWmyX
kz+joYvSf2p9cN+cEUVSmDNttmh6yNcAtS98YNk+cX3+fK7YDqnvJ+DHxY3x/VTc
Nj3YOmfvJ8WKqGIDHOB4BQqEx6Mo/A4fsGI0iIKi+/XC81IbOCjfwnnwgd22N8CC
NXrDD38ZFuXEYFEuIMgrSQe+wSZ3Y/NZn/Z+D8YIGZEa19CBd1VlKBcK6aUm+XPT
LVIHJB9Z9AU3ZmsesZ8Z4O6UBnV06oWqsGJn4O8/Hg9y/y9XeziFxyNtrOwYX5Bm
cMMO3/dU3UM0y9FmnRjhAl/hf2942wdRO1lj0Iq2/8bOLhoAWxEjKKq8YGcydqtP
P2cntqjJsgLibNw3j1miZkgU0+pgykNxhoC1BhwQAOXxyx5M4ET1Xh3KLjEnNpxr
ZCjwQ0hyS4o+Ud+rh8wWNOiNr34S4EJ7VcZ01s6YPy5dCI6Aq/yBCVNsUkCTA0Kf
daBXFy2RhP4SjF84IKWKkr4/PeS2G9RT9kYYHwzzhKfI4tJrRMMV11713aKPDmBb
AQ0sOtZgAVRf2m8ozAb6/lE3BZRagTl5ImvabRXrLay9IDo7t8r/sL4rqwQF8t4v
MiIN3IuNw9jIBWSeqGmsdGwcDoSO8t2wclNzS9PO0w9X+w0SPoRX3uBEP4jhHhUk
YKoCBBwfjs6eKlT3cYEbvDH91n/UAi91t//Cx1/0FLTJAZj7EVE4X9i8tYSAlVna
ZfWsc4FXV5nZlgmQZnH7xSlEEI+Rd/6nc7RHu6bAQDw6WiZez44/k69m817D71xC
midmlRI77ZuYi9O9WOpWhMNIzn53UlGz2elEPxCVQHoTkAM10F3ylcQ/PRqF8YIG
Mtpx5neK3GC0anXp4WFCjnHuOe+VHKMVQL6sQVkO55iueCjQlXbBbpIKTXLaGnfa
zI9nbg8NguBvK5KVOjpAd+IG+5ksS8FtHkXeLR7tDQ4hm+z6Nx5NpISJjpzI5u7A
y1W0A4+/Lb8Zk46dOVmd6TXzFIEdYZlHkcbd6Nse23/rvWZjHfOTkiZKXs2letfC
js4jS+PzyF2QPbXnOnok04jLFcWiFZ/c1fKsDaGK3y1vFE95cyL/lM/xih+hbiD/
VNzqGnOMJsKgUGSqJrS6+nkznmr73JI++/zKdjpMmlpKCt/1/ypB9hVmx+tMWKVN
J1eg1ishFPa8rGIKZPtPbzPKNXMEplBdpUUZv1Byw2eMoGSyAhJFMABA4JDWcfjg
p1D61bgvhmGKF+xpnWf1JvTmJXM8D3fmtENB9KCC9SwT3fgOAdZDi9D9xmTu9sEj
hg3kv+HmuYgfObL4fvMevaj3HN6VlkyR53EIfdACV00ILhLgVp7LjHR0WXTBy4d2
WB0Ox3TjzlN9wJqs682tqdaZGd6Jt/oEQ8OXGOqwwFZf8gAeLxktqMZGj4LGqNKP
0oMRiUjvnkT2zbrMUGZXhzTHnuVC0ilro1a+05UR0mYr114XxkOHpNiu78aC8Gvj
78raaFbiRpejw5dJ5ufFEoWpHh7VLNdfA+kakigA3Tf5YRrqvrFVtmVObfLUQZr6
JyJlSKzj08PV2h+B0f8YMLUWYwC0RBD0wl1xfzNekQx2fXa5Ya8JCMThIUCoFvDW
zMY7b0oB+ufzPCXSPLter+gTFDNH7RBsokTwAhM801LjoupWnSa/PTyt8YcMDhc6
Dt20+I88Jt08YCx/5SiDUXcfyDbnhxwu97Hy6crD1vp4RdDy2f4GJp9K/9ssVMmI
MtaHoWmAgtQdOG2zf+7EVinmk0hvoDZfimOnspclXVklXZ3RlzU1wru5xGzyb6R/
2JaTnmEuJ37nc65U80Y6FVTx2KtPfxaa/PwK40v9g/j7aY3D2Q4U+PMMR/PseZbs
4NZ3v/p5ItmcPdrEUdGis6LLVMJ0hM5JcAI3iXwSzcaYlDTtzUKBvZjh/t9V5Tot
raHh0pBVROu1w0cvUUoJlQSJcFzLkz2mEZ3gOyQ/ao79qvGahmBbxc2aENpFAXEf
xuqiZIvezb0WkkZLHShRB5zSLO54a1AVgZkAxMkeCtp5YFNw2jLpe4/POcblgBqT
iEf5ibayjC5fuKlEJZUfakDhLCpPHOYO2PC/OoNuHlHEEHT6QU4yneZnRT0R0Ex4
hIYG/7m5vS317g/t+g4s1DqHUOnsSLSpXAc3suvRKl412UuTk0Daqqaxita7xyHB
9/0TAixGCntXAqQy2xHg6/V1NgTWEqBFSfu/mIAAF+s5svnawZIoCvXn9+FM45jF
LSuNQOHkiAH1xzATYTo5q9Oa/J2UdYHGdQGgu76Kj9ELJpUiwZtKF8QPBxNWxKcs
Ec7cM2Zcv79ieZSCI9oIgUjeQT3JBBjUaBA7Vy3xR9PPLWZ8HtPMnH41F8udFXNt
ckhnuWl051gFx7k69MTQANf5ZqSszdkuhNgGqdphDr4fHor93nQRKpOR7RgXFNQW
0VQgfghyybLRO+loKHpsUeoEoPTzYInQnVQlx/OOYVxQH0H62wTiFXIsavaYc8eG
CMRrEELxXkehDQim/s9WfYh4WXv2DG4C9daVU5eZEeZzSbjgJnFzMJasJmnAS0Ql
wOLATg0ct3JLVABPp4VBGGfer0UMdZdOoBGEYOolMgFRMWj0Fry00Xu/2KRiVroU
68ZpNVN2qpJG66KzNtE49OZXvqwyTupCyYU4c9oRYwd/m62C+sYWij3X1r7dDDwY
dmzhJG837sUac4E5/w2D0VNoBOKYe4Yd8rUr2Q11rI8sU91aboNPh0/08KcpRQZ3
qE6KMZDcpasbZF0+HY7P/QPW007odmIk0cIaaMpDyPI40FwdOi6MaLu22+AFjPq8
ttQfdDoPWCRENUmeQVJNlWXpMSyLdarZZsOkaYua/OJ2hUKe3AUH1YxhYMRXbyyN
wAxtdLBHstehx/9PVna8VR8ClNFahQujct/X+fHXrkpWRnJAGoGvVDVz6MbmYKui
pROhn1hciOH9ct8YW0x4xxeMhEllsfiDwyk+tO7ua2Fm/6pgYOBnPP6IJ8bI/AMG
Is5kPQyJdupQsq1it/bCJs55y2YMKKn73wDR5qEvZ3pIM+/oZMCoUfxsIYwHnB31
AkHNoqunBuyXMyet800B5lNk+PBxAO46bGW7uInTn9rP/keBsD/ScNcnjvUDqhpX
AQuOKGFTb6D9LlqrqpBm6tJsTtx3tj4J4wVRIU1g9hRK++L4xtIs35k9X13ZrVrX
xVrdplMGIeMapWR4uFywY3Oj8NVKdUDwpfzvubcHdfthkpFvQVrKSvhinkPb0jnb
ies6hrgzj5Y5STRn9YafESrirQrxmXQLLm8ErBy3etRtQCilK6h0BwfIYbSWadWR
vsCK2rUNi+4ehGNPg0mi3E91fWbeCXRF/12SwR5H/G6+G3IXoBf/fJvikQ5vKj0P
Pft/NDIOOo7rdFvk5Bf0PVrXFb72KOKTupnnmUhBKLY+sfcjCTFuc3Cafzb5nTuc
MlbiVjajN+E7no3QTh5UIZAlK+LNYg4povqjNCHm2vW6IUdUfz53dtFWhz7MU5sO
HVq0DwSpWtH19zQ16BQqm/rviYGvtM+XKH6qkMaBpDBdx/ZuoyvbmxRqic6Fy7zB
Imhg+7AySDLu8ITs/8wS5avlwD8YnGRoGoaxDjaHZYdWhpnNGaeZrGK8JVIQrvzK
zk62VkB3RUkbKWdAP6jQjybrWFv7lsV15IRIO6o91JODGgCPU7yrDXy34ilJ2oDz
MOxEGpXNkdkGhuRCVTPVnWD4k3yM5GC05qt0zxWZtIvC8D3/rBrcS+BMZP0X842D
tMWZ2Ncsw62TjUV40uvt/XheEZKC5NogIEmz39aRzHmMFB7HruuzfNefGpV+8iIY
yfBLJNeXt/IFNaUcJ+u7QQZ0/GtNHflm5yTSyA0QHSeoiDktFhaFyVA8rsbnkA+p
uInPxUTEsmMv09VoZDTUKm8pMdNc6YBm95ye1oLN3RqiRdVs3tyLlA99cxGm8Ipe
sLq1z+kBNjsWsHHEPyoolnYjld3YhIfqwkQwI1YLAjG4THEnQVHpJT75M/kFxSZ6
0Am3gumy8Ybrrd+I/ALqnc9HWP/xSBFznVinzoV9tr4Y6ktVVt1ZWJen8XaIeQu+
5CyIbGKpqgPnECKmjH97pMXtmPy8AwatUjx1jy02B4eQNOTlX0TestXkEVuxln9J
Dj0ddHqpJ+wR1Z3WRz1QSmL32u4VFc7lLcq7mkpOYtIQzJBiYBZP0W7qB7LXH95K
kqfIlSt31lzMyLUXEOcUwR+q3BDJwAYkqRmUFX+dvdiv9GPuENKEjpvy/rFtPlif
jdaiGYBmXQ9mxB1iOXbM5RVNs51+SJBKz3eNK6dpDfj/yeVMCrjU1mzPh3Tr0RV8
6JAy+V9g4vhTrqclUtVZaS9PKET/VLBMnai/ClRzMraV7DfgqjbjiT+vjy9NPAo9
Sx/r1Ew1pH9t26uFDJKozAb7NnSpu5cDY7aU9kgrKEfepxmqcCDc0xfdjnrFcksz
6x543tGsfixWG2WWsjM9WOk5CWzK7slDHHc5DLMRgeteYUk7yhkz9ZV3A0yDT86j
Y+Hr8y6UPaUALrm0ddRgc/wTrCaaMo5ZWovr3In3ewmJqKzsfxTN0zqeVYsPG2Ou
+c5znum/WIZnbZT9CjmAPLbE9+a8wnyHJqIwq1TSvd/GZFxMGip44wQdd7o8CEn8
kpx9gjvdmhr5ShgG6ikO43xPfTj0rFz8/bcu5rYaP7O1thlLgqD2qpRVX9X02JYe
E5vWwG2mmCNCX/VmtVCAzXXahHRdHfV16mdlq7ffNzfx5ttLpOYnaqS9NGBAzO2A
SBRf1R2giyq8eEHnZ8gmwBOXTrLGFiy0agqZNfcQPY2zLwrxm+52p/wv8VtxiMsU
jHWQLDZCXSrfdi/rpllb6ZYT8rimtGsiaXR+NSBb2oQUC9IRYLAnuuLGlVR8Yfd5
drBMr/21ZBKIF8aMCOEYQAIPaKibdlPZIYsHl8tna95tZlFdge9ohFfX2We/smCJ
D3TZ7COwGgNAuMqpQeVBhF9cWaYWCr0WvLyYH0ccn3+95GyMF+ZErHXtVFynoNk2
JifU/dEVK9vs0DmgxweKzNIYtmI+/Pv8EBI98TrsySBYxIcMjdh3uD37lp82Hxxv
MUPeJJPliSpkCYQDdThAX15RqEPQZYUM4ExTkVgvXZCdza/mKHeAZXwiCcKKLKgx
H+SmsXOs3c2pQ658mQVXdeqGLkfnCPC+H8S/XNBgQCAHsS3cQhlwF/gdhe7Hk20R
VY2xX7cn9bEh0T9dxXmOL0uY8jIfP7U+RakANR2Ny7iAFhGPNTp0jGBezw1bxuk5
5yM66Ih4wP2v8msczYbWw84gvrjcMcHLW5QUiv0iuj33xI8/m2pckQyb9gwZRf3/
U2eYYgNk/sobKtr8gw6jYu2KWoA0OuTpdMRI1GYrfDaUtvENYg2tdWRYthrSRbku
yaj39kM1DUJiw04pnvXlsC5Owb3hCL7BpSzQx6WJ1OpEGf1VjDBrOMSsk4WjgStU
71ri3zZyX+zLiYtHKezMLZNMVEv219sn37jEmYTFzDxx6SBb5mj0+EHZoKsmQru0
UoG0rj1JPEQtBr+p6KleYXXJJWwLc9SJq+ojutMfcUvocICR1iqZnRytczIohp0W
xmyv6UmA3nqJcTB1tDAg5MeM8A/PFvysUfDUft2JOaJqq4KkNHqBTPadXYk6yfGx
d230hsXnAVa1fLAhKX7TOYzDpfDzEwTdeWE8Xq5PQ6890So+paRi55hNNlz/Hy1J
zTwKoTREOR8gNUQjdGxQsVLdOD4o30XS/ajbGHTelGyDP0Ml6sJanPizq7gWxEr5
WT+fkWOMQYb6UABpdZM6KFkO97VXKSaPYD1e6iEunXbLpRdobnC7i+hQnzhRonli
3o63E+aixzegY7HnUUYB4To5qaz6PznsrP4nknaxB5GIghQd8I3QGWrKgLQux7ya
/+fTgannnefDOVG6rmQdt4Bgg57K4dv6lqw2XholPV1NnOt6Cv0+ztfzW1tvW/OH
Ov3e0r2iGFutdmWD5DWVGDFsCW/k/bFsvAPuJ0geHswFHhA5IVDZKt7WhwcI7ZeP
RlM6/0FgLV7EjKlkM2V4Z7o4hK2aV6fH1Op9PZ612IZ/Ykqy5O6U7oaKuts8zs+J
5EAj+OVkpH++Hx2e/u4c6vpz66ck7sbbUc3MnOMD0J6Ln1JARxxrAZnUib4HijAI
cYbolnJXM3ellv8hbXrO5JGz9fr4J3pphZBiYM9vB6nfZ2g3gL40Q6GzNxlStzu+
o8Bc8tESgk3SVhv3JLjz7LONo4iPaqMXrW2xeeo/QnHUNEk0V2JTP82o6pAK3wht
ex6g2Y8Mo2ix2L/iUo+wMz3NRnl3ViaWg4MHoHwqzkuglJbb3VQJIiZZ6np72B9H
v+FYEA90jhJAkW43N1ySyGQLTOq8+ZuRnSb2CVeMMShjCvER/1epQIFFpxoEqP/K
pv461USKyDfnGKJieFF0xz1FDAeHafN6JiO0CDh8bhSKYktBLDitYCCUOa5Ul+6W
JLbOJOI+24PwvkthRnTmV5y+GbXs/gxSb2vlv0XgPU3VmNGzIjeqsq9+swD3QRov
qYNsu6n5VhPwjnAkbC82vKg7gbfXIytBuXHpFxVmrcTu2/wY+hjia2jVAjwg0zz6
uzz7/zdb43NohINJGYxmcRASXuWuX31uXSNB4fYA5ufkxCUiVt+Spelx6tII3Ftk
JLUsclDMMHsWqat16sUYaDT0jiG4ov/BbthiZDpyfzt8v9UmMIONKD5mqyOF3Dnp
UE0PfBHGSBxD7heuJqz3lOf9s0wsjidCRD5dSKC1wX7fjtncfOxSoA/uJURgZWdf
uRPmK5z0bPaZ3iZBGEavpibuEYeJ6fgfM9uxWknOIywy9zvMQDZTciWlxgE/vlYN
Iuwk47gOT+pxR/PSdhyukeIy21FcO97da0y0UgieIhUYCA1AwO1qPP2zIP+EPPah
Z/Wam5h5yaia5l51FTTlktAPeDXwex+Ti7mjYhyh5oXAOl3vgjMBx908jws+2LfW
+MR29QA2/WzUW05nPlnivqiyqz51eyZ/ATiz7EsOdeUzpbZ/ePDMFsgwarVqxb7X
gwN4B5/pwntQ+nMDHEkVEaxzTiDwjNX7orImgoPc2BYSa6/MxtCmcXHWUhKRhveE
6zvu9IjmepQp/BDt09gwCRGDWihNf1ycYji3hrYh0VJfikwvcRqHI93aaof9rrwr
+RoZpXkmCppGA69axODwSR6toC0doaoP/Yz9ZpezDS9ZFKDe7T2GFlCmwd9WUOTf
V6MQnlheZ3mglykLITRWlWtcu4lxUNje9rHQ3OcOpjlMYVAV6MsYOiigb5LyIGTg
TYdeuVRqjFHl4ZhGM85capvh76O8dAJ779Q8cCyOh4sFw22gU1W9+oQt+9D2uxf7
tfvPqfLR9NeCAXgpT4qdOV9vXqASWLMCgE515NDtEll0XryHtgBdGw6w+7LH2yHz
z7EkIas6lDJ9jlQV+ZxI5TxqQwlfvr6eZZJmzrS0EKg7qetZ0PWrThdnoA/v/M68
DmQ728//3zquFq7J/ClbG0T0I9OhyF9I/IpMtDuuRQOKyXNhkRJZcB/qqjWTPoLf
NxzpbNTPxyRdjpxMVW1BRKcOkUhgGuzlAXqJbaNz2ZQSGBaxtuOpdmTYxfg0qjhL
+otIEfbpeQ4aTz+6n4N3IaX3RWf/8ASKh5z52v5YElV1yeTHCtknF3bxCFS/sJo2
HjSGuafDSjWNEaf29X/XFccgqytlzy/ybmgt+1iPfthScUr2+1M0dmSdv/IYFMq2
TAKlQm3Hl+katQFgk28OZmfG2RNaCFGNG0G4xkZRA6KZNbrC09QhgPG9tqNIHC85
4PuJUJC++m+BrErCmGlT54Y8Pi6O6NPzxXXm3tGBZgFfL6r6FFOf/lZc+fE3msH2
nmtKGuMH+mLnWn2V8sOO2NdTOx+husxjKoCeDVxvW/cDOh5yQwyIXvgetzv4xI27
VDBH+se268+wuoo9Zj449JkyGxWvz/uUsW7jmveUrZZY4dWWDMlLN6DL+L0XsBej
/cNa/Ws0GzRf6OSxO2B32hM8dMNBVtsxHaBntjVQyKQiIw3Ff81TECC0e8tnYaOw
LdWb+Pdfjy30ps+1DevH4phJkgdzu/iuFZIZbAWTFqB2I8EDYIGaBN3atNJLVW3M
OVrtyQ/DEBTf/GpDlMGYyUoz2d5qPD5EMVyugo4S8/T81mlTUPI4r3nJjw/pOjrS
3mITCVHMBMUNVla6Ta9VDEKES96c/ulkQP6zj4wKhhA5S/5eDKyr0r3gMM9hwEqr
SaGGqP/Lpz+iND6vOQ89y5lON3g0vCvjnU5nwNwAWgDjmm2akkZhwv6Y0OCSYCVq
BuncKMcZesgoIJZgKfAQMa1yx3dtVmBqlZHBJ+Goh786pKatGia6IYOd2oGz4vtu
Ans93egyG5kD8lAe7zccexpbII3n/KFZLvjZpIDnxOV0pM5EHZbZXCxlp/2JSVri
+8aFAhBHIm4fF0tzukX4bRjEC3HoUnPDCJnwB3k1Oppd+xwND7Ys3oRDPORqmUXk
F7L0JB7ALbINHxudVep/insbyUKB56E4zzUY6RLXm3IIZpuSJS+NKgjrEEbSAI8v
yo1OjWtjN0vpj0cRQneRkRCEl31MU6ESD3pGgLxHd5NNg/4qjr1Yh3AuIENpWpHf
5sB+tcrxWIxYKUHRwhN2gbZOtXEj2SWjCHVdKyrH40OMBGMQ6Y0Jr1DWXOdA/3cv
HJJnrO2lCL7QAvyWSZRKmvXGK15Z0ACxf3NDKnN63x66EFY7zas4VqggcZN2uBoG
/tdADRxrrqXMpb5M60LzjSuc5cZS9YkeUjsd9wDHE3ZQGgGuJYjdbJgbeA25mlpb
nP8v30mljk/rG77LPy50tBd4cI5YRNUTIQNf8UQI4Gdl5P/ADQ1gEJ1GsFO3zWBc
H6vL3tWe2HOQowAO2UBjidTGMjSDA86aGRMeuvdrEyP9VCjYPpjmPIipyWJAeOwh
yTT8Z6himGzBFuqpxjckOuMGtNFvU+ycDRT9O09l/0R/uNornpZHE8se9GaM5/hu
//wc6RU5zOmYYUJKKWYLFxnoIJ/SCgFJSOsdnRIBnMFLS7NhGwpddDC2ufw8eVxv
v9h+V8DiAEGc5u3ldp+w6IWOybZTXVr7XFm3kzjNvF02MrSUVSyKBIRLOCftRCCJ
mBNperv5HazKYexrneC4ot81lDpmaT2979BAJ4HrbUMkZd3orAvoBhiYAM0ZfRx8
GhTd9b97EsqxrpgD8DVk7cB9yp4y549GYqi3sJR8asdhhXHAimd3S/eguct6ylio
VZStldcOWRbdHCsCITJmjV0s8w/q8vuD0ntZVdAWVPwXs0EZLTLGJWPhMU4L+JjF
XJ7fRUVEv4mXqkECurI00w2UXqLv7nlikOZnMV4Y1mDQQ8IpxEubskSYTCJk0Urx
q1LHI1eD3S/RNDW9On4bWQQXfxcTVtA24K61VUw3YOQJnntikRSuXKj3YYw7bYkC
y+MKEliSvT5+YhFF9P4a0r05BKaYB19z43tssGrQhYpSQgjwCdt8tBrB4I4gQjug
MadE8YPvP0SOtBDmaYXoS+OArV+nEF1U7GySQ6V6QJuoEMbqvo9BCHbkafbXUOaL
LoN/udJ6uMNaDX6njDdmNinE+ESfqw8FFwXup2g0DiZIogza3E1/kZct5F3Dlbd4
JMiie2U7JIfLrV+YOynMKdrpqBYHavsPFv34o3Y5I3W1DBRFfZRmoAEAmbtJShVc
IC1jGYIlU3ku0zqyse3qukXkTA7+0O/WRkYgHN/ch32lmPPxIPKcA9l0PYNKIC2p
NjoTywW3kT/jWOvFKAStl+ggBtGfISMTP+Bo9g3eMbGyX1y65wC1TKXf3Pvi0fyh
swGgfpuuYtfJplN3C5VTY0DxzDkrKjTnAkVspEUvj+TB7lRGqNHPvxTjjFUJxhCR
xpNt9AcsSkpzR9mmnkj8uCv9lhDHBPJCofDRk/CLWnHaLE0iN5e7nJ5BE0bl3ihm
GN3Kt58DcvKm3XDMylffdUMKzVd5ktQbN+X9wz5a+I5YxFb3slT4/CnRIRD76bXk
uB8rhKS86Gs4qMRSWlY4b/3iBaJMCm63hoF8XDoV4aCGmrMIL4FVTSMqYkvdTFf6
HKRnBJ9xyH5jUyJBRiIKDQZNmZ9/h3H8c7WJKX9IZ7ZlWcbOGq0mFKpCGm0rWxD9
7QE+d4ezG2jUQ6V9w0tpTpSAQJRrQD1SdZKIehObsRXTGOxCfIorK+Pwd/iaWsfu
WpBSY3DI/HCxYI+RlxjbuomptL7+g+8+kI5Fg31eZjPfyq7rXRk5eKV6577nymCM
KYti9bgGSbTNJ5Yyd0sCPv6WQSbpvUT1CsyceeLfV8IwnTwRhBXmWrZg/vCO2CFF
K0kTKRuFSbcMZSaqy0Mu6Iqbh/BEwPjGq+UeN/yqdPANmpvE9ngkgXIgXlXJgFiz
HGiAverepgrzGISSlFEV6b17tah5wOnSSKEDaq4xY/GMkd0wIKcLog9sk8DRiFa6
8DSU4x1eYoz6eNOD28l0ZAF++PtvaLvc6t6XUCboR3FL31aeSkxlKWwvpbzzqhoR
WwWs1z3KUzb2TdVe8B0piG4Xkm40tEuf6cIE/75KvSC2rtzyb659K1uAMFg36V2s
pR1Be1P7fPR+mPn6WdphA1hlOKhZ9lm5ci7Ag+ZSAMjUmJWjhoHKZo06xT/134Lo
f1jXAo3nMHGnWvSiVl8+8KUJ3gPw/pud9zt5uQa5YtU0wPsPc1uDGhqs7HLs6fFk
dpwW48VU8c1eN3bT3T02CH6FV2MCKqz8aLWYf99+xDA3a5OGY20exPyXAtj5bEaA
vXpm/YMLzyS3ionzZDiK/60/0izgwhNMFjB7GEbWBOxbXsqKvNyuyieOlTJSWEiS
3mhW6BoCiHNa7cueaVl7/3umYWNdtKt3QpvyBhfTaT8QcmxUfpwFydHsGTI+Ufs1
VUSma5PUivSF0fX3NMwauw0xKYbW2Y/G7DwjtqfB8UhGE4BtOGB1bCcLlBPwCrf3
XTm7Q/35d5EA0EULsE3salycyOJ5SzEXmwYIQx3jG3jY31lXBx/wB1tVpxgPhsLi
pl8BFUmdTmR6sgoIuug34M0Neto9fuzQ7raEiJi2vR7Bkrtc0tlL9we/ALFsfOAl
T3MSZPui51Te33pjT0wDqWNjnz9FTBRjaGFrkxELLvscm2380wMAzBOEeweLg5Kj
wmnf5OViUwrpn9+zFu8fnq3UIRTFiwgBlGLnujqj4NXEoefFbORpZHzw0K/IU0f6
PrWTgITNirk/1esZ6J5H/mCaYr/Rv9Z+cBrgGKTsI9CDvZKlF4zdXFOGK61xI3MX
DEBqFGATf5wbM8TBzl9POQdXudTZa1NlijVTb0/xV8bFGGqXVZtZAOfQcB1jXDCt
8xwof9GZpErOGzwOZ93rxYYETe/yOsJWg89ckvbltmYX9QkCbhn/trtbDBqJ9n4y
DiTXvKBH03JKNmCUM1ID9d0j1rYEv1rG0HlBRWyvOmhLZHd+BcbsUl5WUSI8Hsvt
A3Sw/deZH8WjHpLJSZMCN+4UgR/IZMIZPmWXO3KsoUIH6WmL2GL4fVFSxGkHnbEH
jDohdfQdFuWlkS6fpGrkXZagbMHbYmivuSbhs6K5PzY+NIAEEOt6Jn4mRSlosHX0
+19keo66S8EXCEMBUPgoCX7bMrAhAJFL0U/U53W/jv1lyLF8t5h5CCapxNqmNv4x
tqPPGtVKp4sgx64gKarJAAcKMbzWNv5zfsmhlRUuhzlAGFn7fp/5lP8XiTr3jqB6
hvLmJAjDmY0KZn4RngqJJfaDUINiqb2mjn5je8C7COooT7XYXBJJBlxf9s4nl+C4
iBbwOzn7XF8PgWVEk96102WWYzpMdEHSmKvzkJ+70JYopZDnaDK9hzdzXQLH8ibV
QmV6eqtDPyBw5p833nNelL4Vib/ScjXUuedHnM/XNoAGBrhSCt0L5dP7IbQN384d
TT01GubM8OmxoCcTFsh0IzCehhs/XJumwxErGbL5vLMVaFHifQ7az168MH4w/CEa
EqtVPOY4FDv/YkZGnX6BP5sKg8cLM7pwWxFUIX41CdciK7A9HQjdcVSxQxXlyzV7
+Pzdw3/5UZ+Bc/8TwetaqBEGWFF26rNVDA/tiU/EMPFwdTdD40Perie5CD3ErOJM
cDEVLhW3EMfFP+lg53AhZEaiOoyjzBgNwSIFpRJkLcTaOHssk417UEg8EFxIQeCX
EclkkGTLlnzGwEgjheh+cZtC3bqrqVZ3RGpEZ4xQVjU/9MJhppmEh04h77+W9Hxq
VpQAc2TIac040hjzazviE3s93NfQ6r0G6C3W45Dlqz4GXOE45JPCq2jLS9wK0tPd
92Twb05PqldxexzzOjGItw+9CRgy8wOSnVnuqzweswxU1/JEtjkn1KhfaWEAo1+h
X2xpSofVvml8IcDhsHY2sjgLGgU983TL2HKjOhZkeNhrj0qcVSmyozGAvmKyGy6m
fMt/clvQLPfROGUJwe95LPxaez0cxa+B2tGVXjxrq/g5IZaqJ6N+OyrzTsaSeVfY
HovS3Y/U6wEiDGKBFV+CLELd3+iN0kT4ozeky34gzbP0NMRQDuQnDS0wv06gVPOK
oj3oSNNYF3uH4nAIFZYh+IqMRilmlIkIpxiLWKFbVfMJs7+DWcPSsd6ZOfROez0b
wv9rBi49LkJBCQ7x8xddSlPMSAH3Osdx+XFU2Z9wMsy1OMwMrRdrPK/25vXc3YY5
ioEDPjihl3ErXhu2gleAG1etyHeR2+SK0+EgTUo/qY+D6xk2niOc8rbeXKa1yqOP
0rL+LlLQ0T/fSqmS3HDUCLK0XrzfMYlCXeloDqIV5NeNuduqBLBDtNyXZ4co2zYo
9POZpsR/YdQz+xMmCAhc1LurZT3ldkIZ+43Cq2p+5NlhHS05oYt/r1AIhtFpjwcY
nPLV52e5EjEau5G+MFnYqWfZhxCQ0J5ONd8Mk2tFqF2bkBvaJd4rhqokipLQDUQx
axueC92qwPboF9Wzmd7WzWuJWWhe9Lsz8y5g5Rk40/H780a7q9N59bk/+zkTockt
dnt2d/D4XLdI3KfxR7ECGRVdmj11vLU4JbZON8+dMqrS/Jl6A0vB5rZ8GlYaiDD5
MErmALSVTe3szpJ8lt4g9NYPKIfypLB1qjrgHs1RbznBbPIarqSpJSaU0xlwLSvk
UczYc6Sl94oipPM6JDODYYll+YBbvy+UH29/AYJMldMnLRqQmzaQyDFcWme4HCvK
yLoSTxEuim/gkkLbyP6Zck+SCYoWQVbdOIkHCtdhD3tzIpbDaQuqGA02tYRGbG3s
4j6bt86oq32fyiQGBai5SIj2fo24Dp8ZDucG5w8qrAHbdNYtaQXS3Oiw/YoSYiJT
Q9Ngnu/Imh7O4DW9IjvxEFU5JRv+D57Du0oqHDqccoE4ugP6BbdUV3ayrDYEZUOJ
SVs+0sVH961YeHguGyg6IUsG8i2gib+kZJD/2ZX/vcQF3ITCptVEwrqn4GWmqdGp
NQNnqegMvDSD4/2VlRHvAYlxzxTPgiYJgLlC9VnKCSiC7qZCThHkRthzpQHZxkzP
pwuGiuzW6oW6/jD+s2IKt9TNb1ZHTo1nogOAE1vkllWedrzt17iHQTqKmE7iJhPF
M1OuT2jvATqy0PPuYp1gl2oENeDgfR+b9yguxgc5CQ3GjM6GTuoR6HcIHyO3Hyfz
cKT5NQ1PeJW+BGhrAQZ+g/hyO1VHxUdx9GHMQgx1h1PO2LXMDvIhse04GfZywgTc
xJeH3/AaQQrqlQFkrOD98EQoscemcke3EYxkdNvMn94erk26ON2ytD/ns0dkMJFm
aTAabuA8NYhFy2ixrj1lxD6GNPtRfKf7qB7f7QTNeiF+uAAaiolHFnUjlKKtzhAS
eoTZGPKqOzlPDmY+fD8DAEn1lBF0mGchLCvLSBFmQFD0jigdvmnRwItyIwwAyazo
WE7/quNKIYlNaubBcCdbzllA294dHJJPBAMBm1mHZHto+qU3Zyg3thRrwqFv3IcI
BGmGsAK8s9HsyllDsTniHMQGnAfb1ESLwgrl78nikeJGV/IiId+VfSumimCV/1GG
Hah/CO7AKsJ+Az0Jlw1zij1szsK9AZZLe4Ilc8TuCPEtlkhREwQWvGeCIp758J58
OqxPtcuYWE4kvXJqAzpT+SGb//ul4JcScxssdcXiBliMr4uFW+yvOb4k8p+OtlfG
MVSshjwDh7SiPTwQO33k0srUIUN5Izx3Egbku/0S/bs3n/mIb/QMDJ57UJt0dv3u
znwkZ77DsgmBOv7WIYqZ5NdcwF31rlzS5bk99hEu1xQfdpfZJu1hF8aITtb7b5f9
mCmIKZqEWq8NYZJvsvUVlzK3LdGxjdPoa5DZ7QAr6XAAt0pwcWBlDN+/0iOQbxgi
JmXPfpCl74ZatDXAhY+/7VAlHPVGLMI3anul9QlIj/Nwo/ucS+FwFbeNB4c00KpS
AzHGTXs31y9WNi8WpB3VEArCjI8LoMKmnRtLWB+86bHAwG+aLLK+DKjUGyzs3l5Y
ZgvQa+VORBiyJGX+MUkmHnUBzjYYXI+iPZ/BN8mkGl6YtGI4ciOltKbA7hbaamqW
U0d2+8L6FM5U/Ac+WyihhnVqU5b2aIkKKegK1V9SgliOK/cfwd/RAUACmJN3seBl
Okd4Z7xCl0IwRGU4zQwM9oEct2znAg/HH0WOSWVPItlLg5F0+x6aUno0rRHKE0z/
lpkZxJKxjvmfvWtjLuiuXZ0M/Wg8BS72dbZkkGSDd5jkWcJOxu4sVOTx2y3vY/CM
nLx58MUtdOWrjGaVxgnS+GqunQ6ahzz78SOC+Ka8RaXHwtpjBoVYMftKsiLcBgDB
S4b0JBHpraINjOC+/8cS3BJuyb8+2vPnhjYmfBjMZIjbZh49HtvVHh3uhoQydmJS
8vsxh1FP3PdeQXXpJrHfR17azijyIrmPh8Zcr0Xvr62aS1omOxpz19a5IlYWeVB6
U0zv4hRZHEYcnzJztnEbv0X6joZqXPDODd1v9AR3vImYRBWeA/fzY77WCxnF6XHc
F0zuN5LOTEt3Y4BKryBW+UnHBIrLet3yw3gkKqItnw0tZg7BcC7o4nJb49My8uPP
eW42WnvGfJK3oVwdQQAkqIPjxK53Q2Ab+Lh0k2ICNsY6C8d8GdFdQKe/iOV1nLMx
TyVlaQVrJ00ELCEL8HooBU+jQ6yXEW5HANZNLhE7LAJr/z4lAZ93gdG2eJXkadoc
ohq21BN387h14Wn8O2mXvZtJG2PobtBlyCht2orLQ6qlbuPnQivq1+7dB4R8HKNC
Ym13h5aZepnUiSd2v9SeJObwzZwNC3ODj+m2r6KKNuWLjpqbE8msrRbJ+Lh30xwY
7HXvf04xjimmn8F91A0jPO/AEOMkxh+UfnFNwLBFw1V5KkfJdL51itYTB7+xggYk
d9f+aR0mkq1Xwxlm/tPQTt+xQZXsFLGtWZP58ow7qqQ1GfrrFfSCkxQ7/2xWkUWu
jab06mKrSpttUzwgbksvzX2kKvysR37cEVR8Pt5UwVKfcMtgAyiJFw947IOcRjJ7
WFNPhRxiCG7HW9Wl0NiqutnLwxZOY81rHHA0SdI3pAMejdes05muTcIUeznn0fHm
1bDIiU748sTq5Vnhe1VVb9eUwsIYlypf7e6bibQm1OMSjptmybZHTvzHjq+U91UF
UPr/yXLeV6FiH58ZAMawAUdC+1ykiW0A6h75g21I6ANrNPJeLIHudJoFTUloiebu
fwIljxKcn56+UYv9Dy7USiBAx7CKkxT7UOkN8s4RTLYJse3aLh0FTSsLCKyU00+N
1zpv1B7JvTnVsAYVuScnHnUa+7+hZQMFJy/MemsHjuIEAOLE7dtSjxyiNxfIpPUY
8R8an5Gh7zzzELc5DMiOZnfh1xbVoO9hrA5NJY1reyQizI6tpsFENIkCNMK8Gp3U
OU7wxnbjoV7Ipv8MrhVn02PsjaVzFzhIHltwDWmX7OMtmv2N6yEan7ohsyZAi7uP
s8SbprzFuFia6+pakD15LevaeYCEsH+NDiRE3L46+F6IuJZUivy02b8CuFICLYL6
p9cGbMx+fKiWokAc6nl1LPRESpyVb4lqnWrfxMxfWFsI6cHiPlrt3WuFhFTHC7MD
q8QXGGEgwYVo4gO9qTFGm5Yd/KmYtANopqmVIz4+lJ/wPzK/HR8QXR8bm1Adizw0
9N67A6QgkCBKnnd8OIIFEWPDeGoHizSwnf/njN92LOYAfUoyw6IZKBUUiLXvyNAF
rKpPyU6NP9G1XcYrOkcJ27uU9coZ8zYWY5dSoHc3XrSp06uGaQrIdCi8GCeP9Mbs
X7AFAxll5qaT67sAqOj1N8qm5+Xgij6gOEv37xe0ydvzHR4vJnU1ecZcQ+u+PH5I
qL1LzzUeiAjZPi+usXvPDe0DqR6jNrVI/BdgNfWeTdCfofdgMW0z3ySzANXW+lup
L7ZiKIaRKpAksCGemNeZJZrvIVKUQGZgLCWmK0M58yUysKkzYqics4KAiPO2KyL5
0DqoPurUielxCK1u6T1kakB5bMSTrfwSdg/3YnpXOcZbcm3VWXEHojLZyEOmPkbe
23v1o8Aqgy6kMRvUJVduYEiCPVbwXTA8vyKJUEuv9UIbxDKpcyNkg4v5oCtTiro7
9pib5DWyVR2g9WQ5FAnmn3xVI2Enbx4Wy/bvKn9S/zOTz2HbZIazMlLaA3AwHYQe
GWURb39QoSHJcreTd1SR4djsL5wdE05WLmyqzRPE1z7yxYLnikRcD8DYGPG3vv5C
SEOa3+x1SrdWl/MfZmdhE67x1fmZRW8CeczisyuepIlMzJYaMexeqtvtgGb+rWtK
J8WdCQjyUz22ZdMz6lWrZN0h4XZHysh2h5001umoQ3DL7zchVp6/et/8BOSGahcu
bBfA6bBPq5S7SQUrjZZpaAF8SWvnd/oVsIGGkv7azXZ8RJA9kNiIRirnzuNwp7O6
7oXdZ7u4ebsSPb2rM1AIP38Bqn57JSSq5TSpdQ5qOVzvygVS8/LKxdCqVkmlxLG3
CvBPHORmjnZc6humYDdV9L4TPuTzga79Bh6AIUzLbs2iALxqbLlnftf7SdX8ZTOz
k1fERvldDgtX9j35STMHfVi5aEVMCq/pG4vAbPMspasKY39pPybUxzMVc/eTUHTo
e2EmBmh11kpxlAZsoXjhZ4aI/91v8ILdxYwng5RIqoFNgLm7oiGpeB/qOSAoTUq+
8VTQCSlyhedFEiGQDelbrxDifuFbwSi9BAQewLIKyiRsjw1e4kEqx/BEK+aUyK8g
uB2NQpdLxZU1XZrFaUoGADPj/PWYcAM5KSnPzICSPUjSHsFmPQmqZ+pmBJme8m90
B7+bNRFphF8PTea6KNetaTsOkopb07rW9ElIVLBGdSuiPoxipN3WlnHkJAuyXtPZ
7tZ0Yx6QoybvNy7ETcsOwKVZ3s12HhMG0/brb7VR0Ime534tVP2obqaxzFzoYRes
GWkMKy+QgksBecjCKzc1p8iKlFcpXCyBVBdMfseyw0X6Tz0+f5gGy2h294NjyYOO
E/ZmlAihFxMFwyL+CulDypQUAy4zGd4uNHgAknUQEr0OuvEgvJjWQa4kofbKxt7w
NNizGeVSnONfoTkDznU5XdqZmH2ZoVzMvYSSwW4R8Ty1pX4jVnX0eG1ikydHe2gR
Ri0mUnlsMT4XHKn9SBj0dcWyKslhL/QWW9pdIfhJ+bipR4FeYOTPEF6dyvUn37qr
IhzEoxV4HFTu9wXACmPbMFqCZPtdBpPOcJzYMwmAi7vVMpsWrsO/V8VGSEBFOrTx
BIRnul37rbyMHs/qzBnyZ7X7uyWymWZvIV+OdmpOqjmBZXwXMDfBkVbKPI7VT/uY
04rZEtgTsdOXOB4sCzKozPwtUDcLQVZ16dhvAJmAEJGCqnZDXm+NofNmE9tlbuIx
1yWKerzXhybSzOlWjHpLHMHIERBls7YpV5xOa70HUdwXs5tRHMwNd57pOihBGA4C
MaNoYKlbGYhNluDfZefXf4VJfAyQLV/M1UegUovBdlnY69YDXvo3fs855jFDj3gT
/t9EMjLQxmYpV97SroxqStd4TmUaVCoxokqklJ4YV4BCsLiXwGS8YXirJobRmUxs
7L3cv+burxTY1KLfAweWZBiCcX7wYjYyn3MyKBcGQ8CjU9KOpj+IpCYsp1xqHSeG
CAwU7ZGegvkPMx6100QTrQYabjCRcWxWukAiG2ShscyDYlkloRoGrTYOwps8IV+0
8t+ETWbkAHVyNgiMNXlXpX/LlDh9IHnbsZfLMd5fzvl1rHUIL3/MezSVQAmr4FRC
U6h85nMBxDwDmGBbw22CluSxSdKLbsLPBM3BEdN1cVcA4kyH5LqY+k1pwel/UuQf
b6QABrW2MM3ZxU7cQdFNf4Wv1wQ/Dv7d+Iv7ErqfToRymgBaU+vMZlu+DIIfx5Jg
ubyaE+DCQA4MBSB/239iAe+nFvS7qxxOG4v5h+NXruW6LXkcSd/PgZ86vxkMSdua
mtfWXVTX78lyw7rFKGQnxX0BPGQac2yNmsICRO+jwkyWhui1i2sW0bge/TJ+wJ+b
+QfYHfr67ePb+b0HrSSXU/9JikoPyy62l4JNbpjxrRGw5hWJA3skqnvLBx2NzF7i
w2ajNfz71KRIv7/Zhd8zaMG+6pd/BBnNgY8ySYZpUoo3Pn5wfzmRSDHP85yoVUiQ
Ehrj6YhbYLnZK9Rye4B8D11yesIcdMJzC9oArPsPqzxk5WNsL6lwTAYio1RMzFHI
MxKGhNxAQmd1GxnKIeOxIxmJejvfjr5u0o0u10ul4aBIxQGYSDIf5+EKmDdkzXCB
vxf1OJsgDddgerCo7JEdxJDoD8QVyn2dk1XLxSZonXX6dbZ71ZjC/RGT49Qw7Rgg
Jaj2cjHTivBRgTQb+DP8Hr65gCXvnA9qRD06BnLxdT8/8PsIVmArzJFa4b/NDD6E
dI81a/nNsDvkfsO2hoF835Wo8CLLYIlqvSLSAc+KhhUTUAW+mPz5G2XSwLNrW9P8
nvtA7SvdYdKbZisrlhe1gYlhC5iqmEhoha4PgQ9ns8iS+EuZPKgoU/kBQB2rGdSQ
i/edPqKzH6nSe4qHPJTua1AwgncJzfyCH5WyD7DwP/LfrkISZ4FdVlpI+1vqrjPR
kSGRlIy5kHgMrIddaJx5paFgIUvQDH4YiN0A/oSoQVWsGEohzojHgVZ7+DQdDThZ
tFmzVush3pTSHA6TD6FN5dekpSMf2waK+nYeBnAu8yJ2NlGAGmXJFxj2uZAR0Jnf
qv37kj4RTIX1/j/cuF+JHNeGlFkBrXU1JEhdHKdDIHlVO6TBmv/KymNOEGqeFKcl
1LJRl9GGLjM6N/dBfbQA9G8146I14brsbH8FIfs74K4uXxeQCb1utcsewzZYYJWM
Ao3SaKyGrK/Xon7QU62ZlqGt9LU81YCHR6/f0/vNRt4O0VBB7277OsBhX1Zgxi2h
lZdCnMIJsHs+JZgG2iFTudhDa4I3gMvRzUTVOq56ZtlA/+ukW/gBfbqFPUnVxaeR
nzzMENNVHXc67kHHduYygaKUL0L8Tbn9qJwoEaexpmQXk48Fbi5gQoQLoMZmb0EP
NAoullrpu0lmmAL+U+5L/vek20ItfKamKH5eVuAl8r/llcn8VKO3+daCdZFrYwbb
v6nEtHMFnf7zC/0EKR95l4LvCEnMO5Pl7RHyJLwPjX6LP7X/m7BI2+mtNzkvLctv
TfoXKK8TYMsLBd7esR4gWBDbJqYHGP5wn26zxDlEiC2GKSMHRdEa/DevRYd31yCa
ntv3xdF1hdRi6LJXwwvY0apGaj/Lpje+QLyUYcm8CoTzNMo09fcI9wQ5129azjOJ
6cs4DXfcFvRpFqD/mRirmYfw9XVG0HFaHKKX12xQh8asaIWjuh8YSA4QI8CVjath
GbPt0xEE847rioYHymP2X7wq05jrqrXhieNMRFycGNxvpqWgVzEHApHl8pq+4SnD
K6jCKMxxEvqJyb+hzzAf4rlKPi8tEXHncCNaQnjk1Q5CfU2UJyj4ozUI3g1XI6WV
pn9PKBt3cgaOBHQcQOh9UFp+WNYxxpL+7VhwRBju7W5dFR24hvenGMVBdFBV+vCk
viU0EdbHrf7DogaVs8bDiIFcXVNQ9Eb/NOjT/JGcOM8/hRXS3j+4Ud7uZRFvEoMC
irVo/mNDwOvTzcGCkCAaoDtffGxE7iET9/nhW16ig8Dv0cX2/kobIWylsEizajqg
ueed3vMoG3GOBVuNn18eNqf9cK9AKnWtH1T0tMxWfaT7keg3O+tRwIWMO5Ijmkx9
s8N34zRpKtmKLKwFdrt/fUEE2fTrdoavPc+Y4qI9ud+1ANCjt5Alxd1Efzs8fdqK
LIrKk7FnPxnQytGtjiaoh5FR5J/bqoJLrxYC1U/DQFR3JpMFRErecnGEnNtMBBHy
WT35E5IZT9OlZMM3q3vM61t85oInizLmVaPjdE6/lCaCdK4ed4FCIX9bNRTBynrP
41wtFnErhZS2FlBss0CS+p+21GQNLIuS/lOP5bZgoc614RgM8d+l0zlqDJ05uUcf
nLrhlBrj/t35HalOqEIw2L+VdJBF1G6/SeVsjos16bf7R+NNPGHrOH39UtEzsefF
nHh2sLvrmW+OOuA23g97690fSEKmr0NQxtijD2/0e4FHdOrRWPNd5W/ndOkU7efb
B6bxbShJweEV6kmSWpl3t3Yukp9l4ruXTgxC/mk4SYJTW9VANNsSgOlTDzWLW/qC
9X1CLAV++ZLiyPHoGlAuxaZygC9//gVvI7y8X+2sMVvoDMsmKAaMnnePXKuCD8AH
aneSmj5gk5ynhIkOCvkM+TqekAzRyKrlVFGn05lU/gdgREAR5DkGK1MWdwErXHlE
nI/GKgWd3OTd4RyLKXQzkXUy6TORPn8veBwE5D6wHa6df5c6nQZQyML/WbRFHE6K
rAo+jVgmiy9S9zccxXg7HaPaQSJL8IvFgqdMqlCG8u2mFA5dEys+cWIkKuC/nKKd
uvov/MkTIszyMSazWKFqtZ4UwX363Tl7ntx+N9Wv/oIAPdE1++QUTGPcHVJJsIyP
mTkVvXID6IHvOAQ3FSZ+6XIgD+uk64SF9qBG7dvR6G5kDihv1Gf81GidqL0Mrvh4
uqoHmNucm98Izn0kFopjwMokc2ClW0IgI8/Oh7m5xOOKT00kQEpGW+KiMpPF1b8T
f9Y8ag0kyoAugYTaHO1BryDR6QW1mqEGVH7eMXZ0kq6p4uhVPXbBzltOfsSx/rQS
AuSZOsAiVmuaSh2zMvIcFYTRwMmQbBBkkLB6m3lEFDmikxBr1Rm6G7zfRIEVZII7
K1QAnaoHxktFnM7x0/xPl5SUSE7Fz4cWsEy4EUeYpuanWj8D4Pk55Q0jyJUEylN1
ROTD+D0gYWu5pbX83TzF/lICuAjuZVSMsULNV68dR9aDlDU1cHpnRZy+XZlo5Bij
RfFKPi+GH0cN5xiEAxO6TCcP4iWrQgvmpP/EqMXoKoBwpSW4ZE3HZjomiooPUc8L
NeYsMfPwvxw4GtCWTa7D7SzU1VIxfT8+zKPz+Bog7SO9G79awG4hXhSDbCuBLUDI
em3a6yt9Lx+zC6QL6zWdFRANfFxaLoMKMROhDen9obYxp4rhnD+Po9nX6GfzrCMO
bhKmMgD1/qyrFa+mrmPCbEurNYjUTL2K61C0DhNKkdnByHxs/MQYiCFYdt1pba0/
J0nHVxDzWHag2G/DgrB6odXQ09B1Vph8YCjkLjRtD9An/N3KUVMHvBZuXRvZT+HE
VlD7LQtdj0kJfi7M+ZV+CWfUOrryzDt6TjGjz5EPvDT+VZhLr006AlUycAHV75tY
Cbx4MF0sgLAJrIdGHY4gV3WTrnvp3lLoaKUkDYCUlgDvgPxnNSfBEV8ZlWzYWr8u
Fo4gQ+14GXV17YVtocVbS/4Yt2nzMah2YapwXx4+hhHLZWr3EKLr/jMZwu8fsxi9
vIG1iCqMRx6klLrWKFRK+D2+IDlO5gFmeVoEmG7ccegQGISObAwhdaJ6dvDs4smT
D2wnPOq8sKdIRKUT3kYECrMClcag+1VXFK85pq+Lb01LfCcHVcEnOFRWU+0QB0+F
zx8EHl3mwWyPhvIt8Qeuny/oljJJO79a3GC+l+AvYB4CorukYFF5vyf5erAxGcn5
s59jybcRye0xavFoJBvEGYaGncNZ6PhwxIh7P3RJJuCrBgX+qyRS1l3z2OSAdI7S
KqebDaiK/IWx8JQhCc+u8b8ia+BZWO6UrlbseGMriCkziM7/yy1MfSR9tpwbxt54
JzsFco27PMAGSQ9TZNK0tYGcmHJ9Yc0S2jQMrZbNoGo24ym0cwPwn7XK7k3PmEvv
GnCMaTiVNkl3qczfsf3H71xRJnnJfRWTSw871mHS0OS1KkMzhlPz08yPNt02EJ7H
8/NCsZ8BtBJfgfR8wl5JXpMM+zGSUtTN8RoRy0+HA6Dkq/BPa8qcH4/+eO98pbbX
CWFHMdx3N4wuofA2KEw13+L4YF6GlOHk+akc/C13pmH5xQLM7kJyQqhnBWC1yZtx
2h+EFRLzD+XYVBkOXeCndGYBhXbPayJ6SnSSTmXVjWshdRpF1duznkVK8VvswcZq
HFpsS4buGHe9YAlg3Q2RmBQhw+KBFdxseGwcCJYS4u3bF9cxzARGVfo3zZ5nuB1b
MB2Nrij0LD13k+s6WPC9sxdse2BJPwYZlyYbI7gesDYOMfESr6dAy+pGSz+aNxt5
1G0EaOC2LnwLP/kXgD9qvcvHl7BazaLxIaY/7TvdOlraoC31vswCf8cSXaAP2LWA
YFdZU41juq2A+kPIfDXGfPQy40Z2Q+73oSdpreGcoveQ/nWe9h4aRD4G6O5tSIGk
ZeNRplkQpjy8rE5YHuJi08lqBFmvbrdXxWT7kfi1tf3A5+tXWpSQpiIbt8vfVHgf
`pragma protect end_protected
