// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GcdWha3433JQSewGBLBZ5Eyjpld9amfkhXlLtPXrF6fsK0r63iB6nKHurRtSjNse
Y+LWKnIXD7DFxpK7BuzTFCC3TPdveRzLhPFXXmtzEoMScSVJnmnQezw9qOngXF7+
5G5UWgoSeApZAjy3SKwTIrj9labWAsE746N0hcLsH+Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18384)
N5+toMXN36VT9tdj9qozzYkNJUmauN3hRmKhpmL8WPUOTUqh8Ooob6tzCA+CTimX
F1pMbkLPAsTPg+misv1xLU5uLoElE5ASHqfCgVIB9BTVYwVpuvAOdqnHcoM2/MXS
UVtITjE0j/Sbi5M20ukB+kqbbhNIT3PdGzxpfUd8imZVhcKNFX31+p+EP0Rq8K1s
QFW+DFxw2ILdFbSk03ippRGFPrdZ6ufHuyAei2XUV9M/hCCmcgIm4DnmN8BW4iQd
QMcd8iCFZwsBYpFlC/ts8CfMw0Hn7/8WahjwrlSeKW3im43ePl+KZKVLOk+KePVH
/ThHdiNFGnjLFLaiM7mWCfHTjgVntMChfxWw1F4VHS8S7tJ0QGGcdG133B1OAfvo
t5y4Yrg/sNx/j6kx0/gbfNTsoFcl1zEXHXqHVbbOksIv6BkjFbHO5haeIbFV6u+n
gneeBTZ4LvfCq/oD9BiSd79ZElo+TRKFm6R9OqALgaww6/dzLlrFjq15NYEGd0D5
RKXHXTY94K9TDpPLvNZKR6Fr5crrTfkcc6tM7FlXIJSQvX7fg+19NNBc+GoOpi0c
CwG8Zjnch9v4280XVNTF45SZOt4nW0NbcrA1Gtvn7ZrPKst/s2cp9RPk9jS+YcuX
ayU3scmYVnWHJiKpKl3XBppVIYTTMWcV7ik2IVPNDSqPKTmH3TtXPPNQqJrJNhrs
DHlMFJzHUNz7T4ML0nsIsF9/xqwi/6fU78/8Lh4CC5xs6HFyzj6mFJRO2Oj8yg3A
BKw1bVJdtsnvlLc/wcjR3ycFZYVKoyrN1DUg5M7nSvEMlV/sJCOJaKyv/+zlSCGX
Bsf0owxH/RKKr415akGIqhYuTrBb//pwyEVX9ga7tzCNBd6Vs8RZkvSGqehWILxf
qvgVgOy3oFDPtZUnlY0ehGHq2fUNzTFPusbfu8XV3H0hEfrUXEozDcwT0Tv9uUBp
oAk8nbKKZJ01IbfIyvOgobcBMy2ppH5k5wC4oA9HnLOYTdIZk6aFGO7aWGpG5cgi
x2avM6E8Up1qTK0e4gBWiPXyYDxZR/YOjKM9Zj2MNxQHBHexA4W7mjCP5+30T5Mh
YQ3IrQEqrF346hcCUli0i6hba67Tc0psimg+vEvRTxhFljxJBPPyNfv+9urfcUtX
nWRk+j51hzVGefO7sUOO70IglAT8tsJbV5XVqdI/HSsO8dlQ1J7TczPsB/5mSVUc
Wv6Z3wIfS/x0NWcBOAoF0QvYdAdLyqdCSdOacPv9dCSstdYWndjcT2o9jJdlcRNh
/GLmX+/kkdmV2Ww47PYOaBdXx/VABM/8qiTxeRSQxKDNVCTlnsbOrDa/Jqgcm0+5
uzLkV9utRwA61uIg4SiQWCXMwt9G4gd1BE3kGkImIuUlQFY+/beYYjI6FjM8wP0X
wncPvHK5d3qeYWEVshsNjUY/p0Glx43Hz7BgpKGsst6gpz4hK+P7o8WvM9YRXpit
9Vr8iOKAcKkZJOL8YeDkLsQBr+/9dF5aJzJrY1WFkjS/pFxQ31uQcjpW812P4hCd
/uMsQJexN7jgR00D4cPMe5g/2qc+tQ4IjVLt357q4VeMcpv0nxzapPCHErhdUXqG
gFg0bFtZ6HBeGuLghFsxVgp1Of1er9x936kIRgZRysX404vKNCe2O0+xg9h8591f
4uFMcna9uIt3ZXlVDI6qNHUf+EdevKneh6n6yfeqiYC55inD95ah8ikTWO0vFNet
2A6QnvPDINfwLqG6lWNR9VTlpFk1hGdgXDp43N2nEsVF5oz8BJ5owLhh8EJXfCcE
QWjM9YzmFRocTR5I9iFIOp57UbPKHzUg6nxrc1S//oG7ySpkOgezlP8K15MTCSZl
J2s+q0ffVw9PN5b9v3r/2sm5SJRCs/+99/XI990S/pKBTAA5r1SBPQJtrflA9vZK
lw1gjvV0OeYzIw90wbK5qhYniWDaNC4+mWnOoWBT3PXISlWMkEQa3EVfNjNd18YS
qX2tpgzngK8wo8rVObKfRptj+d9MuGyxm30/BU3LdK5niM1XrHGY18jLpNOAJrOb
wQtpdyDyXhhH3T0dIo53B+BrodLenrsIDnNZC4rUNYPltDwUuYZP9L6godK8xi9Y
LaEvZcqqndpQb74yjetYmUq6IcVu02u/coPESywNzr/ZiB5KY/HrWSqcgjMmUIHj
ESJJ2XkRuoe8ZqGsaMYUNp+0NpF+p2jnV57y95wNa3YKrWnwkKoLpDs11gaTAx/L
zLywiOREycjXFIbxMDFTA4JUdtCu3EBasCELyAdwxmd2iext9eqFN/ZbmlcCEVVQ
GKBQhggEripyp2oWOdF3vCIjkFC/XA5qjcI0E7RyQyqhw8ehGjnrfzQGQd/gxQzh
aiUc1DpcBZVLaKJaPEqVTJogoYCVPR9oD5Qo2M3QTgwDlb78l6pjJAqHOcyUrOGg
AE8j32OB4Vp+vO/baULysYox/ImxCmUpM8OAsPQ87c1CTJFocWLlTUsJW3FWGt1L
R3fez4T7BIXTYxt0TGeCNhkKIk/gISnYsqSmpfJMSuBImb4doDyNFmHvI/pqGtbQ
7QqH06euW0iVorHJxHkJmIr0ysCk//6sA0t8oGw6YHYYx4AXmStoBj4UgXwl5KGK
A0TRNByrPtN54td0BuNTNkTv6X05QFPt+/COv6Cg1/p7SeyBHdCwOYHahmRxZVnv
XTNkCw7nuLaUhtCIooxlv/IOSwlv7jkM3IMJ56QH/SeusKaQCgrGIjfwGCEthbcz
wwl6XHb0FaB/zaWqEg4wANq3W+iiOESYJQhMbbDcOvwUwlW2T6YZ2Ze2SfWhUd7G
vOBAwSlEd5dkF7cXbLo8EPzWnO5XPiZG4Xezfr5xO3K438Lw+NzDoTSk2z3PoZLz
/aQrJosyv4uF7RQZgbsF0wla7r4HhdSpyvD40jlZg2Nbhth68tG7xINPotp7iELG
nTiDGtdRRcjwP4yDU3xxks8QddYuzvCVY3QLp13iiR9RYFkSfOfvS7hAYQLFXIrx
LNB+9lVZExG5+eVPDpCEwPxeERzYlG9MJsZwrIu6v3w0/XvVOOjpe1Fjw5kUunWw
JF4XNHeKuMBLmvV295FRgmUIAFNWLKGhK2s4Uht9J5fKnx4iWLAu4ndGDSZA2NMX
0EVcLsV7BsDNSJ3xJjMhAkPeVr9yvP/ykv6Y3ir48Te7eTst0G3kFuiz3XcC0gVY
Px+SIu4MZZ2fmUFkSuYvagljHj4hbxjDAsn7xT6geeI3vQS/A9AwKm+8MIisx9pb
mXM2rjpJJ/woJ24hiJAP2aaiki5VmSOXElMHyKY8jLQ1rJEM6EfvpAUM18NPQGvd
5gzqOMb9T7YZJ7GYs0DBFs3SLY65gwb8llVS4T+Bgk9VH2EFaSHSbdQfFYxswR2Y
QeY6Z0xb7Czb/PyXTC8Y9Osda8y5UAlk9zVxdQbX7l2MurkYjS3agkohDfjOHEea
oI0uV75eY1cQiAG7DTy0Nlv8WgbYVOmu6pgiCv9Qv0ffurGAO0eUb68a+238Dwoo
pdJFivTry7u8rnWlncSOvLo03p1LYKtsTgcrcdUdBGWEfgAJDlk31r4T1nOfbw21
jSo6aA4SeOXlYIvgmDmGawby3dyDkrc5ZOyHRwfakKaph03Ai0L+wFgiO9Sblg2o
uZ/R7hBafyP/qOT26xsUk2DilyGLtEgOKjkSQOR54ECr+ohpBljOIqgtSMB58lXU
RXKDbhd9d3uGzwMyztQVoY+bSnvi5+SWTVbcCDW59Hme3c8IlSnjiLWn2Bs8FgGN
FkJcS2fJ57+oLWHnx0B2RkDGj5LViv7oAS6rgBXeyvdaOXgTzpz/jSBmTVMM9CS7
LGmour9+q9Xi44BDLLQFbKZnZB2UAIP+kI+IShb5U9MDLATWmbRKfwdDCEFzeHuN
noQCrylzjrdqZl4y32XlSORZ1Ke2d204JpRSc4TKWJ4BChRwd/z0jUfyNnPvTGqb
nHUGy2pET+SuEqwRmzKv7ocRw1pJdHL6/6gee1d3vVljT7yAkhvwk8J/CMl/rMAG
sKksOtqAHnQ18r7L9bzU/WByQz50ZE4a0MVyBt/aZ0QpjOk1LrjI/fjbq1lgxZJx
RGq5ULM/aVjI8vLzyu7LjHjMCtgJnxioYuHf7SLRJgOxepFA5XMGU5ul+jGGb94O
djqIBmBb7b+/WiowqtmV8iPppS0l6AleuMNS0VmfDboSH7OhXWwDidefzp4H+mc+
UifZ6MmEHOy5C6hpnf9WpWr09fCmmI7l7nIGqoeUcrAFnihBDdwwsob+roFgRO39
Iot04+GTMByGKjLlvNLybOuCi2Ln1fzGPCw0/EHeXNf/yEZi7CrfEUPhG7buIBFZ
cZQ7vzCEPiwjOM6AlYljhpmaHol3x0sHKWzOBkonqVXNT6wpaBCNPOxU9c12HRWo
BEfsC2SfNcfu/UKQy2Zk5P2aFJ254O9zYvHP5MJC6fay53tiAQKx3ZE0N39lQgrk
GLvqZPG0QZIbkP+oKOPXyuPgXTu9jlzxxO2fWgvlas2PM8znGnd9W68M/OFLTUAm
p1net5r5RJsSUfiny4tWq3LatiTFZxzHijo4uDTWhwrQsHGaS59fHVPtp49HHo22
lBeQmp39AgNrYxcssLU5Aw4B6bdwtmDdXL5Gh+YJnfnQztoWxA+5skVeAZrfe8IG
P65PQaHOn4ic1tNkgZ6cUCbDjjkgYzA+idlan06ju7W2r2+lIAUmzASNcFJF8DYe
Ai4BuOEUT828jz8uoB4iUQ2uPHlcGARPs30Ty0ImGcHBUIH/XPsLcLykJ3dt0nPR
ukT3yF5kFHSZZkzXst/wBIqrQyvUUHEPH48Rm6sOZvClwrzWjS9m83f6JtjQMvKV
ssUOj4HLItVELJYBLxHCfaLmSujwhEhzC/Q1PK24KpZZmvya0SdFo3rzEo5yDGXB
AzHz6N+djuzwyN2C9SA8yGsPm5y6JMLpbM3VdgxOc/sisXV/XLkewoCW3SS70SGW
ZpHopOd3ckDMTGPZVNRQpOA9fWczlagY9tlseTVZVtXNr+Jf59TGc7NLel9fj1c5
Xrd38Kc+CjiSr3B7nQgoNXGQBlfkzpRuauRyuDnv2YHARs1c0tUoHYIxmVYP8g50
sFykp3GtmN4uoH1nQTrKMl6Mf1l9LQycIVowt5I6PmTv627GIDg+ZzKcmsETVEch
bULceer/aW/oz1hMWRoie8mn6rNCYWQ5RA2AQMwCp79+JbJ+27UnsGgB+aSH/tqm
bP3An9YMSnhibRfKWi7naEuEmWIrTs5YuSUD0hH6hkJBAK+o68fvnFdOpA/2tEec
dth+GCFPj6kGM75ogQM4CluissRoD9HOWUeQjvwBV1ll8U4Vj5MOfRR9fAvgKyWl
/azVjd43ailZ5f59HBDHWyviQ4H6deb8v/d5ju9QYG/VxRN9daWVZR8SCJ5ItQd+
uM3kPpnPgco/CvHuTD1gcGtIHSbUAYbXpBca2Vtw7NdTPdfO9fklDqazEZ2Clcfc
dB+erzYmTS2EWhvKh5LYd9P7a/9rdR1KH1Mj+/PIoC8WDPLP7qbyDcyHvcu5XSjU
8ywtkXC+9c3pjwAr+A4utA7bOa6MRokz+eQs/5icuo7oGCCYzLANbvFIkNwwtU13
Vm+7GvCLxvbQxirtGT3QXAKBo2xgq09HzTaeAbRwXNtm2R1lLWYUl5PghrbWbHYT
UDhDJsdVidQOo3QlYe32346EuAgT1nfoZvuoW4nhyJixeTJGMhE9IlQJ28D9vXjM
7Gjz2Ui+yWHrL8JfGVtHUZYVU4khAanDU4BWnXOBZ5Ft1JqUF5sbc/CZU0E4yhg3
uxFfxR1k8115+Ldc8NiDOASQV4CtQOW790I8wZoUJBBrDIgAAZx4t3qAmObfM+PO
p5lhzxAuM89BRrx2xMjwmTF4/tdqneHz0PIPgssdqtmFc+KPYyo6l5q7pnDdzcvU
LbejKDpuWcl4g1eq917EcEpFWFi28PQer6rODIVTPbtHFbGvwGZJwJlFtN5+HniQ
axUAL2AigwdPZ7vDcZfro/zdP9MJy4f4K2T1Gb1HPNGkjj5De7NkZ/LtlnQCvoMr
sPWeR4FnxffFu1MGXN3Bmlo5V3ymSkitjLh6d4ByYk1feoE8qEepBUO7JqkqwvK+
oTa6mngBFRX0q1cjCRgfLRBk5BbOd7P0guAi9C92Q+1vSxtiosop9KjUUpmShy2x
yDztemG3JLjW/pExk7SXd7NjaN126lHxG+ums8Xjgw0HGWmO4l3ORvUh/uUwqHyl
1tOFvSxUa+g1qYGFwFboXH9Y5oRUzyJGezPeGYj0ldu9lP3OkvqyVnWb6KgVV2TQ
Xyn6nZ4ohoP6VUuuPhYW3wfybbZXacXtyG51uNpmre/Y2oJsafAWLmgYhlDjbLt4
BYUirws2N3GSFhftdDBB+t0U+AuVfB+FRWEt5gSzjcndPwkjeh+MfPgz/SayuGvV
BneAxqImHAglPNsbe22Yc4I3MQXIQbUTzspR7VI1nM8+6LC221bAjSb3BGx1gazk
9X4ypuogfMiFdtFG6iuRimAbtXulYUwCxouf4zwKDgBFHCWv4vieBSZ7UzIwokdz
GjhvZxM8Sx/8uH2EdNIivtUKe6c2JwSAp9nkqA1hz9B6YUGF+u5vge62ckqCybuw
6MFGNd1Tm5LZvQuEnrQJmPE6MVcu8wSQeecpOFsMFSzfiX+v1yPDuXfrQDXEmRn5
PfCB23I3JRDcg07NqPR4L8nWSoNFt65pYZUkVlNFktPCBeEPFDnku17oxEEZPEIx
eD+68NBbNOY8MTDo/KWMM19T4poMMwkFyJtQ4ASYOvJnAZCZkt8yTqX98EHwD5FI
dmemjejsx1iBfnr9//H/q1KfcCRpyXYJ1lExNQeMQiSG1e+JCZGZTxraxJdsYOu3
lA7SCU2aY1hZEO1emlLvwCIKCJLFe1Qz/ROVYKHdE7VgXZ6mvwlgv1tj1Qy3gi/N
OIobVdfP1pLEsx4d+2F/8lazD4wHRf13DzD6sOa3Pv4BaI0mPWiIKI5UBtf2IrI1
O9LiGoEGAT30olNn9OfqZG1igPA0g5M1p9S6yxpB/2oDbEUfMngjb4dXXdmua6+B
5ALqlzcAqtLeIL5iSxaTGqhFxvT8fDfwecfcjuF838WcKdA73UoNwB6OU8HoUTup
3sejmV4EIdLhq+O7Eiqd+jMq7q+2WitxpflamHUB3Rip5Ck2Fr31z+1+OvJKTcn3
M+zQr8QqRdTXlJipbbLFu4iYw0hkL/oiZ+WdsSraE1cTxbX+jVZtKIr6JvHhmNJv
8TOAkocC+GrVxvrt7UgDppPKsK96lEUV1M5e05FM6sOVG5V/O4DGhI/tRXB4FyFl
hldV9gbhjldN0z9F6OqBGz1jPZtaOCPPotu1aUK56UTdj6Joo18jkY5GjyWfV442
BfLcSsl7sGL6WpRTfQ9sTMxcxNaTI6AhHxo2E9aAVuoq3s8uBFn6VU0ogojJAP3M
3hfHTUyzIotA0skSlKiYTdQQZ4HwI0vhCvVn5oQZowTroh6Y0QRuSJxhWba7xnSg
uscHGU/NW3LcdWe/fZFweaNm/1pJCP1otcaFN7AESKXFo1Qdngzt1NBqmTcOkJxf
Aab1JOSyEl06MJ/4Au2tbfS91ROX3l3yWY/fQQ8AW0dNsV76LthUPwJpLoVB93Hc
RvCqJpOqI5lLe5Woy5Dhm0b5lMLQmsW45rD14/CDLBfrFOZYVc4oSDWmRcx5lWHr
egyXTKr+rxjPQxeJZz/Vi/1xM6iJ2xlVRbKapBpKlmqt7jKIVEWTleXSF6vgJcDR
XWeay4uijRYQpcEhmOjs1byg9xF9iotVZ7loB2amKnk/fsOisRrPeyWUNTWmr2Bc
fvxPK+VbZ2ZpvpXJtAXCzBS4Uo+MlnJTg3txOtDlGuRNmw4xombXyVqjV2OLxsrU
1+IKdiUpaDlcJfIp+EJQQmYyZHE+QyIE60JuqWVbRnuuD66aphp2AtU8OwCS2dq/
ZRul4CjILBTZFQkj7MaEQCQo4JbNJ/2xkJrg1tAhnhh5K2umc/VOzuoR4kY3CB1n
K2mTq1u7BxQnHo6N3WXX6QB6Yz8YP3Ip8qHQkw/ARBM2yILvXZhcAVF3uE6Ojgv3
C0xQfJjesUJfDIOXiUDMr9sYWSY7TAX5F11QnyZ7ArbslAFqdXr5zOb4GzJHvOlv
Gj5ORroI8zXfuqf/lW/pxKDQNBn3MNRlU0nn6CquR6xYwpEQFlZkROc8n0fj4/Zt
SNiAO1Txqgyv+zbCFv0J0d+1/yWHktPQdKqa3XGrxLmAMzoaVolS6fxPqPieQQrj
tciJos9BqGulr/XF8Ncf63/cK2wZFLHO+3x7P0PgJroent0t9SIzoU55TUoGZbUc
hLbwFsWPWc6OrS9Hq5EjOigQN4ZsDVZV+nIeTcnYNYZ56Sh+VBT+z991/tu5h3yi
zPNyZUfJnBChKKTUoS3iAGl7wunh1JvN7DMGEfypsicMc3tvipWqgLYaQ10oWMX1
rFdF6suZfbkEX5o2c8xOA5N6YEvRoNrr42JyKOOYdPjjh/jI0DpNKBpWLdqdxE3l
mTvyRIEqdrtZ5hiCTaPLD1esVj3hryGbyjt6Mgw5sfhN5JijhBdE4gPK0TrE4S8F
ogaJIhOot6PAozZ6/bmlc+lclBaj37x0pcVq7XwTME7UsXZxjWnxSzz215yB4Xjl
WKWvevbukBgN8ctV/j39bQg9ipCAlojIgScUO4HOWierf3OiBMbCKAWteACr5Hki
O8usQPr5xy8SXTh7EDcC9FqNKwA2rT81Yr7vTXbgYpHZCl9JbvMCnkUted3pB6Ax
Fe/gwo9GBvE8C3oRfRbv5Cpc974aVBCzuMb5tZ4LqFQ2fD+aDeQ0ZSvapxfKvleE
wr2GDoqz2ErBkml3rVXJNnajDSfacIBc2dyaClXUKTNQrW7Dou8D7h3fBNkdVGIo
pkeA7m/vezkpWlYXcfjhg+tSXsJfTE/yCTwJshWABqXBCxg3ZMBWqKQ0PVCtIp/l
LJN02V7mhbU6+eHs05E+eHbdURuPYHH2evcFfnNk8sH4SyKraWI6VTijMdqmnJJA
VBfl9lAkQtP9hG80IndwoVwmQwXW7S8Tg7FroVCd77kU0K/GJUoxyonN179zMRpo
r7biNZlMm+XGDPeTWcqADIUCcZgNVpjd1+ppXhhEPozNhY77zkHeAAFEfShBMlNb
/MDYAYw1djBkox7DwkPdsCFwamg2EAcWEwECevx5yJ1D3XIcK40vieZzFhB+oByg
h9Cv2xeIZ/a+MUODZ+cPC/CGL4mSoBTIdKLZvQJYW8uIYCaIHyOxOyL7KVPwC1Wt
0RDTAfO3pr18y+YjmVSitg75sEn7ADXf3MyvHvYeenO7KJUQTrTvQ359XhD751ja
yrhJmweNTyogMljr/LEryK50oUNGdahMlvU1bWTAZmiSTuSEg0UKgJX2hSJwrYyb
RadLgWhZbzF4TAm57Ze8sB3B91wV85pAbxOsP4I7K1WUhzhXBNDObC972a0+YjRX
CZQB1s3f6yg8aOC5DzH81DrI0v77vxG9Tnsq5uOvcvEZymqfIbNyPOuejfQ2f5+n
2FEgqvWP3p/mv6OjM7tey2HosiT6I/ERwkTCBVrBuCFohyE+8dWIZxLBrCllvFKA
VJAo0hjy1lkZldIsLsg4EgJ8kNpRrwWPxqtJuP8Pld8GdKwXSOT9St3UyegLq4X7
Qxsf+6OUUm7jY2nC2w1Q/FCM6odQYWvbNc7msA34nRVOQXhitjszBtLizN6OB4RK
mAEFD+JeSNfR6CHujaP4JYk/xaniLYZX0MOgCQtF2zVuwc8E38AROrX20MAQ0rmo
B0WPcy96y3eX/sGRhGqJBUH5ZfoDzrUxXa4YlfFRalyJiPL+QWX/jfs002yV9YG8
tzUYaFL8iIHmqccutvthIMNgMKK1H2+S39He86CqBis+LugysD+bi7V4aUFOls3Q
dVyXJaThbyxgvHB4tG5vpth9VLU+2pUycKgBlN/SyImmOs2MePhY+ffS58Js1BII
iEAKJpJZp3yvYgAt2npTSGgEdjAeReEEN/hRbCLiv+04CAWaeRGZG7np5HNlLyof
z4cMY6XTbHfL8diZv9TqQXXIKTgcTsrzO/z42HFzHgeVnVPYrHtXMOgmi9Ikn1md
J/jPBQ3Rz+tOppWwcVc25KRaFL9X5o3scq7kJP6A6dMSO6r4sPi0viX2i7di6yME
JcNikNaq+eTht6pd399KSzzdWyXDeANK5clWhUe5mjW1UHlNJnmDBqh7GqpDLQMs
ul6bjpxgn+SjHDAHA3HQZz9gU3IHZgUFtH3bvyjT40CP58Mo+nPtIonzRxdfQ+/t
A2A9N/gs6qocR+1oAkjDxNigBbbqNOLUWiTXfMOo6NV9IjFkxrjNrPWqv1PeRQfP
JV4SmsN2VoXorHdcI+tFRmgAJMfms9jdHy99D2VbMxUJPovIw6HTIYhKyVrzXF90
06kxZkiaF8GAaFGJRl8UZoXxgJU8p99nTPQElwk+n/SViApj3grxhIfPV8DVHk8k
6nhbzFceCcacPoIFf5Dqdd2qL4qTGK2XDDQCQ+vHajOCL16HSRkwFLLiglAKkXEl
u5fRcQI4+YzBa1Hm8qgpD0UbWBH455zw909tuSuU/Ubk9MP16gwIuD5BU8K724CL
A9HqSRp/vCY4oLQqsTQ6KldYd9JpC/D/OEwnU5pVoF7MPMl6lWu2ZDKd/iz09ase
NL17eyNjCkRZjw0UiS4ZDtUk4UWCCRb/5mDkAz7YiiBVDi4EQAxjD9E9TaxiHlBh
wy5+lHVhwnxFBK4y1nsF4iOpUJgNdsNsucbaIak7ah6m6K1Oe3USEYBX9Da+Sjxr
X/X/deEj0A1aurDjLe6icSbxm+CkHeyCoUKkLbuYLKsGjLfOgMKAGMKFofXJgl53
20+CK+7JfwjMLeT7VdHM1GH3P4KZ3Ps17VvzFKKTKlo2ZxsbBTyGWWi4YhuKY66b
VusPGxPx+HDHJFXbLRwurO3ZEKCvGKowrdWZprdLZP90efqrh3wqMWg+A4N2vM5v
kZpqJGGVxqvF1nGZXBzBEINSmAeQqlBhA90GuWpPOiaInUjzEn2eEFZVaDqDPFak
3eBEiifjOAWQMNI+tGl1caEvILJF9nZpdAiX0SUVbh6ZsKnXgwkdnUds9VjAxudF
5limWd2q+PfV9ZWnqDySnAPP84tT/AsO/V5b93cPS0bL1f+kwbrTZVw431NRgZ/s
sZDRxItvyn2O6esNCaZ3lTyaC87vfHrMIQl+TxRXnZcfhqol3tIkoWj/L8W7arNQ
rkIGWO1A8xPcX6FyYYSlevqlrlpqDx2ulb8jcenlHp+WQ6H/NYfjFdXQWPFbesgk
IqsTVmE+tEwQrNMN1YL+LKhiyrEbzkDNts0P7d4/FO9Gd5uBNa9qak44gucVlHhL
Zm4uhPCMjDzMlxnaoARiB3CyCNlORUJ+FTe5yHq1qZC2AXZIBNwntw6UusCZB52c
sJ0P0qimfDiT9vljeiKowyhFjbdCqytH2iwHShzL/3/il+bN8mdHXvTd95u3HjzY
iirAXVXvW0cMntU7atD+Zy8m7js0+t5y1W7k2b8yzrM+hzuS8EOyvoA/WJIA5Wac
LDS44/2PUD3cXUjc47iAMX/o1UGaWVIi7pKmqkBx8Dv0/u0XULFMRz2iKW4MZZQk
h+iXaQ0U0ALVb742M1xa8P+KvVixU5rBPsQE1tZxRE2UbNITQRN/uobKv/j1hsWt
7dqVOaEnBaRifC+F8kCPl1T59j+gHwbcO4emrrGVcZRSC8yEP0EmScMdrsjm5Fyv
v47MJzXMSn+BFx66GJ4buCGRK1CmIKr0UBl6V/Z6DWHodxEqApS2Go6gOnqG0EyK
UPjA+pCvFjSi1TCeuIT5lBD7nik0+jbxwIPbtjabhAQYkkwf/leT5zLKqzR9Lmhh
ECsfdN+xUsmmwFWN8KUataXYNP+gWQ7fwpIYio8WsElDyId4eKh+ipZBXk3E49bI
2xukj8TI56xJqZfj0QgZzBPgHJxE7wzy8iHgdcX9eBiLg8VHNk3iDg8tmxFD3vXd
3KTKRwjC5q0Iyb/0nUJGAZnbENZCPTf4GCm/uQzF7AGcvrJwIS8VuJafeMTFq62e
DWdbS/xd5yo8aDpw8eM5dIUIoTGnPLhCzhgK24gHYCqMjVadwdIJqHp8eRqhCnf1
HTb0eup3a/HyvgZ2XWFnMu2h/wdKFrm5g70k10UMBt3BDp2InAIwKSkqBS3/KEL3
PuRWiWFJqgIIWuaPJgl7wegx0KvM7OGKo/lrYh+eX9m1GTj3LeokNduuSImPIwhW
R1eypz+RuHZGDGiRWLzCJ112AIlFeo4vsAgy5qP4YuFWhfJlWzqKudiGxRdUlXEL
9nlwE0gkOm7Ec4Wn/FkqqVL2D+Pr+aYaTzinm7dhw03GDswMjqUSRb76BZCLgA6j
Oa1v9snYP2Bz+oFe44Q8775UkbP6coPx0QxbqGybWm/eKVyhE+//qim3dP1jq7Hl
OYF+jlw6x+/Uqe8glzz7BQlGB0LMsqEnHDuRNjQwXMaIqduNMRE2kFd+VV4twuRl
vO8TWKiM2aZf3A0UgD67yg8pp8qs3TmZUFwZDHDo404Ppz9EXVcq91P2U0SmrbXC
lUzATiOJK2VDeDNztP+eIBBuuFbPeRNX2cg/66E8q73krXIqp0fniJo6bHm3B6R/
pCSua4CO6xMtRSXLmynL3KhsNfwQi30dOpeeEM6JNS2mkKHuds4jEYt4obiQXVeA
X4M0cfBdkkusH3hqgbqLxbYLf3H/ikqy9HU3fyfHJx9Gu5EQJ4H/S4gX5DD4JlwK
cESAAc49UDCrmnqNKsrm7S3iTY2nXGHwNfZgEQ4wF9gBCVIAMY8LquIEhcoiP/yS
qwWhXK+K1aWbY4Lj+sl0/Od3NLEFj/UQQqG4fmKcXmygF7aeESdHwfAIhis7SQuu
kXzVAclhExAN9FtvtEO5G07xSqPTQu9P31WsqiFziD3sj8epwrgaTsrYdw6MNUwr
WtEe4WifKS92rOZhLZd5SSkaUrDEZ9fb6tzmJ3jGwrki8yZg4NlFXyvgmOTbbIKj
hzOKTwgi8xOmn2Sl2Q8edHGraPcaMZRXty+yjf/jel4FN40fwiIC98JvwaBlkXv9
5q9YGw6Pn9ny4/k0D/YIR6jp7O/W2pIWmVtAEJ+gkIzgZBJKjQnoxRLLyrv0y9TN
Z+bmWSp7ZXwJKbW4M5Vm5HRToG0hpmAyPiNj+ph0y/+WRJ5t5We1Rph4ws0wra25
y2SzzHhb0vDTB6a7bSe6Otzygw6YNNeLjhiDxJcHPAitPGqqrKSjhOhebd0cXwR9
6wBxxqFib4E4zEM9Uq0nviIoULRXIf/Cbe/sISQUUfDngAzmUZKS7E5En/IolPL6
eNKyWFNCnNstHZ1SSoveJTBG3ttDM6Qfi1JOj+eMYojPsaVbwuq72E4UYxJ1veci
bhMhqnK1m30PVHM1DKiNptpoHtmQHkQtrMVa/WCNb3ikzs0pUDrEW0rplIlbHPlf
K8qA+CXTY40EI66M6ed2/RbHfBfjY9UGbmb3hnko8PmxuOLJpOxytQskFsB/vAwZ
tsqPj5hq64PEMfDsZqGFgE8MQYy1d5IcEZqkTwT8D+85NRXkPLM9Stxd5aBE/kxI
Jj/BIx+vta4412qhf5bSzu1XgfT1B0zbACSNmbO5DC16vKoXGr26Nwo0cZm+OFPb
sluRwDcVRIbuvmOkKfBeERkXnJ/ZvysPurBO1rXmssHqU3Z0OsOOrRkIzT44Gkps
eUvyKsaV7kSDW6yMuKvzm5gnbDIMJg6ngc4FHSSKtdwDC7xL4vRJ8OU4jz97D7wB
HgUYtkn2OZZ8DdtQ+24uPaoNt25nThQUjIx/czz3RkpuNjgt1tBd0s06TdJMfaO7
WGZKv/ixPxRID7L4mpfAWGbuj0Mjic/lhyhmqiaxPPdbTU55E7Opuyjkkq7z9Gh1
FcEY9ZI6W50QFq3K8nIC5xUwpMuOWNYCJQ9eg9MQtD6gfqXP1gyQYxLOHj9YubOw
RoDHHmH1hBt+HoVirMULbC7LbuNWnMEKwkQYKS/W4QDQlPgl1lzgqRjbBz0wddR2
alzp/mYEe1YPqVbtIIaeu+b8tqSTYDNX6vLlxfpb+DHiZ2vgZL6dacGgHW6Vx42j
hIfA/pS7GjfKDX/XcU3BKkOPmUElBwxu8HqhqMqT+0CelJJ2cTMJ64swmsa0EK7/
BLcFrO1H5ZP/4W0NHv9hN8h3zCAdBIwZHiAWTUgtwMiYQ8kHMxam/ySxx7G9pvLm
PhlW/cpgevva0UnDrIyLztREoLm+GC2Vl3MDbvOoUnHUqB9yCx7FbGS9DeQFLXVw
NU2zJ8SiYn4tnZiGfgDhvYo73UydqsqSPeJqnOezyodLZFaB274rD6Wtoqv1816P
rlMu19otka182f2zv11h4IKelNFm0IfY8AufapiLruqIMHTLwxppPxnnddes8e6d
Oz84BXbypTTDIQ1wAMe87PjnDpLmyBydYxtvKqbzKUQlXzgRnTK8/RW0KHkuTK0T
WIfmxbcf9C61qn6bbTv53TcS50nNfOwN45oX9NndYohf3EGhiLWhZB3COAcY2S6z
ipAdqplEZJUKBzA/fZ6wVSX2aNnNdjWy+ACq4GKVs5cD1NrJ+ydC0zVHNFnMYdbH
L3pLdN0ud/9FvWungCcdoGCzn1vCCKWCWT6mUtTuuVOYwo6/rIFy20dGVLy2LOFw
doVXeUfvICGxIHPM9R7mQIT52PuhyR5PdZVFKdsTQx6eJTsU6llXEu9aQrA8dkg4
dZpPLky6mo8OxIjD2/xdWQ61WdrJf/xFs9S2m3Al7DUiOnrZ7862LKTOHRysHoBK
UBJLX8dYBmATe+ESzhhSf+6+792a4wgGwDNMBKNDMt1sUySBffypC9144gx0MWLe
0tIvogV363zEVucCtdFzJAg4P8ObcUOH0sULK/dJ2GPpEjBPxf+/DlSFWxxNbj9+
+sZHkKDeYdso2+RRANMiFFdTtwSNPBWYlzceJ/BMg2zgNK9U9uL2Gi9j6D8dju34
7oE40EvpLMYJkxfqKD+RBBO7CdTtZGhp7In+Yhl/01SrfhbDTvNHkxs17HZkNFCU
ETwbJSrwYmfmIaJqAWUdl8m9ZapfbiJ8db/mBm2G+l2nh6Brwn5lvqPS+pUhY2lN
U9UybeY5n96gN+LwF2dlxAOIhN1EiJe+ogy13DfSFOqura5I6YwJ6RO/MYsK3ckr
KUSS+HdFJH2pXNp4XLUefB9AjISuiqaMVn3qMTyadTj5rCqIKfLYenNV73Qsk+Yf
iwcnADIvXeAvUnvk75sTZktRz9yHTMyLQ0yiM39wj4VbDQzxhHg2IvjY6cc98iAk
Jgj//s5yaFwiTcm8ji9rp4Ln2TJv1Z229mbTlnOkLrFFm3/0aFibSxtCyJvcsK1c
AgUOihZUHBiiOiy5W4SzJhvrRf3x+4INJ9bZk9pQrwDpjL6kPURDTReFcyZo3UDx
5vy6+MN0DZTGKx7yenapBljjZBBEU6hoJttM6ivLKjaHgaYF+4X+gIxxmGIA1id8
fOnCWMXsHmtINKqWjlxohDKSpiSMIjmxYsTnN7W1WG4cL6hnYxUcv0evkuNh8U2L
pb22v/jt0ffPdc2WEszxZEaPVJZavWNb3iSp8hAzWQgBg9K9psxp4PWcEP5fpD7H
20xD2EDB23eihx/mppVnfD+D4i8+QDaMT20OHO9uqoeYP2VcKPIPNcxJ0yJbVX01
5qQOTlR8KHYHLP2nTeE0yeUZHZCWs3G+btBhyPyOIdX5OPdD5YZnJkUEjwDNnCOG
4D1TMkWC11ln2ric7zzw2ljjZhVJazvGLLKrfoYrudTw/GPdSlZv26zxeKWO0Bom
rtDeea44cSKaO3fGrx9lAMwlgX9Bo5WFSaUI/0ypv7e/ZxGijGiNw9VEvmzBsVDp
JqGrDwoiT8NWFtFw7bQiUyViycIvDYpD9a9Ufc+zcFadh0RHP6fHnoFhpYtcgBxz
usyja69NdTWEYyg9AGkCmDnoE34pHPzttD9Wuecp9D66ouJqzIe/O4XAlBKob09x
/LlEddjHfzxpFJSTOMdCLLFBzsjNa5nFuE0yOaEGrX114DJ526oPzy/VqQQGZ8GZ
KSt3aEiNR+cBCDMovhmBDgDNHvSbWvf8H3LKMexl4RHZoWUjVHyyyBhd3ZoffWhb
9nPMDS0N7p0lfrsIKqsbpXTKzOrsLDHDeJHny8tuelg55N3KactEO2poP1quKNnW
hLfaPpCY+gE6gY2ZmLBYl4Q+SLjkoUlZQ2mRX31l17GcGEuSIMIVsRsNTq2Q+X10
m3VG9E7a4O5suywrPknhi4yrOm75CQ4ySeMHDFHeL7zaFeHF+2+rHwJG3jVftdni
2EqJqP5p37hqQM40aptgSVW4QP0UgtR+v24/90f2aN/i7fLqeAFRw1FDgMiEylt0
QU2iB4zxzHzoH/lzjdQmrp38bLFYk+hjVWTTn/5LS6OdvSU051+AfgqyrK6Hscyl
5WY2pJ38srfagTzqTh1Jofr5L52N/gQFyqMcYNtnoQK1rXDpXm6NyT6c4edqhFyK
esojFCToIuDTqB4GoIFf71Gd7DUoqD5kuCYgU8d1y1/hCKc/jvAEPLi4fLIIzVXp
qfD078aOnGXYhx7X2DbbV1/izHHcnRB1BrlXSC0xaKEXgAfWY85L2SQnT1WAcjBf
0oq/XcKzMKJrJRaWYG6eOL8qCqf1iUxVKEYNTbUIlSlhUrahFSnTt95UHyvcgMQ5
SQ15Pfop463w8vc3Aq1qAhrnJzmLXpHgLUekCNf6aej0etRlr9he7BvnIO9lIzPE
mbgsJzQqf3vDpcQaLwbZOghTPakHzNEsdAntMhc+S1bphJWYbavLdPvMQknbgp9G
aSPTVZBVievOi1uo+LcwWIGqSIH3/bhOah+WM4G5NgGDon6OC4FElbWBnsH6DfN/
Z9ctjrU2iG0g6uRfYIISDEfstm+QtpG7mq7PTfY9vhuncQtlOCpPBBOOyQXFLXjN
guneWZXzi5r690zy32ZkCEoGmcadei7xE7Aozyp2t2Jz+xES0D5XEbAC8EVu1qTu
YxYe/IIlN92e1MVETEERSdTz9AuVJ4zZ+xClyCLNQcCkQFPJ7gWNysSLJahglg/z
0+oMQtCX/PmLrhMciqmuFwE7CM6mXOB+NToKFM/+FbmPwTPvRFITqC03Q45e0STu
fKCX8L6JFVlkTo7CKO6rmzDLe2sUgzkG9FaAqeAhNOFWa/MMWymBNs394rA1y9t6
IygNrsT7/HoiHzDI3fcO8qf5Iv0YtTuMSvd2fuvdwuel0gpDzUUut+wzTlJrvLKo
SphkIBlhrh3YbUAb7DntvfmwK7DrTKa6kvvWv/zB+8q6E0YkiFArRcSs41vjJxpy
eFg60JZgzvIWl2dq/4szHrTGAJ1yJWn2JY0Myjk7kaI9Tg6J1SZsV3MV8yDHrewc
pUrhTJxq8SCgYFj/oycp/+PZh9nYrUmPzJ0dpG0voJfwj6sxlrhS287nrPucPvN1
Zq/wCKLVRYmMDkE6SWvlqqLRlTQy7r2zW/3jF2PrYcndw71ZSiDRaLmba0POSKOY
Tced2qZad4tiYwrzGlyuIrQWn4PdIMUhvpxb8ZSlRjvBtKTNwXOSEu+qoh1grN9s
kB8YastCcxi8y0nFumGAOLf0pyqDmGTdjIQJtdTmI0VqIlHQdA9lAS4nczSiISIO
EjX6kdOjWf2K9g6BSwfUXe9uxtpU3q2j1EZNq2lmkEuNfYLn7ThHoQM+ECSL5RM1
71Hr0+cFLDHc6ICUsgSbHhNToZUsbhfBy3iY1v3eNNXiRByicA8os7ZPK0OF6FFd
IlVTP66YK//SS4NOw/ugfXI8Fl4rJcEvSZDJyKp97JcrdIjZa9Xb7JYuPBtLG34c
OpbegeR62voBJaZFArNKvUBLtDHdvtYbtPBwFwQaB3I9XSyC+JgckGh4HYHHymZL
aaFLh0gf1c+nmgpgh2T5tmF7OXjWY+YdjdL/CEUHRQt9tGtPjDeLLcGcMW+vXX72
TkWcBcyWaLf/VUKZWsT68zrGMDARLSdj2aHH6p7SXK85FjxWEMF3+2I/mVaSM+s6
wVXR7govn2pPU626IrgQcSgKOcqwpO3vJxdvaJzslt+cmuM/xfEDND0RSrQkTg+E
7/V/o7w0UDM0sV3quiShfMqXD/rNu3+KDDomsjuzSDj1ZJupFBtzhxE5xAt3OhGA
b3y9sa7a6UAjjgP2fz/1rG83di5lN15u6Jvr15+tuM11YqXYJWb92iNVK70kczj5
Nx4XgMCLJPe3ZKT6Xxmh5DCb5eG9O8C+GIAQXLIFAIIXOrNd8TbbZZnsIy7cJ5Ws
HAgxjbTXTNJTNXoSBSJ0nhVyy3E9KP40+w9lWa56afw+WoWBWwIeQOvLST/QRsdn
k+ZFNkG2rZ4V46xGLNOY7WjLmjV7nfb1fPvKVmzsUCdJ/fpcyF+KifgArwcdApLj
mAoBAUwLQVzt/rf7TEB9E5sgI60YRflW0Zo19+3TZhHRpZpPbHmFpYfFtjSLt7PQ
xHypJxBaP5lxJ47dExrieYCsIDDj+WaukfK4tnNypb4lTPscwXrdLiA5MUaB1WH+
/yiXLCMqLiVkTHp0TY2n5iKcnXmAEwlaxUv+bhC0+kNYsv85/iuGPEkofy4/cJMD
2tSW8tv1t5wP32PR/7uzYyNIAcMyORTNv7XVVyAZ0/pJEunvEMhaSsdUQX8Mg8YL
mhCkmjE4qpQ+h3aefDBB3+4DXp+HTMfuBnJt2bt/OkYRVrtYfJHw98oF94cqwxuz
dV8aPNxMJqX4/UMSA7mker3EP0nNorkyjiXF9Gp/nTYK/ZKxW9gab9HYqvpaWHbh
oL3oKmrUXgqavcxdHhjfo0Z7Uh0L8zYXeVysegalsGlT7eTtEzhcPceT1OLhFvmh
AVbVwe61h9ZvXo1LGgJ6RhxMiaZrCBBZ2Wc5yTKuLTZbAzE1Eh+85ruB3BidLeRR
06g96AiUxvEU8I7f+e2DICO840LLo7cdY+vk5l03a3+SzBGRbfzv8IaYeGXjDj0n
1+bM1wiCzrtg84ek6Lm9V+yT46ESEmFZeowmqhsEX3bd0d0M/CDTKtjRD2TIYTax
Z9VTGYvks/xXkoQKK4UaxfP9A86YWgdRCx82yQmb7wfKoGBcZydSgCdFRq7sT4Lc
E3ZZliYpuPRRO/Hp3g7K95FVilTJ3W5Vo8wPgz4j25hJVZ2UjZ1mZHqPkKCem1WR
6m5x3YJDGOtWaSO/bX0x7iev8rvzFA3mMcK2ElrZVoSbzlz5Os9Xvw7JdE/K4ipU
wS+uehf8G2gtTMD9Z6T/+CN0+ek3Tbpp3WV5ddB6bEL4h42po2kfyp4lwkfwHfEh
815QopdgwiLbJrjMJjynAwbVSPq7pQz99LN1GYCko9teEfGOdnNp7Fsn1IuWDEzB
ywAcPn8HW+oLUEtA2JGS5Kht8GeU+DghazZBpnysfECaZzpjM33gl/uEkC4/ddVo
0R/sxgmY0ncf7NXVWuIcY/KZhrpaQKUHcKE+2F7+cI1bYw+PjLe6J5fU+GGDBrMS
OE50h8kVBqTdegd38xH6OLGzR8NDhNU0C2EhQrs7faqTxsPzHP2f5SUYD73L5oRz
YComhF4kfEtC7dwLVYKgAOoR27gY4OVGvqvVkg1qnVSD433zByMz3HerBqSEjJeW
jhB9VF7T3aMx/yDeUskSRMy9lV8bh9d9Vajq3AfAiJ0brWS3WSpExae1o0NtuaMU
ru+4HavMcImQoW8++OhCdZJITAMNwbgWvvp6dgcwxu+QWJE8MwYuZn5w6lxJubZt
xV57l0WStHtMND0qI7MwgOm8gDquQ3fZoS2Du6SjeEhYz82omEjLTwBBvXvzjuJY
OwN0jFiX9i+4MoPd9O7PPB83AbcF2+IeWmbxgmmpb9bw4EV6LvZIYugGAaiY0zkz
Cd4eoccYIn9c4mNvzL0gqEOJPUuKaHQeEwrXSDXYMa2zwE3LsfqlnSaEgBYTMCcm
wNuw9TwzJJkU6C9z7VEcCzJVd/V9rJACfT3K7/BDgGbgKXTv5lktjBV71uqqKC6p
GG5ywq7DvtSLu4qBfgStOmHUChJlaEAJ4lB+eC9LIZLjNf272S600Y4rRVrJ0e/v
HnhyBqk2d3o0PJwLc3Eou72SsztIT+X0MAIRswf6JNYVLRV0Pt/BIRbCng73lvnX
gmc3FClzAKJZuaAvmRNK8xf4fZQLY0gUZntN/rbvE58u0b3DDz0sybnbNvcOh2ed
iLqWyrk5wsyF7kLV+Croyf+46oUMRkqXqWcYouFZQ5BqJaLWfiJsdX/SlOYtJkbZ
bAR4VvefMwXxXZCP/Xwj4q64Zk+Vpp4ex1+91C5w1n6qrdpVJRMbKvgIVAvEEwPP
vS1KTTafSbHbgodqEwFyWKpZNxFVCSg0bB9qi0oONhsXrtyXRYNCZlZdfbF/viW1
HKUTLSYWxSyZeaEFoxIKbRHLicQ0qHEk6VyPoWAqvPEJEQ0PqEj/zHR5AwlbBR5M
WH6A19JHQ19JAgy2crnjVMIVvJSQlWEqnFaM7xq+tIG4GtWtm9X/cGKISWcD5yxF
xDKNTjo37ocqTyW7NeX4SVPHuOM5u7AtCUQLS5kn6LRLH75gyDE2lAfp1FSs3Kzn
0h72lCKnKMcgs4OPE3J2pAcsT7I41LPho18yWdL9X5rzGQ5EuAG9uypKdm3Si6NX
ydrm+9ruO6UImWAl6HeknkBcu+D3BVAGje18e1U7IHLo2lGifuzL1aZa/JDRA7Ws
HtSeId6QMl8WLgGPGickek0n/mlmhQ2IBwhMuTyl1Rf+CVRhncoJsgskV1Rd+W6n
HwuDqERa798+syn4+iNUzdEp7DCJR79nuQVjk5FH9jya8JdKtnYxDckq4tsaHjPz
QrxstORYUUNKbVrLpJ9KLAzuzXj9TFHNL6OB1ZmGziqm0sLGZPCNsmedpgn+MxDb
yO81p3Q41oXIisI6lhS9XbJwsFGenMGVce/bKa1IVbcytbVh9v5ofLkYjoH//qPN
vASjjTEuOVW39kU3ztJDBj7V7yJfd7TbEXmWids9JRB7pdPO/DHQuNdTnGko+577
5LFVaW+HY5t/SWBqsEK3BdqUlov/vmd+xTB+BwV/dRwVdhAI1gxTtT15eb24mEWs
iOAFZtRh4sxIUzDnMEacw2QlRT7XdBfxII5yoMYtPJnGH+l12bqexS6DCJWOAghp
qEeL3ycll3ijwNPkWXnn8PDYQkm3HuDWjLh5dOD7H3645WzF08yV6FXVvXJVTYg2
w7m3WCK/7IZ/4gr9SE6LNQsknjiWJPBxjwI7+1lsL71RGbuCcUVKHhWG+3J7tob7
cP7rCa6P/fsl753Cixe8dkHqIx2csKeBUd7jtwI7feDoEI4EWE6VN6Za98tmK9BB
q8d/Fmr2HqJLwBE+QmnIclP11X54BebzZoyjqWEOjijoI1G1qv8LNeA9XPJwADk4
Ns5Mkk4qsYsO9pZ8b2k6v7YAULijWY/uniX73nXOLKM7t+ftrS+hz4opvifh3fig
NxQ0qlL9NDauA8SQvVaKXMrz7kNeDxpwz4M08XPyQH5lKmY2dOMA+FJ73kc4NjlU
8A2INgC+jkqmD+EedXyn1tkH3eG7hyl8Z/1alh/TFk1q0sY84sB7lrENG4Uo6L2K
OLxm9K2ad02DGn1dgT6UblxBY5tyPuGMn+ZmpjfqI4IjSy9k92svD1KfM84HJIHk
k6+/20wYeObnUU0ibLlSBrdM35J+oWbgJnnAElrqqWyf/YatSLHCSlUAvj5sVUg3
DzzaBqio/ZWB8Hhgq0I+0mwVwjjOsYhIp3SVw13FoW3jHG5+AZ7YONFe/IfDMabN
k7QmUgDDf6udIxqiHozdy3CrJBp4CtAV9RFcQuLT1TIbPlmxZT6DDJFZaGDiYEO1
Z6y7W3Vxks7X3clp7rSh+QApcQMhBEG0Q9vYAFbFXWXXMI58l/6KLStXL2opdToS
7FvP9gDQkYM+xuwGOc0yuTCapGHlnyW2xcgGckvBCxS2rvhuRltxHmg2WDDx6mMR
kwPSwFDCS5Qa2TlclOVO2PBWGOxPxklcCVKt+563dQ3Hr3zttwQdjRWKYyGqjP68
BMc9WlFPebHErZ7RuXaH3Kdfui/eYOL/Y9E9yE3ku0OzHysUU+96QnFivPpH7gBn
w9YnIOuuIiSAZE717x7Obu3fWYZgkCmJiXsITnSIYzhuEg0Ru6hF7YMruucQ3a3N
gK8mxTFQ3jce6lsojtd1Hx4f7dwXVA4VmDQeRONNkaSFiCX8udBEw810hVU/Q6c+
4oLxC4GlYMEk80B8RRiLPEDEt4UBkoZpBULsCkIVwyJgih0ndgOLBP9HCluX6hs/
9oPfs3ZCH74BZo+3Ibp2i1H1mK386Mm7DB48cwOZFfnQl5nsOsN4GoB398or2VKp
gzemlPFCasgurLOVr7uSlvS309w+0x0Xt/NShSpkA28gXWt/EzaVloCMFQLM1kFW
SW3Efjx8W7R+9EQrTuJTAQA0flcBoyD4TkAHER8NM6bMR5ZHn/n3mvz0hnEek90M
g9j4hObbujCk62ggx6TS4bNgRf4qbfOpRtKsxp5U8gyoKWD3FHW0ynKfJm9szTMt
6tjJLglc7MppJ15UhMCXrceK4tXwjjDJasLt92Ug023ce7AMpSWIIKnkdbUFXXhk
O7fgt/pkrwEpIXVqP4C59NbHU6GmYJttFw9/jcFxnfRHrBhRtROHSSFtIvUeQT/Q
nB7fm2A3kxiAqFEi+J0F885z71aEb3qz2Du4Fnc916JzVR7rXUnhpyY9xnR6+n1L
VzQ4fCL9UkjdmhWbGzbShhJpGewDOY6+3KLc+IIRrFu3Olg5bt6cpspmgs4k5ctZ
RNpJ0Rs/P/bXEDCcFNkYaeo0cfOWi9SGUnHwpJEIBZEEn65aWKZsaIMA5mzSnDim
iCzQ5PmPqMXpeZdRdG50CDPT4Ib95MrZ5Sxid4vbMcfhwzAFy9Lec9bs+JKsxm76
sSCBY0+dRcfdc5kau5oLO3CfM9t4lv9E9sw4bMeDtIMP62CpW5yhcWNAjF1R/OYa
ge7E2UmmCmYrfJfA0hikmS2AEF4vekR9tXiGBW/d0pqmCVdHr9UmNTcq+oFYbMbE
FJ5SRhzKgHzCQ2Z1uMYVM+bsfmVc0ulD8DmbBaqeo13uObeElJEF4hrjFDrWkRps
qRcNIKA8jWBpua227qbEJT4BbXTyWnk7ESFva0n9DePuPgvSIUat2sg/bvK24vXE
q/EykUcNkC3p3Xd/yyvLF4v7Hi5MOpxVwmoIN87z3vmxsFLUtIqlIDogDMZgy0bW
4e1ERRzTEa9PtFSY9tlkTUCRVGQsPO1qxwlqjij/577f759lax1qWrnmMjpGtfjU
ZczReVbcYf0QQNYI7QWBWWG91Z1eEe3RNceiiH4J5P3GhVx0TcT8TyO+bU0wNtU1
WXEXP76OYHSpCPLa4PjqM4MouzE9mQvP4GZ9qBMtk5VbXuhrprwl0ptFt4tv3y/o
9ClJZYLqT5oJpTb7x8zggQwG0146Yn6okbrPmX3DHs3AfsU2PJrp3GvF1exirGhs
9vEzJzyCfboSdrIoq3moRj7DfkP1v+sO2lLCRAHvCl5TxUHCKcshl3esVNxrd2aT
0TtrUN22oC++wivYUhNdU9gP1Uc/abyUPPigObpGSh/CfgqgD+026Evng0MA8ux3
qzGC1v3e/4IYpwkN4iJSTYLBG4OStvq1YOLGDAUioOMPVJ0CzGK8jwmBmmixyS0w
FdBN26LSJeiZ1hPy58h9T7FDr9eETvK+7FAcsVvuKBaIwNd0NPGqYlfFjr3gKZ4X
5tp3bkAcc8QgwfRfMUh8wIr9KedHQDvYJJzdCaeROM0BT+d958ughfOJBFH0L/P4
gOMhMxe1Kap/8Gm7kKHX0TVrn/2cqaceXCpBiJ5l8ijLxXyA9ntJigBVgKTu3d6d
EfaVuBLE0UdVUNAgImAcOHgUVXK79XWOb1Z8RBJAQ7aJCQB4MY/J0+kiGjwAAQMM
HmFlaSTJcdJWzZn3f3iB2GQ3CH3zaLapn4dBVpNPk5oCW0d1BIHvNs3W93dvfDET
Fx+75oRaR/rvMIAMfbs6YmnluhPt1dLF4kewXnkzV1NoESnPMKIQREwPMB+qiGsK
8jYGq0+uw11tl9Pkceyfy0vlYED9+m1eWyI51LYa9j0KTEix81J4ldhNK7DcP3tz
r7cD+1cuGzwBfNmDqxPgQQnb5q8334Ai5Ko7bJsrqRCFKCquUgjXSZ9WPFi8Utqh
kPnOcF4dw6mEeOq9I0KbLqEq0vHne+9tpzkQAYgnDc7LgPKp5FPeG/0RY2ZTUrww
UoqU5y77bdOoAxX08KQSCzSCigiC16i48y1CypQNjsnHN5UOZ4k8eCONTP5R3OTn
`pragma protect end_protected
