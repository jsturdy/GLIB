// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AtTnGn+18ZeA4Hp/MhSgN23BgzbjJz2Y00rJ+MTow1X759y8eV+wbQnk9P99ZjRd
dYXcgIc4nAwDuhh0UjYPmANFYkIzGligyqxLGn4K/cdJHtCzvnAiEXR8RH76NrLo
aOsM8hVEH9ZPYgCgwF21e1bXiOhEyWO1QN2Beg4K9Wk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3328)
U/9JWffmpkEToCO23fgGdz74KYJe0nZnKyjMK8GUEH6drdRyWGlI9MrV0jXSVDAa
iKZaAl6Ju1StxecrpI+XW3N2geeyAi8eYP5AqMDVKUo27e9HCiQU2kQngIYfXagj
W6Cb+S27d8lac8tzdN75mRkFXUvSAODhXSA95dGYc8IInRAMWqjRimVdF/ymja8G
4bTrbpJj5TJgeD8S3GAfuAuYBWR2Dq4euOo+DxPpLV5BvJpyazxo+w3+96MqUlOs
Zm6QNIZU415Myw3YG6wbrGu5r1Dh3VtVASj8XLaZnAXs5NDpA5PXhfVuBWWzzmnL
L71wEo6lLNudCxAhhoCOAQBDaukZKY30PyKkVXTgU2LdQPGP3pV3S1QHIZeWxe2Z
cYq3MMsvjN8ltlYNmt0yyATugzRAaUEeg/RCxdsqSlNmqfma43Q9UMvCkf42yRxb
Oqe74qTmBBexCW0Ru9gOBumF91YFBShPasGuWh/g+L75ID2w2l2wofvA/Nq68SWU
zwtP+ivznirtyFBA4GoZXeb9OPKTaDk+Qc+KrMJxQq7o4babMQmvWe5Eudm2/sfc
QaBtdz5/nTsFCqYe2icNXWaFp8I1vGpCPcM+XrCkC/lnQ7BHhYOz9tmjtCPdf4dr
cdvdzvSjMEPydlQdNx6ffzBO8/XzLBjPsFNBrN8TaQpydWhawp7yVFsu6HFYFe43
0X9QPBy6YEvGgoMfGvbj120RqdoRXTnw0kv6DKcTPiiE1rjqaVPcnnZHs4UWO50V
P7S9vuoKqO/MEiCzXfrB7RMgLmxyjEKgJXsP+ai4O2rJjOCv4D+5Fn0p6uZuIrXi
U3rTpVnz2sLeeuK2I8ZEoA58CIGJZ1dwZr5Ht1SRFjyRHogrQCdRSEMWJE252NFB
SQL/p4Xuee0kQDmaYIwZg1dKmCo5f9HXKSkvPP63+dJ6m7NQfi0/Yf1+K+MkmoJw
sOAhQuUOqFZL/uyPOKwwEHiJDbiB497+RRPoBvHkZud6B6uM8DvWRkfmHZ6oDCnY
qOS76wA8pKcJWHxTcF5LB8/D1vkHBvLW+vPS8ucRRK2frb7Q1a1TZamsSCpD/xSn
byAYbl2afkgybdiPrqNjpuY7FzjYXIyc7xhsM3eWh7KSShDg9SQMSUX7NnZlLR3p
7Jc8nIFSuPhX7d/m3bQENxUbBEqB4wQtxmsBG6RK3Q4NtHlaYRGGw4eGBNG/v+2w
ysneQ7C8gi5sfN3a72m6DoGxnKLLsMzKpJ6DuDsLmrGjWcpp6Tq9owP8rU0wZ3zi
8K/R3ZozFgn2jMoqBz1gf/KdxuhtHKT5bJTe1HRQE+A8m+fNY1JRocsw+gy/8meE
CbU5pIBBlhtD8vCS0Y/u+iLRYZB6TxzBAJyL5FSAK4dL1B4kbxW6LWXGcGJCGRid
YcdYeV9+aDxzV2WSu66I5DGDrrA/8daf5oIf1c7OvJfXucB54SxMRN0HS+p1Mk7m
35qZlfyiBA1CbYm8PCor20jVrjjz9CkhMyvbSJJaGdKpVxvnlWALzQbAwV0BO6nD
gMpeYKWAKVf6P5Uh4Z7CPUVvSTQymg3UZ8mMzLOW3Z0OuDrxjqyvATvF8N5nfi/4
jo4hLldpx7/HiwgjkYmb3KfhK+WJWNdUgrZ/fM0+hQET7p4j8tSTDJ6Ft2ZWgADc
qtFUDgggci+0HiXHYaqVjVVYE4Jya2Meb0d5Y/NdRSzJZz5Ipl9632XNSLUqqiUd
N1b+1QQ57zfFT/LIkEH4XKRSLjR0cM+TZpv7aKUhheyJ2ifc28uutnzReHvKJ0Mw
nkz26hm0OPxSIEhULwhOwj1y3gHXZvP+Mlmal3FC/+vjSfBHr10sIwNwcgxQCK3C
bpWDYnKzzfcPtlIRBi66F9/1cJK3SPcPV2cEtKwuxEoBGkIVtzgZExd1VWv4MfSk
5sUWV6ukwbGiU6EVA2PGLQIrvy3xAHJmeU/1SRRnJrXO80VyuC643171y/hYtmbq
fbJqzizLRlQ1h6zU42VTDn9X2T2Wfg3uBH/FHB7y8feR9U3bULCKJdc00f1rGBF/
sxh1MNiV0LUmMcohdFS8Heo0KDox/NNRR7+KvwyZRcBZ+5XOZUW8xO91X69Ss6uu
TRRlYNfBQ1YE/VyH66Go3UP3VkyF1W9Li0pfplGK5ozzsjDCOtIk5YwPxcxufjOo
jOen5lGIgvoNiv/cH9JZ0RXECmExhkF0X+hL+jS7HrPkOcnpN75brVdGgHLoeEUQ
wXUoqF2UYpSKe/+w5EFfkOCkOUvRowplnzyrQukcWyNLEyAOldgoG0PeGSGhuyr/
ko5pk1QB1zJQmko3DO7Ca9Qysu3ny/fWviQSqEx+EoQckTdVoyA1l6vERMbgqgU0
ml2GFiSfk58cfwSygANGXgiQnFg/gCF6UHR6rSUpHgsjDeU9Pr08rUQUS6LGlpWs
FXnBi8NiR5lduLKRs8QpMAQY4Eq2cUTERROJvDNEU+Y5d/bTtlG2mfmcG0Gq4IrI
Cd1zjlMSz4U9zIrwlEWfF5HPsmVzmWUW/jysBK8ityPQUZIbPaiUBkfsutpJ5qdg
I3vQKOSX4BnRMgDVsfFJ8UBUM0q+EIGBsyGU/VsiBPE/5WtpOLehF7oESyNbBgND
sEcwoMHVpxFPwgFGXUOOvCevsbGCwqrMif/c8it1lEm/QTbosDRlL3SosujnjFCd
XzY9DNZsWb2DlpP9MeZHdZtO8EDCEl4lt9ToOgzHKoDXLdTXZA1YAkLvkboDMWmt
irpDOFacLFN9C84HrwjtIBdF74PIo9dghKLPdcphbQfDUAyxYKDDtMLnpAYRupzf
SW5YCvR6rL450dsWJXsZ3ExRu1S1+Wb4XMmtoCwJw53zwiGJMiFOdFhZyK6tr4zb
mcpmgwFbkyboEcDQQ15H5Xr72/4BVTjRbqoSYpjc2uANhloEcO5r48FFrAknXQPU
J7uXikkomih0wGhb4eJHHLWU7JQw24xMdx8hYI+xru0rLVnW8ulyTdhSBF8Mjc41
e1nQM7JVh8LOB3KfkN1Z2OuKO88qou6M9HVsN/d26syJq5yjDECdXExGI1lmxaKo
nQadSqT1joeYtyZ0Qf4p3tW39oXBHNlco8ajMCgumlhz8ZFB5wZtIG2guSrj8Y1r
n1NtRYM7qaNIfVOGL7y+EHmTxDnynwcX22gPzs0gOGMEiTUdYYVaIMPnPLEF+Bsw
8HA1aasM+pVI7URXSiM0AzKw13oKf+CPm0Urg+N89H/OeitmkDWUn5YxVugvByJz
pJcbUy3btSghVJLmRy+uik0lIQa67+TxsRpPax2arn5JRwTOydi+u+5tovsMX3mz
LeKEhP6bvHvi7feGI93D8dyuesK4lVGeGSSRBsX2WfcP4c0q6PPs53pVe2YCAPZR
eXPABhkLPbKB5gU72bnn6P5k+LExubQjRgbIQFqMyLh+SxJjDjRTQ9Trfa37hbiE
p02Lz0LJDH4q8hYFxKzIOKfUjCgXbPl+/rOPfrvvcxtwWeRZUvSByyynoYeFoc+V
tNxXlq/hXdu8sGxtIEfkOX0OqUAtJvT+2/E3gazXKSwmVTOsEqFxzFAdZvnf6GyO
NZFl7fuvxaRLzTKGxoiZe0Dm2RHb2vfl98GkG/9lAhZ4p2mPeLThDwwDPqJqWFDD
vBY/eJJWvtrtg/AlOzO/cLrBVVJM9dVRJByElduVCcsX9mkwBKXu4Ppza/3mvZLB
DIeh3u1lIbzeBtJ79tNgEwI+GzrAfdndWNDTrX7CanvGPje9h/oBs30PyjtPnRX2
e8Ljfpq76bOkdayfJhkuuoFXQOwgBTOV3fwzvo/Jbgk+EXYRk0/Fhl0zLMF7FAUT
w7t6Yya8xNvQACbz9K81zeX4BtQBvSn+4M43r5Tz3op+s4F9+ap/E0xVhVVjL8ED
FHFl7OG4tZb+iu1M6bNfVSmlAVISAA/KTjwaXE8pyH56CT+mFLbCmO6oSO4YdII1
iEqscYkZYId8mA2Y0KmnFY68bvtZf5t1Hx04G7PZ0J/vjZXjPnX88e3aGyOzFHA5
Uosddvf/OkJYBAHP/2ty1kf7bn7mz1Gdyifo4i0o9bWenxx3Woiu0scmwBHOk0Ns
fNu5vUsN5A8SyVvB+r3qKoWip1PLvHE+yWdRyIwHB/gHdPC0Rpj685W4qZTpkJdD
7Lja932+QXK/aIhT/J25vEx9lFku6cqb49UhckHHiTSB93T6uB1HKBvpFU0nKe2n
WcDfpQsOjO+4G77Q0A0EqDP6j+Bj9CuovVkAxQPDA6W2GEEuFOzLmiFtBgB4BH0D
JMvyyL/VzLOAh59PmxMoSXVI0vu3hA7isb818wJugzM/hHe0+IiYr8wi8Gaj3LkS
3AZzTuzdy+ZusvNRk51QE9E+WhSfji4bCpt7VN7gLfzwkizppFBKzwLY+vkqSsKz
IkJQgzxmLwIVeDungO3Jpw==
`pragma protect end_protected
