// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dGYlfFjz7C62oT/wXR+2dv8aS+3IL9z0XD8iZHefcR6SI+TtBK2bUxeJ9eWmCxjy
8hvbR1L7+tg455jby4Z4oIjgxUp5oHomrmcXB+Feb9cM/23MdZLt7nTnarMZMvQ8
d4NY61R7QD55zXIjz3o5wUyVR7S81IBiwCNEcyymfB0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16752)
hGC0pVEciqn5kAEmbnY9DGmuO2nNWi2o00pypWRM7yhzzzIYPhOQ5OdMAR0De1g4
XYkB6PcpoW9eie/SzuyxSu8Q4RkvVVkQpAAIRf3aBdFDZiho+7y6uR0HRkLqOH6F
RkHoLeiC0X9CGNaQmtLGWDmsnfoubg880oSuNbu33vD2axk/dc7JdLdpm8w7/0hD
1RqveIGoO9sjqF0gXo/UVMxOHxXKjt+2AnWu/xQUNjh5/9NZJ9G78ZAmWHdbL7jK
4eiTK1eEPGmxpFSsaM/wldVEvg2snCaR4eqPAvX4psfC5qBjKb2IZvJ/79qcFFzz
PBTaYpZO8Tiwpuy58Mk0MbU04kr2atciIFfWXS79bNyU5nHgejvNU67CHdKHywEK
0o5f5fvqgMf22dS1EHiVLTZuSJbKyEH27f9jNynnt4AYj6ug8fYyOpSMko1Cz6rq
Z+oJjOB9nt1Z3CyyA1Mm1KZAlwN2jmBKkxAAOWroeqPHOSWpgpqQ5ElCB/xzdt4j
1NyY1oOgokOdfHUf68qE26/trqpATvTQmRHzPz0PDnKx6fTpKsBYxEnuI4cyTUSU
7Q5ETLL31FTY9ThAGGnFYbFPNDjApAsaCckru3Dxr/RvuhwCqqZEEmVjX36GyjQF
vo14Wo2ZQO6iOaWk5mzu/ISYWVJLDYPXLJ8Zavl8imjoXdv6vP3Q5jJG9o1jnF6h
RwLy/0FZuhFMFVy2TYeDGXN6sR46I1N8fFI3DOxsj3PK9wvtCKU/LcoeMn36SZnQ
BWIkCYNY+OGnn94sFDe+zJZYIEqbdU3Ox7qaHwQtNY5S0htlJ36B4tXP8jdb3ghW
J8Dlzl8uHveZ8AsjmaI4tw2nO8uGk8Bi9M4wLZbrFaA61vHE9OdeqNa1Y3HgSJHa
HTH3ivoI5fbJOoAUIdIMmOe4WvwNAEe947ljkw/O7MXwCRR7aChGM9XTTMXguY+e
DCDX37eKVjX/BPokfKsGwADgyrCG3D3OeM0WKCQfKxnIYRPevCZOR0YgHDGe0j9A
hcp4AXOGIwHRSn32rsgt+ffBm6JduPtH+/BoKaqwZ9JPMh9tmU4F/AJ/hfYhyjcE
hdhQO11KZhSnKUIIMtGyrSLWk0pYTwJNlgauUDL7VCEFXU6awYjyfv7JvxHsBywl
zw52NVlX8PLjz+glJatYjXTbrYj08eHvlJhLu5poz4Fe6UV6UzhizT7EJzARn3DT
O/pvebtTulkU66lbA57AJc2nWk8oT2JRRQXjdBKavoXTw1Ga7qjUTmwIVmkE0Ok1
X2nlcGMzSAJnOEPNb/CDlB7L9ab7us4PhTFHvZ9FWTKoetwNJ9wfbowoMD5dffPt
OUdzJvB0bEx7umUyhAW/1UUIy0fNavFi6eJRETbw34Ybglc77vt/hdiFMX0roO+v
ElJc+Fw9EHazjdl53zge+dEcKaAzMoG7LiwFYvMhHnlA9Gf9J1yzKg1PhsjY0SgT
Ul7g51xL/LzyeBJWTXwn4tGkwc2NTSzuXjZNN7hHjWwAQhO6mbaIn41IV5YeEwce
SGOgQGtDnfiWSTSaZx4QKI+FoRnrc4ZjRMAZ9SPiqVIk5WOvH7l8YODphiiANx0r
XvUEDQkepkjZrbM3Ux5SRFcIr+Rz/VtIyfUEBaADrdwe27HaDBOvBimbGLCPWDtv
ALDhE2BdQ29i1hQD9VcT7Nr0PvshkhVf7FTtfQi/gU5WUA/z9cymNtWcQcNSiYtZ
oRs/Pmo0hLwudkveszXHlUJvL7w1CbkcDpSgWtr9I9ZmpZFN9uqS1gzosRlcWzJf
9HPxQxI+1WSFxgcuEf/3xyN1iNsjy2wDS7v3TGnv2UMDFypnNKjrPEg9q1odnntu
S4m8pQ+wZm+Qk2uq/b1LzZsH/mYNSmpM/dOxU7MYKdWLyvhH0Sgci7rF8EWarEHI
bHbTu0mDO8tWLzybP8f9jbgtCOWwum07QMCoOKbvXs9jQXq2mnzKJMadw3jn8eQT
18lc+erCQQ40KNMcRePsywrgRcyWQeHGh18u3TLDxym00S7tnPpTABaopW6boahb
UBj4sEDoj6KYNHZaKDTJtwtW5ERhXv+RzWUosJpbPEkJcv7VQk25ObbAy5cFhI/o
9MfW7hRfuWEf3qXOhYuIlNJM5iyPUxF2JlC+nIgG+xzuQIh2t7q2bbqFOuYvApBD
OuPMYiXckRwLF0ftdUN/bZBi1A0PGKrRfVINdvrWrS1GYFVQ7aPN136trOoFj3lw
I1WmTFHZdsGRI0NZUDjDUtnG+a+z6Cbm0DFP2kinKuJOJGGFaT1eJqq0+yRF6AHD
+ol2lQ4dYTj+ZCnwU6RYHvYVa7y8ThNU5D3ozRFS9zEoOQ6+74yUfF9fW60uhxQk
Gz+ArMqwE5HJ8RTKGAEI2pGmsGJN5Y9Cx5utuPSmchqaVNClfu4WwREoEuPstczo
812N2+tYQ9wBcq6oYLEffyx68CnIQVLBHwGzwI/eWd1FrB+sXKN1Y7moQ4COLCyV
+orn4b+/nIKOho561cuXKDybzHxu+s74p8QFpf2bgAF8WpKd2O8i+7RrrmVYjh6O
Ashs7p3tjt/uqNY8zGqfsO44FBtCJvOq/RKiUwcourhn0EC+Ns0e1aXEzIrLO36M
jp5k3gPiscEJByXp3YnSFpzNHw41h1tOfHIFK0nKENB2M5hZAygpHgIHknl3QdqZ
5dlF0dBsvTW3mEt939bCdVtMSRHCVxSFlNs3Wn9IoWRxIALHtmpdruxL+a23Qrai
ICAXcRZk/Nc0vKdkIb5LczfS95+D9apWbG5aRYHHsPbFScO7mgbyzIgUHaIZu1Ui
lSwtpsBhGYom4A67k2mEhMpXyzJpf7PAVCTnmu7HruzNTOxwDNKmd4aGrDtWgBzh
ZYVYzgnuav+1P7m2cmZ/ixPBi1GkBMVFSJSsvJMK2wWbho2XGG61rQ+X/K3Egtcq
YyN42pVRJ6ZTjYPYz7GhJjVfd6YaYBuAKo7RBAuRJTiJIKy6Ghh8Hfda7R/l1moj
jwfmmYGm9wqLEl5jGSrZDCpD53SqyATaf6073Me3VLrsjxRHZ4CVEVNwD3Q0lagi
DGOGlkOjMhUxbIyhYIUv0gXRCbz8CCC45JDcT5ecUzhCtw4vf4VMIhocHppBPHp/
ESMsCrSgj/ETfEJcqWJlW29tTMVZTAgU0F2byvKgWSnzOFuS3uGkfzGpasiIGcWq
CzV5aLskIIjqAUNsiqTou8uX2c+JXoeNFppUaJKtUnb1eSvFqyGqq+C0FxtzR7QG
sO7Z7lABG5cCVWLs/ZXzwvYuuLKAjI/rhrHsTWGu1C/+NN3H89iifMis6QJ5HEDM
Qtz2tO1TnZR1SHb43rlF9AI4AWu1bJ9zmQJtVVTJbWQhFdiAIrbeSIrglWTtt7VT
0QYpinTgOLBh710TN/DTtxJVFTj4myJXQAqwkW4YgHpNDXwLCOY/REFk8SiLziCE
6RkDjc0U/JLAN084qHXyybcUdMxc585A5gKPaL/v5VHeBWN0/b3BnX/BIGY/R7DE
KNTIBA6SMtHfTFdCJsOvj0ic/tryeC4ykrP9VsQ5nlmWBs7W6J+FCDH3fLqGhw3V
WX2iC9r6rsatZUkH+PLRmNWP6yP0vUs5bery8KMWv4gysxiU0yV4Cg5HjTRtQvxE
YkdHuwHfblLVLROhVyXi9VQG/6cdDiEnYN2iXrha3q/Qar/I0qoVpHQHwTMPe9ja
txD0XYa1tiJMhRxVU7zS4lLWn9FHOj/6ZeBOXzh+NxEWoaNa2IWarY3KNeNurMBc
16A+laiz9mfguUprvBNPfSykn8KkOLheaLH5CaBb4/JDBren284wZ+ZGBQVM5FSP
4erpTQ2nRFO3yVjN7VN/DvOusmRwWwd145T7Yu8Nq8U23YLZ6yRV8UANhBs2faw0
YyedCiIlnWdHKAIR8FPQi72xGyRWEZ2iav5xmEXE9tGij2sTgydcBbjZsLju3XZe
F7rlvE8w+usbxLfzjikAsT71ANadE2X3XO00KNRJhxyRuMcYrmnQ7/dsI4mc9cxU
2p/VVeMmdml/8QNYovpa/WNKMsKCsMoUdPKU0i4ZOMSV90r2gYjvlFuEXuwkGe8+
wMYZD/Pp+ZDYsTGXnAJ62myRqTF2Aj8u4fT2VFnmuIfiRUXM9Zx+cRXfa42wg1sC
htcxpLhlffwLNdJc7v5EyBxYhX+ej2nMNc8qcWel4f4ceLhFXC6XfOrKtdvhCIhN
guXZrY846Q+AOyXdxkKthRCnLmZhySo+d8Sv/EAwkUAWeodYhttAbUXrWSFwTNn/
bOz9ocaWki9xZXEl3JR7r3IKuIWPdjGkReQdDWMWm2T313vYUUBqt0TMRoukCgt8
MCRVN+ensMCOVYauNPsOF9wl7oW4MwV3Cn29W0BExc1ioifCcO8DJsnqx2f7RyHb
Ou04EcUpxnrK6Piihhx9cjnM1b6et+qSXcXTbtrRVr6H6SGtSzzpW4ALUMiw9Xs9
W9I0RoGSgzzQgOdapKFV2I5tlJkMnL3DnKBuuw4mTIjfpvWhEn9Yw7Hm3apJF6vQ
cjH9oL7A6oI7eXnzhQwimcAlI70+II9ZxNlt5a3gypec4WsMzZxObGyulMvEyoh2
LsDHXUM+sqIdyVug3VFT/YoEweDUOIqym9AExPbdGk2KuVECMeVNr3ly+N8ETO8f
PMiI2LKuULum/yUYtMMpEQW7+FoMb45XXvfyxQ5B/8RV65ReSRBjMdnAnmocZlKB
5IKZ+MWKT7Jsi/Ormy9nP0BSkUXoeCHEbAtYZaUcdpU2SwOd+1b7qY/0ihgYtuu0
6gTrDinqyrpNoJkwIcfn2HYbFKrDhSU2XsPjvU9fbaS7SgjM5P8J6/Lc8rc1qyEA
vKortPS63DsC247O8qXZnOGw7t+bQY/iCgCwsiUKv1Y3FBmrRUb1XiQbqW+3OGB3
xmCm4IMKZ3VLmjo9+adG/BKBikKIoORfRYPxqgAbQiAU8S0+QN7S/+EmtL0g8EjE
6TzxgRlHip/OONKFbRYhtfRPqjZqAQYh6rOp4fTm7N+2uj0p+mCZ65/ClE2PrdAT
NZ9iYAVP4AXNtT56jWTOCpNpfLxKRaf0+vQGqald+mV/ODOvXZxjXQU6wnPkfuKP
thb2w0lqciR3r86nCHIDspghKY3+60lwh8RmisxmOiUr3Z1sxl/QzLcwWcxG1HZh
Yu9k0rbjQCrKqN4jy5O2y+G0ltgahM1za+ilVTJ8+BFkkHvS1Y0c9cZSP2NJS7Yy
mkPtKi4wwkLtkZnqdTT8jJeXu48Enys3AHaFmgbgr21EnDJ9XPsem27V0SiYsmjx
022dm6fXXESpp2we16TKup2l1L3lLgVhxXzRie7nh+WBmH47KMH9EQakakJKfOhr
YlvnElFZTmZj98SY0X+RnfxKhGvWpnn7QHXTba4uLWZuJJzECkRN0Xum+jxsEvYF
lnozzjl1Nbc3PSxCOphdU1ujFTDBP6A4L+OXP4BgBbK5wBvXvKtW7hlPYEzcd7gA
5d0tsGxy7a0GRTbzqmmFM8HIzb7aU0PIa6XI5m6vY9Wfpb3bhkR71QAzJPg95Q6i
F61zB+a9rImQuN5+vqmjUOooXcSbF4D4yD9aOmmnRSidGY5jCIlDsMpTIrv3rdgl
R7fQgVWA6ijIJoFyVOKZqL3utrkS2qKbH3ZGD82R5JT2AZcWXI2TPTBU7+hSDT+t
6Ex17zcvVeL7EIXqP6bburKI/k2kb9pLPuGHRQU9xJlAQO4NNoPvSScg8ZLdW1oB
Zf5YKS/y05DAVuysT8ChWjyblhbE+r4TzXDFeDA8IHU0aYgXCBdrYxK91lfsLE00
FO9Wg/OLF/5f3B3KFi/Xo3hNL6etlScNYdSK5tXBPAQO1oB4RHzgNLx0A30pIjgE
8JDhYod+jTk0v4VBTS51HHlbGH7rfy/VDUa+iPqUWZNIB8DScME1jYJgf1AWCRgd
JkWEwGGcKJVnYUnAKWI25pG0FOwlgxOvQ+3//sy0mdrs9va9BvcZAMd3fOI4MvY1
ZHy75J5g6eUbQF3dEWvsDXNcJs1YgvTl85iIrlbvF7WtWdjyIjRpPXpKPa0wYdbJ
TAY7WVqCT82+TrRGvEXQwnq+lIlz/dQFP/GGPlQC0HiGtRVq5qamhI2Zxs+N9UFu
heJq2AuONCRURjd1Aj/CYgr0EO8H7WuJACtxgxl8yVH1UYHvhMM5o8NDKC7ZV2HG
DysH4V9bTRNpmoVWW40xRDIjqfm3Yqt8ITeCKPoo2lg3D14HMyOqeF4/eNWiThiU
QzE6za8P32Lg7hUhdfoEp0ddagJDUmmnk4GA+88ht+tZOIMMO4PNKilkia7hoFeC
RP1ZAzkeFgH1uUCDg46IFoPTSd6IzhllR1Qft1Kv7hw1QFIOe3diiydsTUxXqxVe
4MsBHfsG3l9ksLwmqmBwvOpitQT8sK8CLq8UVoPj7vaFOap/f/Ja9ecQgbnXl43V
xipeNTaqjYqv8FTmzv5k2G//2ogj3fzpzwjH9ttOWTL0G45BxXTctOgeBOrooVOu
sShj7ptKGVM1qo7nnjJy+KQW/sJL/IBkLEXuNKemJg1ufb3B2wCJeZO5O6Ys8UTP
Pj4ZrLEkr/a1tv3+yp+DmHwJi5PV795vj0HBAdHioA79IHbXYIW9rG/O8Xx3R05d
3mES23tF23q4BX4/Sc7J7PxaY0BVfzhMMPG8vXVLL4fjVTczqMzSial8B7I6UN4+
cimNo5G85zus1Olc6WxDBWd8vCOxUzH+C7E51Z8/EVcQU/ibVnoMT3x/f75i2Ulr
xE/H/StDV4V7QdeMlaMVyUJ4+M+AanwPLVpsrbb7Uda2mBchwEWuf9DMPMiL+MJL
RINtOWkplB1FebCgF0AhjZ3/hcfP1aSxbclTYgNAHVoD58E2cdyJaOEr9IjlBgQB
TBMWlvYs/pv2EbnhFJ9QAGXCEg7Q6Hiv/+Zi1XSLH0TMcf9uPWSgWD140155J5WM
rRo2teaV4z/qUCfWxSwq0vaKGthSxC4Sqcg2B3Mu6HCtP44eBcZqCF3l2cFnwELM
RDDlPhYxVJozI2bbyuCTUJ4K6RHH8Qqem76WLSx4raTuUxquEIUUql5gX6KheqpC
vzq5vSbOIntdZ4t5NUNLMew82FaiD3TLKL0cPqFOpIy/E9oE3TDur2iQHCYCiMkt
spaa28ttfZ5FjjmeMxQPHiSoYMnCcgXk7kjyoQ509dpXFGs+dlnEFEumJbyMjG3w
pjIcnxn8smGRW9UZ0bHOroyXkWudwbGDOZhlIqcrKh6GgbqH/GTxR+aNufB8i8M/
CY+fION0UlXvCgAN8hLi6vXZ+B8k7am0z/x66edhjJV+R5eEoERYlZEiYT6fgI3W
aZe4NRhNf/+dvq2ddJPB8nKlnsp64MbamcYJLOiBakm6SvJj2fn+bzD+RA+mvKpb
ZqQ7G4xxXF7k18wrnc97/M8f57tYcWh3pG/VBMbYBvp6Zx13OZFKYMq8N6PctxLf
oqEJNZ43bPgcFjl9OceDsooDhGXIVuufW5WCySaP5XSp71GlOCeMScfCJeMBcTy5
mBRenf+jVuo4tbCbbDGFqqVUPQZaWARnheCxOdceaZX24KdRwOTbQD8JBm6GjKiK
qCHQUsDyg4Ok8uPtOH7fDBbGwxf7428NdptRvuSlqCe/kL1DNHqGNZGrol4vWr8n
iHAUBTk0fKwGbHeNptQ8LfszHTkvekkn7PBGvxrtKifbDGGnG4E8G60xSvWb/YUx
27NXCi8EzuICcRsEygTU5SAT2FE+1TifJHk5sSNJaFLPRE2vkYLybZpOW8so0ZvC
wRfcxHsTy6dbRPlIhoatx4MljbxdR3/Ia1ny6PF3X0uoD7rIfVl60LqIn/fnxDMs
nMRsztVS11O8fXJBY2Ero+OnB+YRRgJSV3YtdSeznszJLBUZxpYyuKI3J33pT85l
JL5UH+o0uAw+3jnkBYoEyuv3deNEQRrrq8BIPXXOfyB481iXJTbpYgnyzmDcoRnr
eXr3ez4aHtiFqEOabd5myMRsqNpnb4MgIzEo/94qNkDxmfojScANVSwSM3Rq12Ex
8jw+jIZTXLeDBgRplR5GHCnsadzJaCvZT76EvY0fNMnXZ/DpYdoq57GblOzo+gLe
N3pKGQ0ZWNHhG5d3sH1PqaYv/Q6ULm0FR8XnfJISIld0AGZ8N1zmFgaEeKSa+leV
OshPwj169afxJdi1B7AKCBW4GfOBZXR7hw3et8dE1oTY8DP9fKgnaYxdu4wHUHOU
ANV+fqwbxvzlMTog4v3O3KGO8u3VujHVK/RqD9qbnbXNAZLwIv1ko3mHqni7ZScO
K1EXMmncZZvrsEzEuZSlsofMw0tFYBwuw5j7X3voVpkdgBIARatUB3KvoZKdjiJk
0fJ/IdSTRPXnNo2RXtGVT1M33ZmnmZ7ztrudOxbgDSW72Gifsc2rI2F6vD3PSqRE
Ua2ZdAuSq4ehayueP00mw8E7SScn6laGClgtNKB0CEXE9oBQbsP6WZMbzQ6sI1hG
AOPVsNc9rGAurfxsXu7X6CarPdtGsqFCdA2IyZJuuycP+m3gZj8d8svo56toqi/S
7mz+1W7WWHHi5jcG0DNQ6952tcz2315hpPx2/re4LxktvipihJovX+F69jXaRvjS
dV5GFIsLDPaQXDZDxgB3aaQD1Gjt1bEhDZ8TgsKCpayiAF9/VFQfZBIWyi8CHQ+C
WtBiUpm1leFxCaYn0+TviQtKxeLkl4vZPoJzgJu/ntB6p5A4fkGpF7eQiO051qfx
ZM6OeWc5BnlmB8IMKYnp2jyDDkcbMpKca6vT7kiPLjJI7ZIuWQEvowNd7nCS1tR1
VrAPzzSx6oyFwnprF/gVbU+6CZu4O5GwcR4eqKFb/OxAnUrs7Ycnbl+baAUDnzsz
z3geDQ6CIdDyzbEvXPHiM2QXRQCZEYVzPJJmr1WY7+YN3E4TyIer3EhJo0MzHVrs
1Jw2+t/QHtZ+/DTPZzvudO4a3lKS6xIauxHXULZx2ZBU1eyqsRB/4RhIBOnTvs+6
dZcBF+vKQ+RVJu0GxlBn/2Z6diIF4y/Hn152zDbgim0srGAlM4M5AJDlWbxL/LmZ
AVCj2kShUNovaJUN0DVJrVh1oovPKwfCsC6aVtcy9w3v1fE623sHLh1vn+dXXDY+
akZ61lBoI8n8ehvROj2VfC3SVXtDhld6btfW9FkCHbWHJN5ZCYn5+44iUy3NZ32O
3DND5hBXFFtbPSJVFxA7U6aVdHWKO3gSu3pwR6oIq53TF5tcNscp7KjjR3ypsV6h
iiAGiKbNkE9qweEbfWz4rcGlNVUHpuuPFpb2Qrt6wNN+nqY1bt90VOiCuMNGV7y4
edIduhx5jWQxRntt9vl4MZaHShWbgHG0wwYN8xQYyPecQq07r8BR6BMbfDZeSQkD
GjGqRhZunxRvGp1lGCnJ+310PJaZH1mbDWfsasIgEZiackvGJmOzEzToyauInGnJ
F1UTNkEhDHOz6EVlZDX/BXr1NbD77zMBYb46faPAyCXKs+eWms8S4dQ3n8SfxrN3
w/2l/fFrglvfts5KV8H9ZyKuArTXNExHYxwEm6LxA1vuKpAtmT/yWnbC9CGUagMv
jndnfTU70BPdedPfxhrGc6GQxiSTEPj8H3NrmdZCgdreLXyzMejg7+6d/A8+4mDZ
0T7L5cuhi3bnD0e10/kYSOk7N3uhzsuKVp3Dqe+B/Ecy9+WoJTG637Ijf5neUT5p
Hu++8nWj9aJGiM6h0cJICQEZbTs2dY9M59/DFJFCDtQDbecu9f0sC9/TgcjeGK0+
vLoSijuWepnfH/M2JYfZInJjlnGUU1EPMqJaqJa2GP0nRRhZdOf1ednfDhgrAr22
3MROpRAmiNtuH5rFApd33PUzSesdkyB+AqYiew/VAk8QsGDgEelWYELuepjIGclh
ZtcOoKZyUc4QtcDmrTXjDpY8B4cnIOyHmvUCoz3IVVtDLYG7K/HEQ0EgnpiFLLh1
oaTcYavgqcI7bEgjbHssMIlVu7v4sSQvtHddxNnveBsRhLlbukRdfIqZKfimuY21
/BYcZn7hEfa7/QhUX5+mPQ0x3ugniueQysyoh0oi6Za1s1Iv05WYGFSpaTo4juk3
K8GALJ9SaPX7HWzCES5eOhQ4ICcfQZKQUYBPfkItYNDeIaUWZWCgyVR1x5IdnCtJ
yX4TV6qTraU1smmR6gu3YndaeJPyexhsJFzrbmezK2zsI3eAN4p5YFSuF5gkFnlR
zLE5anrGWy3r/waMRN0VBwpQSBEjuTp3Vwj3p/nX6jley9PhvSlnc5W8j9cd6mrm
J6CQ6glLbklVKslY5WmGBqhbSzjumsoluLy0plYoICK0AgBdpeJYzu9JgHw5lhQf
r8f3+CHx3yRZbV/cAPBXWYoRsKuwbgTrLZsFt04MQvDHh8Z5aIHLugfCi8tnxg7x
wvmR+XVZ8X5gj8OdsMuI/qmwcD1+MB3bcl6aqAiYx7//KTf67N4X3u+Tpb2GceVv
9u3KydYwldc0o83GfoXduL2sUCdIH+u68BevjGovBoRG7X0/UtUiQpoU+55Z7K7g
6aOZKXvZ3J91u89a1EGmy3R68e0cTQKaEn3Xz4EtstpAfaHYI45aZlIjT7djeQ6k
oTOuulU9Vdwy8BqxBlaBpzJWwxM2hPlly1kvE2DOUp3+plke3gBV5EYiOgH7Q0HL
Y/o3+6La5gaTaEM0PIXfwBRAmObUCzd0kXKxG1Lv5wDw3bBQmVTmFD8xVGQx0Maj
CIbMEaLlQKaMJJSO0gy5UUjxHQNOyhQOnY+BCxbv1jAO2E9+oE/XJ/keEBVwcl2F
vsssLd+DfTh1XLQ7n9ESqj+yAQE4gLq0CsG3/s5ruJRurGDqJUiI9bW/xBU6/IKr
Ou2SywlCLyiTXnqw6XaCsC/QCiefJb4gM7Fw1Srx9phqRHDF79MkZ58b2E49uQoS
oAg4exDO+LF+Sm2RNzn0pqjDUKBnWWc6yw+jiAGCdBHX3rF+ps9lAAUjmQ0wbMtq
+Ctku0mr2zGes8sjDmkE8H6bpomy/ZyMIb9YucPAMcfqt9n5e+7IIZSFIU/T4DiV
m/FPU94teC+V2PrHwyFhPt5Gku5v1CzHpoqKSvutJm7ybgwd7UnTaX9ex0AQhylq
ToLHkioQk/eD7XcfCpLxHH39OvPq9gvXvmj9eVmzTIoEhRPBvevBkFlqKJSyUzYN
1vltd4WlPs3jNOIyH1apzTRXSn7/LaLw8LNTXJ/wl2iDCotc9Ti4Oej1Wgr4WJnn
HvNt2Qy6nLTMVNP2PQeqSFnorsI1tNn5nvS8BWmsAALI7eNNRSrsWDOwn+k/Q7i7
L/kFjOOTxJBxl9GaAonW6XH/wbiKOMiGtAeakwQt1jagMwMsMo/XeHBAdiyiuLUK
A+ToExnhgfv6ruas5uVcXnxvtJKO+kaD7oh4XMvK495elNvxtMhbhpc+8NwF+pZ6
Z2nniG7zzFAQNBgf4cfrk5yeJ8IMDjFTQjIGP6CB7zQtLHOOjMUlfRiMUFUvznoe
sMfyb/eCL2gyOK8HezGwlD+GVtvAqgQtgBBbQ0UrcCa2h//qTP6a4Y7j7R36B6/k
EOvwzNZ6yNsOguOaxj+TRvet5e1BMMEUDNsPe4UAK8lAJFEcP13R4Wx6i71iiQhy
Pf77TP8tihF4lLDmgEKISc18iPSbl+jlAgZ8PpBLM21cLKfuu3PtmqT3N6tkIINN
lsTCA0nkd/YY8ExKBmjaVzmuRoEQwR7gh0MRyI5oHRRGsatpqqn7evJ+jQJZFI7C
gcCA25W2Kf5VQ79spqYyUKDF+Jbh44M/F5J7tGoKxaGj4ocPgnYeoaHkjzKRRihl
m2NE6Q1C3T9rQFdinGbTfudsx1asrwTbfFeFt3pyrfvMkzd4e87IhB23ocaE2N20
ReoZzzHVRBDBp/n+IUmOUdHwIDvgCzMDjFOgLk1OtJS6eZkMG/cCNNpv5MVMAa2D
tFURwgQGqH1uuaMQ8qaE5DRnc55kWHkZqGlkBALOhM693VojZF9Y42B48e6we9G2
pOq1ZJkXT4zKltYtWPOv/jVqWpIHrVMd/5i26VNnBoX8QXSHCejozTV0Ej20E/wn
za083L3pgpW15iG+kQAdMF19e5XKE18iioCBQCwQ0GQ36Ej60oaW0B1HSJeJG9z9
iUrQzUJyTZqFCLVHRgx22R7x7yUoLNx7OTOkdAeFWBiUgNZ8uTbdokDZTyWMY+pi
EqnABbhq/h7kL6TtO3zN8cV32eHGRp89tvHEgfY5oS3Nyo4ywI4NkERFarfoa5XV
O3ikd1dmczAMWQqJ1fGljH1bvFmUFoLLace7N95bh8LBzaivhRQNybzoVLXRz3MI
10EbS/7NvOotYdy7QIZLi6tI1l+ODJV17hi7BtdOQMhkPAC8gogJ5DbXn3nRRzWO
NANaE95JUNmxYG202zU4RzR7QFDr2sfnvXUdemUsPvjJmAT9nroKVcjrmwIE0R8H
/sZiv6wq7P8q0m4Fiwo1dcviz16MvlJyB06nQA07ZcSoy7vZlfexCPH08fk6Ezfv
mdGX8JXn/6xYEoTAXkJLOHfRNLzlBtAvCMq80E8Q2fWWI8WsY7Llfa5ssFOLRls+
tPOv00zaTLAc5WRb7ZeZEVIQF3flSGqw1fL+Fs6naDL4FF4XWA5AHuhQjN/HX/ig
ezTpYFCgZTzYYnKg9QEzfpj+e/KttVNixP0IDhcqAkDoNdZjM9TfCAsmrsDTN1Hy
RvJQdho7B/AOCrGIQ4oTX65MsvmbcZc0uGOBSGWJ2w4kyKR9fQLNEFWhWanQoehP
79uNCpGIVuoywScYr6zJ4Ksh7b/+/R8zwr6vwa1Ssol15vAA1L7cLT90cezN2NOm
U0lcsxi2SYVY16ijoPyYR7OC1HOmnORnvoXuTaRGQ7hoYhzUmdxc7HKSVnV6kmMe
XWXkBTqYhqal70dO8YT9m5qgK0hLFExC+ZO4YgcJDOwyUDtgmNgc+n4TJX1koAOx
uJesB+Lk/1t71TaLGKy0DgobtY4PxO7RxRrGcl4cujBucgOqLnD7LrbNaYse8dm1
oLQLBY4+8OWCilyuGk8ccXfGRNunRlLOFYX7c2ZuymMKR7LSTo3Dhb6ofiR9UYuE
XydupHi2cACWVPAq4yVL86okuoaDsWWIuHoFE1BZbNmnw1a3lwAy9efe0Unvg5ip
HfOyiMZMNv6uEbQ2yFx9cEhOoo5KZ37p2ZtGB1vzb0IIE6GxH06hxoRsz3MAus0N
RBapCCTJyFjwq0n3RuOEjkae28FwsMS6zc6UI9NVJl8Ro4rGAxOoHd1jEPPRjX7b
pCMZeygQqiOtJ50jiJjaVgcJNp51qOvh5XCQzJuEQ6H6m3rzdzzOTy+oFfBFyZlc
cjBM7e+I+En72vfAMVQosnkt1ITAI3As/nimnTc1A0nGF+fa5pX/u8P5iBnnkUzk
faR+DaVr0gLnhSke+J6jb4DocHuWNm+ziQqlxoMuo+ImJCXvlvHhZrsv9/fvIvkr
RwqMPNv8htLzJqWPESP+CUXj+i9ihbWgavxKrNfuaPeAeNmef8m5+q/o/+t20GYd
DJyppBv6ROEMeRBMJFD8/o8gui3Rh6U9hbpKo9KPeznnw1LFN4+b+iWAH80K5Xgd
2vdxdyVC/THLtnGnJNUdVqq3HGjXdkNjXdkhZRzkFCZ8yIw+vFW7tFK7v7c2QlXN
oMhTRvvyTzZtHBFs6pStIT/pGAtP/f4mcsBtHTx3Xs66BylnMiX8enJUunQoVe75
CObgzcJiXVLB+Hyz8A8f3K6y5XCsZKE+B30djzNu52PSKjF9zQjwbg602bxxsHIz
CeAutmBNNQdrzVdXcjScRmrcWIopSue1AYSp/XqdQ+JSGjTZyzNwAWV8YYUtsc+g
GIbmJoXpyqkfCW6iLqLOL/QHR4zWdK7AB3CQzglCBfgd35lHVvdkPCr8beIPtRQf
vlMgWJS+JkuB6Lhatk28nHp3LjH3fo7+cw+lLhGX5O8g6IfmFbNKJ7k4Oi8FbFq7
WmTpblFRhrfI5Oe5hjUgpHMc98MtfmX60sLlx6Awu+y8/FKrhDOj7nyPqrRJ2sLn
DhF+eEuz8HwFRQdUJwfNOsNuNq7Gwg9e7sgQeEkoCYErkeJmjd+pzVYdQYkBcdc2
cyP4V87krKFXAYrZ2DP3RJoH8KlCesC0A/U02ACTBpLejHdMMAry8rROxb2IxGis
LHF83EODDIppADGboP1KAndfT2tnBzAmWFdd4+On/hz+MK/4JcSsf7gG84XZnhq8
jwOFjkx3Sn0EW+JXAoGGweoevs0r/WnBqOePC/Ucl2NSAOu6rK555uLxO16LXz4l
lWumeJO4xJcMqcJABhrIZ8h3Vbnb/jWnAHUDw4NMUqfRSlEGO1ldqhtFokLSeFH3
Nu9X/BGfwjnWBIff1ykpeHSIHcKL4s+ICZsETjqe//MIeRSaeWK0PFWY/D5arwUV
dNGcXW8dLahH7Rs98zg8wn+W8S1Svk1l4w5TD48fjZ+n9cJV6n+jtzSOUitjuAd+
UrNxKSLKxWKk9GZeSg62xlPOBxPmzBxPM3C/6JPcpCWo5yVd+i3SlnLjjwtQm7iK
uRrlhpXFK66x1VqmzHywKz5+EzpeN1ZIkzaf3u+oIU8sAyV9Fvwt5A2IRYDJpdi4
HKs3tYV45AjPIVdr7CrGhVUzzK1ukCpTgax8uAmDpWqBZtTKcDpetJDcwR559LrN
yOslx8j+aMlIJAF4UyznHmpSOlpOvDZFTcwEf1LUxMs1MG2+U9yadnJuR94hJOYs
IMiwVtJrzrBbMGxYNS8q1qfnOnZ57Stwb59ik336XXj7Kd7W86zv+Yj7HqvkK2lR
p3KY3ESnVoSsajo1tdJo0GVY8NJc+Tf6+JSp5CFMj51Q1Tzv8nl5O4bnPQg2/LBy
/k+hRnRD0DnFHqJvoADbTtr1Fs+XIxUyR/xbhcT12M9254KlF+NNCDnbM7kP067F
gEHeHkIFjmXJsYTr0gmRIvCqDJMnedenk2OpeZ1xy8CMvd7iQKPVK0RFukApNZJ3
KUjF1rq3XoTEMZFrRth05Cp/5n8g9GBlkcW+uGA6D5u6UYT6PcCXVoR2GXD3qPTb
2l9HAsqULRvu4fZ5e857C2FkaH68LVBdYfdSP8ytCUkk94bsjtVaskwNlVfSYe5v
0eDhbsoLQwQWzgs9CdJSlOGkyHOeRXY3kk1xeTev+xP02CCoVU0sQldiSp3dCb8X
hptOyvzO8s+e7DpXfXJczCnmlrZQpq/yRTW2RkUAdy52mbdhvMk55STiUY6nWBT1
ZcS1I8wpQgC3DkekSoYzFPqjrogbBGkJ4HDXe3PhNltQk1qx3TtKRY8KzcGC5W4e
/uyuTOl8oU7Z9FgFjEJ2nr5nBwKCKbG92h5DuQDMINA476oaF+Xz4Ekzi+6rpois
eAKK+4Z2L6q1A0MHr/jwMU1IryjKXpmCV9QztnsNsxPiXdEPfmR2UVl9veiDxoRa
q1c4eBcWdG8b3SYx0jV8rqaollQIcbCItm0ntXkKu2kPKflq208YqqfSHuNangoa
uCv+Rbqnh8dHt5+8U7vOU1h5vtD6oUeKMw3v0g0nTjdF78OdJW6gyAdMoKINNgMO
Bio6hGR8XdlLuu6Ih5qoffgF44W9ZRWSYE3CFc492l0kuerMWXszCtOXXzehFUEY
6g3L/vaf1H5oqrJUJm31k59EMDNMr7/rvhKJSl5c647133zX0k2XKB5LylPQqBbu
5IVD1cv6ppRsKANMJZLfEmrRm9/LQGuWscjaXR0T+vfYKxoAorPhJ5gIxca/ef9/
8GTUAuM6kMMr4iJl0xl457KAU4hg8A+EWPR5ceV0wftFwj5/wasMIZ6ilIA/EeJj
6hwX8wbig0XEnIHLl4d0RVSbr/6M4OyCH1MTx4gWx2d+1QZt19BPReQCvndb5b9A
nSwGlUJJ5it9kLLbc8okqPJ0IqOajCKwgnaO3Ug8eNYE/r5rYC6szVaefs2ZPmfu
rDkC3VYvU3yf2q96g9eLjeqffT00/8bBg3sfy2pxyJetVwuYQKHjbhFc0NX1tO2D
F0SVq+fJyT1+609YuZ0+dXR0ZbyGmOEYLWD83nknV+OSIV3QHIRS47+2iy/c5mrF
Q9WvRukAd/L0v9iMX1fWcKiM8cYQ9A1Ba/xAHtGxCMBwzqM1dNrAeaPj7E84QVk7
9xHpNyqW4hsBy3OcCeEZnPvif5HteDsCZ53T73XuZXwviDZeYPy4LD4xqUH7YINE
n+hP3fWZct5IeaKE/hvrfkSvJ4EwQNfZ0WsGgTuFENV1oxapMmoRbkwxx2VM+YnW
Pu11aqIIJKMrPCJa1xm8j9me/Idygfh7aD6IyOI9R16/23nIbJgMT0h7N58CoQFh
Hc63Oi6TSpjbBT1ZTXbLLlXkze3SnhRJWG0WMiUTRrtBRqmTJr16ZXjKerj7rq2D
k/nyqLejNfFaOnc35E3J9gMh+fKWE00NJS+ApKpHJ5CH/UEoKktnrY+14x4FrDLK
wcqx2LtgpdzpuHUVil7WcYyJcaK0PKLVKZzVQrCb6KpJ6D5HEVV3eDLtTzaTcxj2
7kFcWNbrFrTRjzcygKy+m6bQUqo2rs01+mDhxCmXIH+EweYqGQWsG2QzDMdcRCZv
GIP2Sh9qIHnal0AjgG5IHWEbjMkXaxvDo1W0EayqO2xFk+o0zuZipZSPR9CIL49K
io8/MRYDuKI5AwicYe7xGbwh2E1VM6rfEHQAagPpdoUTYICEFAtaT4QxAVMo7HMs
CXu1osZSudz7RtTNHiopbtBUK3k5DIBSRKuCmaKS4Fc/2/99bNfYqzeBhK1LhTu2
j68atkcg9o3WwFJ29sopetRbT/81BlXD22b+kEzKuJnBNVBZlkbXA3mGiXzAE1N1
eWDURqzIsbD0BOngy7kpraemn2/l7qky1/+EcudUF9sBHT3fl/T0Jl+LAaqHK5ft
5/0MHZEOdKaxkAU3XbRCFK3ARfgO5IVDUkA7GzqgXySLn4w2XZkaFXT7heYQvQZi
WZn8EjcAC5PKGzHdmR3Gez6MZwKG0g+8+UkKC9qaz6Sczb4R/ou6or1J6s68F1Pl
P/PzNqW867+wRN9EZb/az5snmePM9S2MnqirBW0lXADWjNE9z7VNCOU9mSigT4Vv
g8AC76ikEd56Vgjal0nUnCA9OyZHwbH1EOUsGWHdbdUZC40UUurLKWg861BNPGul
doSkw3K7duihOpKV9zEeRmJlOZKnERKVbl9vbBWnN+cxKol1EMWXfRcfmLbJ8W+U
BhBy2IRXqI9cXAs3daDtTW3JPQfX8A4mEu6TVmkuduFulmzvH37h61iyhEKJInBM
O5/NVFELcpoDGEVonKdoE1OfzpYrRQRTr1K8HgSJyYdIRl2yFREBsRxAkr/zjQOP
70y7V/LAiyjJ0dQCqh2xXMv7yEs4fANu5TVQH17alLcsJI8Ng0Sf2jZuxAJqiqGu
yqyOh0QpQ1+guiIoZRoZQb/KPlx8Qf+2UEK8B8z+1wNmRvC7CiR8uK09TzMBL0TW
ETQxEj4PxAhacBI35Y0oGBw1vE8fdpwVIWC3A72uj21ZcSLmTfGOAL79e3I1JPX9
rnbTZ2o13otHXxYu/UHP1Zv2FPQq/5Mwj+WFSW93QvZEvw9tasL9ZFK/ngnONVCH
dkuJQ211Kn06U43EX6jJK1P9WxnhH11BlLEnLFKwIVIXHBaSiuayRTW2YVKEG5Oc
7BNiok8LsDQU72l8gHGMy6aH+goD8vNVo0x4+2r5rgWL5LOQJt2lmNLE2Y58o429
a6BglzaxoK/niVKW6Wd26wBmJXIM/ZwFENROwQKTGecSWFmHNlz+sDEvzb5ageUs
ZyDXjvP3hdPAxe6xr1u+qwuBkyFG5ALOfdRJPrYo5YiS13ZrIXgmt5b8yg42ShfP
tUDnIs+oBzuWc//dmkLYKkO92Bl1MqXPHKSIoZp0WlMfFPeGGdYTMYxGNPX1Rt1A
0hR4DUQ3gIWSMIemGF55huwEMENQUU66im27GyX7O0lkQfhhhmd3eU8/Imu811GW
DAeiOPikd61YvYf9zunhTFh193eexuvQsWjXalxT0u2T1540Xthu/MALvf0NW5v0
jYuxMiXpIMOLBA2BprE7pKL91k6M1vj7+7cvt2NPY+Z8zRUp+09groy8KC3EO65/
EejS7Ard7Gy8UHlNQ0+UeiZkeJtqNjG5uSfon+zL/t+EsbFK3mPUSWzFZG4nRLrz
flheBlOHDaIL8WEQvvQHv9icJOPDk6EqaCsDfiNBV0GbT1ONyqvyuFhDOLAD3ndC
vmjzq0BYZt6AgmXHQhpyMEr7dxUzISA4+oromMVaH8GO+GK9kiHS3z0zRKF6OGjc
RAkWm9LIG4lvAVxUe7yzNBRJzSM3TSxY4XdMwqeDX6JYLUmJAT+RKBD+apyrh2nW
BhlXizzJiqOcytbLPVYH0Ph7ZRfqwaUdQcSQKyu/zF3SU+s+1o81aJH0YWEWx7pf
mxpJI/nIqQWm9NWgH/hKavnAy1jIMZDHqiIjN/ipoym9C0uzEuo5IFFISZ13yV9W
O5RcchuO8SSk0FQDNh02n8fdkSywarUTNai985DLZgfejMxrx6NtbJfetHjkJa5U
YNFqhqwplht7iiY4ZduBDCHxDTcNUdC4ukcFM7eX/o3C1Xhz84wpCsr8jwFGrHTx
HezoRJ1k76oowVXtt+cdzwb9WZLTVQzd0eJ7vXDtHFs8Cag+jGxX5O0+HCPZlxEG
N83HfR5x5yrwHFn+GqY1UVOgX60+Y9Q1TJw7Z71uKFmskTDSfaoEDFUfciH8JKql
Z1lMnVYtljyaHqjt0weBpzxtqOV4KtdsB99+/TrdU4rnQZbFYbWrXj7jDlEO2znV
7B7OeSw4TXyzY0DPeL18gR7KRkYzQ4obt70nykU7tq1AYdoDWXmYrrPkV1lHwnrP
f5CpCcdWUwN8zIMn7o15lSam3xZioNl+gCXWomuZQqeJvnWRCbibu9KLAiD1Adoo
75ioOuy0ubwELzAnVZYZOeHw5wt0K3nG+Wj8o9zJeoj1vARzxTgFjkiPGibN1WhD
yPgWT4DF0IoSqJC71/zXoehBAvs5xLSc3fo+FpH5wnL6xH0ls3LXbWZmLF9wo6+5
wc0iqoVNr823t9n9X/Q9sxdhNT2KqsscH1kguY91buSbPXtfLSGxxLwqIV/PA5d/
dyJKvoGvFoDTdz2c976ByB+f6qqz/ZT9mGzbYjiO4LZXSOe8Tl+T21IizgWBfd04
OJzCAfDAETZxjoG38vwfYruerrQRw95Yjv7IoKiZD9rcWjmtg/hPBc33IHffeZXx
56PYya+mxnQPGFc1qI3Hj7LZupCb/icqV/dQKiCcWlffMndgrzF+DExcsKmgqYu6
XB9OpmJ/VVgTQSaWb96NgpvJIo3dXSSYr4xrs4r1Z6ol0kLCb2RygCBj6PmIsa6R
3L8+fxttp11c+rA8X/8MqxWcEmpZoYkZVcVautAfVS5mM/fRdl+HkmNaitxG0jmh
oPjIe5wpyVvxISG2TdIAFVWsaew7enGFtF1kTljaakupgs5y7lt+sjndr5UfVD+Q
gnZp/9vTQwNBYCBtGSnfIdCW5mEFelMriILkLIt+czfCi0o/I/WgW4ceUfIxEssL
Ps8Ov8O/cnlw2vbtcKZFJvAxdIuK9oKsjneX9EiPxUymzHZOGz/yg0j5ViSmqAC1
0I/fhfMVB+ZdOvuFZ5RdCYi+wIQ5ZVTOFkJch9DdBlAp6NFLXHlLxTd296HwCQx8
k55pvndxetM/H1aYLoEK7xzmx2ank8XAidstPe3unB/uEc1m1pEFvbN/BWlieVpt
Cdy+HNBAAEeooKdSojpJ+GWjqVXgLSlGlZvQlsKoqBLDEVl5rogqjwlTHLHxS+95
eudqt9Wx8Ig4IBKCXeztfVRCwaU08RDEAE010B9fsnh1YwUZELxcEqU125+Aw2Fq
37BSuOGLIufI2FUfMAOMucSx6f1XEUnBIyfRYpdKl+AThM1X105ZqGtSTSOWEJhd
W40FhgqOZEzwFKYwArgcVEeRxjVlnbI83W4Bn62v9+QOOiF0VsmM40pYhTimyv3A
Hx4wikTIRaQ5z7Tk2uRWLya4KA2uDSohllqS8cr3RKy7RBKYfEgvRAY8tgAnDgVV
ploqHSpFUK4cY4yNPEZ62448LKwYuCnRyRLOdrCacH4FTrbCXbWkL22P1dZfgscy
715O90y4/JwZs4/OtUMVOD3A3nfrqr/OSFr6NAxMDVBqdAMG0G9MP8PBf+6t8W2Y
oQiTol8tKlb2wijibVzqbwYEc5qXYeX+d5T3izOvLl9Dd5zClygvE/0yOLNOtdTK
XYENWMNFPtOxZOBtDQ6kfrLenOOHhJDAy99Ev/TlmyetnzNvHq1iXzGRWX4mOMxv
xt1GwW/gZDtzfqTR9j/jSnH9wlYinNffYt0BvT8RESIrdt39JED68YfT59tQxEvr
mQwfbl/k08S6Fj9HkIo+CEINwfBecfqFQZK6pmfpW0y5yPaM5YfzTCY+i/2bj72H
gAppgMj2Ds57d7oioAife2zkzO/dbO1NNXEL8fpBjXmjbZCM9g08orDe85VXUV5Q
xAHUy8TItE/GrYorY0e6m3bAGX2e0EHwp4pOxqQ2Iimj5SWboZCVfTHYRB4qamg7
qOoEry7Ho79nirXZmHY8qFryHrhWEa7ujEgDo5zMCQy4UESRxLgk8dIhWrT2Yj1a
B4tfq7xACsryhaJCZpJj2dW2d96Hjz/tXgW8htWyprgWUv3OSQHMt8SsyWGiTw5w
+z1QxBkJD0WQpiz8M0LfBd+YrogEUbS5/T4S/SCg+RREmGupL1659kezTesZdRsD
Z8ji8wyvpfxk6EvEn+vHna3Cb2gIHBT46Llh106aOXJwQLnlph2MF0qXToSmoSY5
8aW1hgNyQ37ydEnTj2QVQMlzZ5f2dat58RkypCM7zUEeXGR+3S6ZoAfSiOpUfhi3
u3Z99vLePGr3eR17rpMvllwamT5PwhNezjPe2JkaAs6sSrGDh9nNS4+OadT06vsW
5iG5uuqpyTcOcmeONfpIHueYeP/mFT5nSHBN5j6xtFW4FvbVWL5BJeCZEu3HUy0j
jQSZxhlmPezBiXm/7X/Vjjili3UiVkOOgX31pcdhpKYNEOMUl5/euIZyCmR5WnHT
9rKKLkcJ1YyHvku5+VbQJ3sPWzIm4fRodrs+UQ36ow8k4TgVv8VBBEjSydlg/s5x
sdKlA6vj73R3ePorj7TvexU5A8ir/4gPyTVOaUVDs54O0Xdt3TFXiDvMCC0rYI/f
Vxi0sX/CtkYG5VPJfgcSiA0HCBeb5O0KOOuO5Q+zD02YVR85d5gepGZvg7lsoTDq
3lf0ghPSefXKG+gBocqHcCHbvtzsjeH7lXplgVFu1sbVcsLAuvjbuM8xkSVyGmk9
gQGLoUIyhBSbj/2ll884h39f5HBXiOO5cYC9kiZD242jD/nKJjLqhk2+yPo+pywJ
HOcdzj8gDHunLX58BWsxbCPSqxqLEUlTBSE7YxTpSRRm+dL0p3IR+FX1kZ2D0jSP
MBWsHqRThvJV6V7j/xs6QYEZy8PDSkPr4RFGas4aaXBGWj5BDQY/OXZW9cW+TAle
6WkZ7JsQhm5kL780uQc4GSnLVinc4KXaoOsb8YwMeZFMZITHjA3D3hKJUVxWR3AN
ZXepl2xAzMULLQeSriX0LGfqDaANCRvxK8LFtYUPY5Fija7VmJFTveejQknahT1y
M7sF4hnSALtrF+cHHd4s+M7aoRZ2JlnBa/8n0+BLftryFYeJS2uy/PWfuFOpParR
9CKDhCYd18Hd6rSNWX02jfjQlbcuo2F+KIEx747hiULwDBVWidngu4hXfPfwuHh+
lzvPV4ggOxRBoRCCKsFY3oOIdsM5Vlg/bctHD7Z6LnLySIoxFZjkya0klYySJdsU
94QuMm7nP0/Azp3aKk5+RbXqUwrdcZl5R/amfTZ6gvYG67BUEi4gDSvj+SoZa1ZM
dTIorJBI8p7Um0EnklaDE6ITACOeQsI52e9tsR/qObuGgNPHIdVb+4frjElZTYPr
2jmo1ZqSpJbu7n0/vtecdusOx67PwHMpOwewZdmdfwDS1yXDKHI9Xk+GijmwvKou
Wx+zA37ZZYdza6eT40OAk+xr0UrkSUGN3Y8ZCYvAMUa6A8VvveLxO51dlWz/S+wo
Ll87xvvXkxWylLCyPXIgoh/FDuIDkFVO4qpqpYfLKwgWflABBTAC5kNciZ1SY5Xq
N4Tdq+AHiejZUGZ4nNrUqpN9vepYGGBRHUjrguh4e8TQKZvGHCUrBnBJVe2bMFLT
`pragma protect end_protected
