// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZMZZxFkc5wHtbeyo6YjI/XvADNyILvf2mfFX1LCX6qZURs2fzYKcJc32v6vO/I6J
dMGUwHFDbqBLj6PRKDMewbVc6DQYQqIakibLRXEh6fntPqKUOgtNcq+dti7T2x9P
1IKd2FLnrE0E19/B2S0OKIlcjldVvJJZxJpFOs0376w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20448)
4T/ISEZM/quBKzc2Jb+f/CggQZ6kEOLMK6YIxzEvtPJlJPKukfs2Ah4j4++KLb9a
443oBKJTOiiUhi9jQyqMSYMIfCi8KWegRrwsjbs6US5O2OR+3K26ZNRt1JqGh2+y
VTmZVH03AhA9+KKUxlo/QlaHVPiGerDh1aEK4fCD04+KrOMocDT14BLFe+oeH4VE
2x5l8OUnBoCCQ5au6/vsD4B4B2VOthFod4x1oML88srki75kYFiaiDEnVUlzJ/5P
aWfHuTxZovq6t9XWE27JGKmvS+aMSfw5RPJ+XrmIn3oxMCnFYOsXfHNy820mXjcC
CLXHyuYvj2yvvN4sSihfuy7X+pUUdGA+omzb84F5UC2ssQQ33I1GeiyBCiZXL1w2
snIJ9IcxH5R06mk4zYrFlWVErcxLEpY072lMmcg7LREeqn3wBx5SJxkAEib5ipuQ
hhu2pNi21g8y8o/Om5kTTICedAEESQ/LkggOXBDQnU2mIKrJRJy37z8wKmWGH/VG
VefLnAUMawO3PJ17VtWmKSmBMhFR75paStor2rIAJdZ8KJ3+5mlofVIrxrXW2SK2
XWvmpGPVluUJ/DA7tmmLYN7x1hCRmyWqu6FaFiGO1LodGzOHg66CvMbYpuSgw3GF
s4lUrOIpq0PmbE3aEMpYcv+U6rmgpCdkHwP+peSxiL1qSNrM8H8HVACGNNs87KfL
UXal1gh9MpDuV2aiU+4m3l0v5E7HR6ipxkYyFk2v7nmgpjFlcqKEOplUly12zet/
bY49wccOhDYCON0+Z152vbT3DMIMhYLFA6dRI2E7iv1swHLe1IyMm+iNf/gR0TEK
RMrZ9fnnr3aHl824XfI1FI9Dx9S7J63arQKr0hmj+ZEfNKuCvLrjPIw7WHtQ+BWu
+kSBtvtCp+XpeMv7tnpOhNnA4U5Cjgr+7pkM+wiI+wDp9xqIsONt5ATfKXIHvBuM
EPVwthrqXIWKI1ao7ynZcoigUJDNxgjvxus0ZXrS9Zs+m87692ejzE0ItDuEISn8
Eq8WBJCSnRSCCrQJHwFfi6MauVgX6n/dROE/gyTuBLOTQMVx8sWwsxqcNDoq03UJ
li0GxAU2ge5JcwAq1WC8iS/ml+loCKhnNMW+YfZFqLVICiFdwV9HYWiHftBJAiVl
GGxlLmQFTUCwYQyYihrriyr9vrTLNJXU6k4w/TMkn29L9t2J6iyTCkMWtW+HrqWd
4auuLp6AIA5WP6T4PH4uvP3WukhHs4MIuh9aRt6zHHl8WAYHpezRQnCLpqFjiMFa
FNWu+2yWIdG1lzSUoNGErObkKfoQ8BuNexLdf6/TdL/4fQuilwmO95IC2qCP85xB
KPkuPWfVo5kayHwW9uvt9MfM4AUv7z93Qu+z24ziH/Kvcs8gJA8GKJlfTTAi6JxT
227oJL4hhVH5XJuRqbnkJqpprw4WuZd9baN48q5TRvttM8/ni4LKxyuT+6JP/ZVV
/nNWGKvchgwXty2xmZ83D1lOPtXm9FxqFxNxoTMSTF2+eRysAhx0sT5nOjulDsPC
7muXa8aRJ4UKlb5D6yn+KE1HMllV99oz3ORcRbpThNw8C63Pk9CWM+2wVnwxsCKB
k2reAsKcTiTzLq9Hnpn+85M9wIb5PGVdAKvL/M3y6XBfgFL6LTpORm/LPThoxFBt
L0QVDfuMM+3ErRwuOKLfOc4P8Ec3+G9+f7CWW+LoJjuJBnPuS6FAEXhDXguYq1F2
Ge4YCKA1/QfiJBa8HTHHCchjwW1pBRz2SPfvjSd3wgvtuUTA9prO/+Hz2S5IQ8Fr
VvXK0hM8rq3ZYz0nZdw5A+1Uz+t5m4P9jxb84KsW5wzHce5rrwZJWVlDDtC+QTyG
OfZeR2zMouBnkOuWt5ML1C3v725IrfziIqcDSoklwwO6QkRBWQSFzvCnS2K0w/0v
Kczo0O8158btNGtMhq8Dws34YfvX7JREfKI+r0zbkKhYpEflHVGbrmhgaq/ooL2G
1tWgb0ci6MRB/u5onwMhQiloAx8GZIDCCwextXyaKikdU+6PqS1ArEYLG9tNofpo
u9lGdmllmdjpFzT8WgK/Gqslbub5Tx6ZSGnunZYbYshnjn2UnPBs0/fZ+mcRDngg
/VFaFpo6DSAkHQPnqt3vUxCkUjsaZTZbffU+KMDXvV+tZiLWLI3vHiPALmvjehka
AhCBUMzYKkITW1q1J/ZqFKitjqQ0hBRcF+i2QjbcFBAQnHoVn5wQmdPnuwWWuFgg
fW0W59EYk9BzACSeaJonWZI/sjmq0fThCk6W+I8kVQ2ADHglNTSb8nwVZEADdRQv
enRdpJmzYt2W9fH1jZjfMq4pWO/62PO5lbx8x++CgXy1X5B4DFiW2TPuUwRLitVv
TwaDNFkwZi1PV8fAYCnFeX1psJpYGRklz4jqzWq5ZV45KNCd3ZBrCiO9h7bhci8K
Z6nFUUSLjUFuB453Q56bxU1IudYKsa5PEPVIT6Ka4vdAnOKqLZgTAvLcn9GQqEEO
UvCPo26ztCbyhvtyZxIJJVI+eJNGHED2fUn5eCUsq4YKVQMVDjgEWhEBw5/xa47c
Iq5Rr7s2S++a5WdJral8m+0WJVjzjNH7mUktpX/FXLgcyFgOPJMQ8zN4dYP6DrxP
H8YXoTpwP/Iy39q85JX0FlczK04SBKNrUe3sMfFFh6rXk831RYYyBJicK0HtCnEO
UPg3luqX8iRRRqQhUZgHHWoSf1c1Fe30YvFZXrSNN9ju8+tvzPJ22GMSmLfQqGi/
V+5uve+cWkVAqw5LBQvgyRfs/KQGbi+0jXkMpAp/NZNoSWYSTMDCtQcAckuhNcsW
2Yrd7aT4ZXrvBvE2oeb+9CyOJ57N15teqLPoOIFi/N4V3MnVf8KyoEZ9FNh+UUzS
HXiTEEUosUoGXITV//l7ptBY1D5rg4EE9APpZElVZR+hipZgeVfNPYo7gV1/XcBM
7YOtLDZhAGYad1IgUieP34Id85AjjXOuWx6Vvn/PIhdBPPUNpFcRCdkcXEGygiPj
fmrRJVuMjbXXx7OSOiqT80IT6G3j3t5U/YIYdZ91w7pW2fQDPNL7JVqs/hKdKE1i
ILNmMP7pwP5kfuhfxrsZi5iJ3XqfuQSfAI+7Aorua+ibAebWxX+kFyc2lzJd14hH
6+26UUki+9HRhJHJ7jjh/1MIVeGTeipLtTSjFNEzxzje+OLwJvIJJiMpZqQTVVdD
qHSbF8BVmBMwz8de7UhxfvI+P24M93+xb2O294VuaCSpvQHzGfJjEoTIkukZvYbA
ErcJkWNajyv4rX7duSFr+62sCJaSlrFnPpJUPqHz2hDrJw0pQhhMrRIsEUT3eUIV
adH0jwhDQvsusFHWnzYh7RIk3cOl9+KZt1BKnBoiZpJaogKViXOmXPDHH4HT/r1q
3zcs8RyRsYGGHfagg/EJbtRj6KdhqXJp1vnJUJXHXeWLJHG/R4ZwNPrNpwUhVCb+
JgGMGPiPpNG/HkZZ9QSD2Ipzee55mrlT5jBNOvKj+3L2dkVR6Gxk4xWdgSpwjced
NLvDySL4Pqz5UheIldRWh2JLaUA7KFyrJQOUDPvue4/VnxrE6yNR3aR9KjL70lDi
Cocs9vrXx4LDsOGc7M0FEyw7kB+Ei856Yl1T+lDvUhhjjEmy0jIq0EbnRH9kyx5b
gj+F6QvREMI3Rvatgw/s2ZPZjICd9l6SV7ieroP+2GtO73VCaG7oBQiUhhee649s
uXRu25lQgv9joBs9cYPGjK/Uha/yzb1Og1Z7e25apqbN7wz9/czY3BcJ6KdedXTV
Hmyx3VJliYtAJzcuodTI95ZgSiNxs6L9Ibjn4fhMfEwepdml97uhi+P0MmeFtVK2
b0uM7whKYHSrUY9Lk1GhCmKb+jqZh/gJtK7kvbnATACb84AnziRZ0IVUQT7A8u/K
FAYUgcY+c6tnjlmoSUTOkBqsqHCTNktWo1euO/2i+2cjIONyW0j9gD0M15F8VKjN
JKtD/de+cjqiuWx801A7HZ/cUCoNj76J5fXQFxG5vMmeFeyRhQ/3l5Bf3CKnSM78
3W2iM2AykzmE/l2tS/EY5gfA7uapbLEbkKEdErI2BDFQN60T4HiH1sEjjsOVyFeB
QzkQHcTAMLY2ykS3+GXx3+1tpFoMrMsB/y8nhqaa4mZd31CkplFx0IGSqZ+/rrFi
yxnSbbq1DG5ByY4L16fQZpTMxAHnxabkhdaWSPm8qr8e9vHqmFHcJ9aoFidd5L+I
0pXYp7yvGg3HT0Vf1zImTyv1nA81m5jbpndHUQn35yb/v8aI7HbfCZcjqbpAMbI6
SwqE5IgLweQMbvutACo7kGCfWb2UPb0Vu+tDidz0O1WHNFKR3eLfL2vf4Axjcp5v
+MBC0JU9JrjkVdTrZOu/A+1IWFCA0RK1RPdCgaaGtq9fBEAQHlBOEDCzn3rL4zX+
Dg5xMkT5ibRghOFilubrRubRJXB+OQfDRCVMKLvRw8OY1vXGrL4r+yhm+ufAe+zg
4rJ/0Pvl1jRjfta0tx1qZ5An+K6/wD3RpI94VDV4R8ITYoKAtF9nllq6uKwg73bU
RYw94j4UNEWWQlVG7OPk6uH20rPJvLGXXIa3xsGsQA8dHJz4CY/v8sJtaneQYVMT
dPwLNQ3EUVOxLgoARN6FWBYO97uGBfNBBBggf3o2pBmBGz7ZPAJkLxlH81fHwKHK
w5MH6lxxsNEgwaEagJTSw7i5wchd/qRvtI/r/9AtLsZoZG9mS1jLse5iDrUMr7se
L9iosBEBGKpKHj1ZDPmbdtzLXbeSmPPlfNEp2QB7O4bXyUpGWGctNIIhmigI7x9v
xgv1Hq0j+mGf8Vc3QCXal+EGp2suQHucml2MSX9LJ/b9om7FWvoC70N8oN+UYSmM
Qbfyi6lK1KJqDKuGlKvsETTXS4RC9vw/Gu/jLYD0c6zbZlFCE4SzrrUY9ZnU7TCO
WOmSWZP8aX0k+LDLxGvMZbod+sbOsBlFrLvPf/CJAHqd0BMEwKKotz2F+zBMtyqj
4IloHBByOO+r1zMF3zkTYBNqmfJx0FWvXhLoWo+TG0YWUZuo3sbA7+3usFTbIwpe
MFNnDCDf1mwjP1vVqbcdZLXrN0CupVmuYWH50U9YSmHSl/rlqGhrP1rkyyEXIe+5
iuTvoE510Ajb5ogwngCmvF3cLfd5tFacFUgpLACfTvifV6bWDnq1bO85iQhrU5E0
7qku2KrZQ22TneNlhcfEwir7Dlh0GseLishm6AKBWxHLyc6Vlz8CroPgZdeGWYPZ
hrFQKajnmZXqEnsZBvKGZzkqjMpM8dUqdED9OulTAuFswfKrL3AEW4G/0vj6Rn4L
K+FOzJFmDrkNe9foStSpeh0KdfuNl7oZp9aX1x8o2nwWTjFS3G3OuhfNXkKCegmv
haRs2okiasGPyLUFzB5zJg7XNaJpoQVxgWX5Exzp2UlEGgrVHvpVkBo5b/yHm+A5
Fnsmo0ehGLE3erGzQrHfTPvEmE59rkbQzX5ym+o5KREfNW7JilFdUp8KEdDMKbI0
QKxH8SX69D9Cg6QurxlB8h7s2P6pzlVDPFYiaO5HP6My0HMnzYILUzCW89Ek48dd
ntvj3RXhGp7Lk+Ez6z/JadilmKLwrdIqnR8lYxSaAp81Xg1giPC9iBe0YZ+a0WJq
PWL+5uCbstJAqqnIRiGbUQyjxllTU63YmDuijdf4vMjTxdMYzAyhm8NIBdH0yqE0
hnMKxDz6jDx0Pdx7cnlH3Q0Ct+33WTSP1nuz1n5U5EnukI/37ZbnKttucvQO4D0T
c+POAQBJZrmDurSGw+fn2m8UPJR7BI1KOld+5TUTX12t0lv0rIoduRPHkvvuHKkK
5v7geys77+ybdgGR8Tt0Ywkm/wN5/Zc7n3Fzs0V/hsGJi7sgIBhNOgaGxyeI8kYZ
wL1FCy6tXW2aQWPPCl9wkqsM8iK+VtZbnGrJJIRGqYVWBundtZ4IDIunjuPRqwPT
r1CXw47FTXyoT0rX9D0wBhx39M7PzbnpUvige88gbKKwX6azpgaigrAgYT6PZ5zm
uXG/ZlGdWrefanxOsacJey+9dvzS4/LQTLMG/JqgTibNij9SggWZcxGLdALDuQSZ
89MYxn23AezYiiYQ72fcpKyRlZhh7/d/lFinHiMkwcgGoySgVok6pQQ70L4H3D7B
15hX7bn7OVtWz8P1Mknybmwtsy39fgHIsDyiqhVoSNpMD6BJELM/+0MV0b59Y2F7
4P6CCqHq6lYkeOJdoRLejg+tUvGyJ4eW1xLkO8+Wuo8UDP5ZFBk8CMrUf6nezTSW
6EGzXX7fTGOrcVwd5IhIX8X7XMLYkwriBPXO0exFB/IUIHOYQ26AQFL/5pzuf8oS
bYGbI6wDNHfmQSqJGn6q7Ye/VC9Y0FOwpetQGB3tiFl4JIu0yDcPzg4Cdw5R7saN
yTaNWvfaBMfKm5YwHl8iU0HZnZA6rzWhFEUMGcA3C7Cte7IHZKavJLR1HeDvZEvF
0mKkmF+5z0LbE1+hyzOxKNRBhWAAjUMir1ZGmDxi75ZNXKIA09vomcQj2eLwzNha
bCZr2r5S2UMOnpfoXHhu+CIgwqbiNVPFQ2FD86oxS0kXmNeLWdjaG4O29+YBkkWB
kh2UoNxc5EswqhMn68deyH09dhQ/lj0B6mBivG0KjMJ5MYQ/JRAdnOeYQJkK5VHT
WBKOAgQctjxVp4OrF9UedQL02XrLOaPsJqUVixrhqtRmy1sb09eOKTGV+enXWgI3
8ci8QenZX/TweDm9V7UOk3lMMy+zFro1Kx5U8adDymWyuBPIgGtLTQKBHyRKB2YV
OXH8adrTsQZhzHJuMBoucPve500VsV9B2Mybf6tWCjdBk/dAuFyipeBWqCRDyu2h
7k0G25WQVfpGQpDXcW8Zdu+xdh4HC09Jr6ZG+3jIu8EIoQ1VCZtF8OEUPOK2AvoT
2+fe4dQdaLQtTVJMmfqOx8XwRIYlbvspTcoeSjFXr1Menvpu+5uVTQjo1qIaJPRg
2/muLz/BXsCZXtQ5JBuGC0sYXS2Tke1eXohKMsBj/LWuNiaok2eki6B2Uh1L0nUu
a/xsmAOLelCwRm7OUunTrwS+RAC8cdrsxIj27drNyVHjA+I5RyfwThTCReJ4ox3d
vR7+J0fsyBTT8+SLrIm/MYtdGFTADboyeHIZXgi8oIQ7EXVuOMwwg+tJT+NYFyUs
Gep7jYWvjs2ZnxVkbkDYCbGYaMqI7rVo6kQc0UivLrrMuUh0zX6Ha/X4W+HNnEL8
2WPkkQ/Ni4nwAptipJJma7W69fh5HBzCp6VEoGqAqvQtxDzeT81bsOJMhXzjSMBZ
8SPjGjk7Jyx+4ujt5zm0NM7xC8ZCCldXBYNzOrbhD3wFGdsfjNKj65L+2mkKsD3F
cNQ+oDa0ZCX4nPWaCRuB6mX4J6F7LNF4iF4oGXJa6HPToPK2I5brSEQirmlCf+y8
BXGpxDriszvqwbIirMHahpgxxPxs1605+EyQ/nWqatYW+J6Hfkc6tR1ByEialEA3
DT/TCycWVErPcGbQ2UJ+rS8VqubKiOzH2KY5M8T/eWxwMM7XkejS+ydXphg5WYBw
po78Lg3eNABbqhdYMBed+r9tFI4lT4oCj1s4vGZWXmx8eOYp7APu2h1pX8THlxAs
aP3sG6nuVRdEW1WvQCrCjjnZnSZC49fPaq6Ba0TI+jxA/A+IKXGLsblkcfp9qGKL
RFR5D8fdcSw3c7FcsoJgBflOxCzQu/I7qUeyT7xvHywRdZOMT32jU/QQM8P8+RyL
pbl1R7d66dRogejKb+AGclMtgec9TsLAWE49jc02G7TsXcF3ntCIhsbReOGoPV0N
3bi2/ZJ1lnCxcoIQdfKV/AjLZjLD0s+72f0z/BJSrsbgXrA4Ysdwuk3T1Z7ERHeV
4Nr05XjpduTQEuTM+kmxT8FLST+vSZouc8tdVNmKqGGrYuP0HttU0Xv9rhB0XZ1U
OFfnMEn3EXqG1zUrZixoFFeAL9C0UYA2csxYO4VwIIa+0asaK7ju0Ex1imYXEF4q
ST6quOZfMi4fNAcawAnPBAEiF6rV2lvIE52Uj1SSiPQTSkxcY/9Skr6lp/+k6Ch6
JDt90Y4x47RWXt7DduZchT/0iJJIXR9BeLXeTdArYxD1zlm5p6PAl04H1xsceCJw
pYfiO/IH5pEY4Gv4G/sOBTc838/X7jXCgxNTB3qhtmk0cjbh+a7JHDbcDghT4+d2
qbf4aa3JapwZnqoQ16uRqUYpX1UJ5nl9RNRBxbVlV5JICs2g6jEZW7tQlJtaathe
dvcG8wUpUU+csCDUjOCEgX/7Nxn+IDfmYGRrP3Ro4ZOXhbnZrhh6fEzWHoULkbSB
MJSf/WLFBDXoY2A8E8qcb5u/fVlOyK3AuV7iSD/cqQD+uZ4q1/gqTyTEp0JfN67l
alf8ybxMMPol8bWDzOgvdDkTq7EKiaiW3UQh04DUR84HbERzvklYTurJRo9FaMeC
tL6uPx43N79VUgX1eztuYJehprro57dM3X608mCjOgU2Or1XjjAxcmije6JjvnB8
GWhqZvkxzVyQdWezQ6/XlaWJkZK9YKWhAU/5iNKAheX9irvnTCILSGVvdKmL1tYr
xnfEUr84iWPrDgYroCNpaFOXObb3R+lvvtKWfnE9XIb8PH9IO1JmpGYVu/iH6IAx
uZC8X+ipL2PvGpuPO6cqQb5cswfVgo7jo88NrqduavE4OJfhzsn6nXd3jzPn0RLJ
JEyWjUeQMwQNlJBKelE6vY/GBi+1/sr5hGDJauoRSFYk9tztZh0rBlgAiC5rB9ud
N6we6ibB40iFrnyuV+wQl13CuJYe3ygLTBkqAi9uL6PXfVYydUmW6GULOc3JhuU/
6t6C3k7bVu4x939phKB3mPjGXdXlZDp4ocMR5YRN1gMr1DQehtAMmSZ1W68aFOPF
0I6xzxSOqUAeXBA3wO8w+GH974n52enTQEyxnypASumxdSqWT/OTTTKeV6VOMhpQ
wpQu88Ur4XQurbbamZOnCWxckhdR0fdtQT9mQQgGG1eHcgY/6losh/oducFVsLE6
4bf/igP5CF55FOmV39RcBU1SJUMZj1ZQfeK6LQ2/Po1wzy+tlgxlmE6JD1B8KBzL
3Cx+FAo93d5NntXs0DPTdiZt3+5rVh4KyO1hY+QO03l0fjfz7afCbvicvar4soBG
lex8faVFFP+PxcqHFDERBzXlTU610+MY4wO2i2eeRw7JAmDbYzTiywC+m87XOupE
07KpP6OAga0ulVCzm6jWS5g6T0KPJUMuuW6GuI4Fsb/ICsv2iAYUr843Icedq9oD
u5iQu2h70mWk0kgzFVb5DcX8JwVAaSqWBqz2cIUGb9l6iAhnANZBiAXBlzumFufW
pa1VDYUP23IahOsCIsMlfgNSFftprkCm7hSbX8twAOoFbIQyi4ekuH9jIxWLrteB
rXbMPqxJ8duPryTy918cSAXAmPuo6IwdBjGsy4So1t+BfMXbrl+rjnkPBIvW1yGI
3IU/sHNohU9zJvJC+UPSNEYDHQLaokJiOFf5jvww11YSek4VrhC9lC/FuugN5ZmF
s5LrlMIv6DCespAWqE+XxiVDqijNLj5hKXVP+N6UamCzntmOs+KR8YDIzP3GzPHy
8u7+lW5evg08w3JVrFcnt43Hgnx3sb9gxE+G9+Bh+vQGP446GdQVhefYqR/GNOin
CX9uWojHlXv92MZmBSkDcnMcT30HBLf38q0HV/r5f6PxJIC1qFMvBcIJxo6Sq0r6
jmabtzPNwEguStsRCoo5bATgQuSjCYpAMf3WWIO077JZNGxjuQg4VHdacphXTq/I
O964+1RSMcEo15BiZgwrTkkRKmeXUfSNLe/imf+pxRvNDKwKawOa7iN9hv+4klKc
BxYfurhZmMs4+VU2rYfLMi5OiWr+2fnaIGZ79AZFrSPgoedrdB5Ykg0rSujLWAUy
cLu5Pp246idfK4yfz2hT+OW5Auz2UQtE4+kWX5fEDY3HbKGffzuQh9hnQ1nWBZSH
dOr1wVFIc3bzav/M0a4kTCKYjpwtE0VFuy1p6CUE4GSgQExwIEtlYU3rFMQLttDh
rvAfFIH9XDsAUeMU5S5BnRltZy90mwB+vuFqRlcP+RrOtbrmXri8dIW+O9BVmORZ
q7aeX57HWXRLCTL4u0EdEPJjtxrNqBmC6c7bs3XNc2QsJshiAtNOlD1JLARgHUzg
8liPIcCWO+N2hyA66xo1qHbPX5XlmW/AIcaqAMzyYcXCpl5MT1KxBNe3pupbpeAf
cgzoccGfADaHOnCHG6Lvopn6/v4wO8uA7KLQWXqUD2NGZEVAdyOdUuKjhh9xAGMU
9cncBfF7IOMC44iqrzH2Uv2jReiBGafvpUn+pPCf4+B2ZvC2WXXUFpQoQZ5rRSml
OKEv0M9q3R3ioSlL1jz1RuRJ9IMLmV2F26Kd6+5F6ntpUE2N5iCMy/TSnun0LtOJ
ydPkFWJ8rR0eyXDjvZAOETES8NWCpvLhzmOHed5Q99oDLIwbDVXF1UhYt6NzJG3D
1004P97S+dMxG6jeR1h9KsgFqhRUrm77LEbiI7ORKHtjIVYY62XaPNZDkWHy7+J0
FDcGhiqy1b1rnArc6Shq8Xc6y+AxY6oTpXAfNkRH1hLk9lst25Hrsd+cXqcIoaJY
OE9/Kla4GTVbdE5KBTo/OQ9DrjQO2C08Qzt9QbBao4k31vDsYNVeynRBKqUc6jaj
Nz3pjGshtg2PZDefe+qr0Z+7pHIM4SeW3SuujnxhcHfYgp5b6R235jUk+s8Lbhil
1ixCLYqX2dMcdlFgxptyOK4T88Dnh2Hle8ZWuPU0sKZplGovwVh8HoGE0CVSlJNj
ZGXPnznMVUEBaRx5hnkWJiVk3ufKKBIKpR4TnkR6S4Zfjg45IOkX0bpW4pqXBvi3
3H8Wkylc40TeIhc8wpi93JwTms1YMEgIGG2mfBP8sWP5X2xM5XxaMmiTHzdqpb1f
qVoll406XBgbzB/L2hiYOu99CWmzSs2NILnl/9+dfSsFIhEVYfmMALOuA0uscxXM
goP2uXQu7ak3Kb+1z7AhKgG/Xu8TzbM2oqrksCKq8+/qjTSlh4GGlOpM0BGGJe1/
XsWYzjzOOENhG12+t7gUFkqYOun/ALdZMEbNw/4WifITl3IPtZMATYdLJcRgDTVI
1hxL2lVZ0q8AIT9Qw1HuaQ6LVoSde2LoviAGX7RzAC9bPDwPef1fz8rsdFgGsiU5
wQJN6hC40WCWZTm0VyOY4FnR4F47UtVWlOl5+cMJdW3JYlqGalk1QHxWhsYn6e8y
7dB894/jHvTbTyIQzU3BIAoXu9H62xfai42s5OlPlWuVhPGU2R7Fsqfj4BZrX+Mt
euc10Hj9KYy28IemVMNEBfYgjYVpJlJg3uYdgs23du/Db1wlSPuWtFfS++uXhAJL
dP8nbnQ9V/fzQgnvEcbraUw8IqfAB+k17Ux5Ni293mOEkf1Q1c75nljaVfjKXpTD
7jPjYfpdReCGBdhCXEaKv53jv6k4q7AekINKgdroTY/BrkWV2M9Um8FiAJ+1XtYz
Wqo/tI033xF3G3L231cZyCP6NwEGFl8+SmQSoQ/yF6IL/ys7vQcNRWcmXphmFwpV
81RoMpgPhnT4OdE7+7lA86D338GHHFz2yuoOyLYsJjmpCh9hm40tEcrzFb+gKrUZ
AhyGGJZ0o7Ct+dvbA2ZYOGoYaGcZKcUKo3eJ2nbBK7KGKaVYpWsJAZR25sobOQGv
7ujnNemXtxtEHbtdTfhi037LHPyBlqQi3fyJL86pYh/EBqkahuybKykTCLuRk2kQ
bOYN8beDBpnXqgMXx3A3f+YjK7zTFKKo32/M7CgkRq6f/clroHKev84xZkZRR60y
fVohMoGZkv4uN85juaOhE8/+bigNFC0hCfj7l3rgN4Ik52l2gn3oNqcl4R4dMhfz
4rMDtvW8+YNAFP+QEn0yXT7e7E6ZLeowXdi4Lk6Y2zLwkGyYUuUinXxU8ZnL3ojp
Q2YCppzrLts/SS0q6M+yGHK5IWWjnbfT6PWXyl5ka3zSB57To4MEy8OPCW2Ic8K1
KVJ1BHiHqeuUiNpOwX7TEV+O1IEOVEsT+lYtY7IXy4j/A5yGFj2PfqGv7djj3/zG
LzliQwS+LNdcIWwc6XzfgjJBbX6aEN+q/W2rTdyP2WvMghHCEDQzc01ytatrG50R
ipI9S17+L7kDihV2UBEEpqo+IF/3bII+QLSZ5vFl9QOcBW9+WbSmc+rjgy7j6235
iD5w+D9GyUCYXACqQFSw8Rz/n5c6Vs5LvuJBPnAQoXK0FDniyx/iIa8Sf2998t2V
tmDT16HaO4gYUW2et3koQp/Q13B6ttvTnrd5wPdYutxJOia5iWqhcRHYJDiygY2u
jZio1SUBvcPnoEPuj/u3kkzMwoeUrVfkKpYYEAmiG9gmlSxRsfrGyUsTESo/7QZU
wNQpJX6l7jv1ultr6hjHRkSGWW8CTcRzxfPkCz3U+5UkGhj/LhnsRzuJrexUhDyQ
7B7ebz++hhfMN854kFpSoqrZw1jxkfdwHBX6E82zH8ZEj7HmHQc6hzKcIku3Q5BZ
cWG3MW1PnY83sZgl2I5dNh6D7pvT7ubjOUvQSgNuj90PL+sLjhhhLEsqbjYmCYzb
0m9SowxrGpysfv3Aq1Rq1LrOUSoYEp+6oN1yk5jL2noU8MwlsrP98xLSRR1XoJVB
EQc1xmVkCv1+iWru0s/bi9RnaLs3qECwmtluRetTf5yFQQDs6Rn09oyRxHr4obDJ
v0lIYRaSEUs6+Wy5UJEI3HDnSCn0ixL4umm7CoqsqOnz7porPj2nRG/ncydg4+SU
6lP1bVcIKP63Ozon6+/tFM0rdKwO5bC8zYn48LmM6HMa5qRvJMSIXyiHkiklHbh4
H6m9pJxGrt21u8JN1MzMgP0Fv0hBOZiMmhCekdQzJEm0TkuNOTIMVaI0VMwCygUW
fvoOKAXyUzbwcCF1yMpzN2358r4OHJW7Odi14b9J3UGcQAt7CZIXc0Ip6Wd8Z3nT
M6bX/Pc7LOiyMSFHW75DHMkQv4OXhfDOHH/vuyNPR12PpY5f6UmwuV+wI5HpiufH
9KRwLkyAxo03pBl/DJRGMIAOMucrvF0ZlWdY38z1W8X387sxbh8j+EqwDIib68ii
G373Swby9upUlPFp0vVWx3/dSFY+aSjxzvi6MnmXPH2va5pH3/OqK6FqRu6dRXLK
q/I4b+wcZkkjUGwk9wz2duCEDC8iT2dKcHIpP1x8pJo0D+4B6xM9wyV3RYGU31x6
sLx5XKzxmyUmeXf2FryKKIf3rmGS6O9K4RlJeddgBKyQHOOvlqUwasmJ4hE5ucTj
IDCBUBUQZR3bQuhx2h9EXXRTRNGi869QBmUyL1QqWPQpCK4wm6DpWxUBiPjI3vKO
7u4yRsS31rjeqM+4+LUva2UsRxBgGO+eI9rICErjU/fGWXf5yRM7+6XTzMl/Elgc
YvXjcz1eXzW+T9p5hpeUQ3jsO55/w+ptoN7527t2Okp/lxSF4OnDfe3EggYaXspU
TQzxAfo1X5Egu9fqgJE/TuEjFSSajwIn4IIoP58iz/Q8ac6KnSmM6kuqOVq15XZt
GZSxJ4SxtKRa15f0njWKrUIB0j2ipu5OkrNoRODYcOsKrAumgz8ExkDKmBKcNCTe
2DGnpRaIP9rYt/5tmoXL4XOyuG9yhsvxLRJxZiTI1yUqYfw+ZNH2YIhZP4L4GOsQ
AM+U9NPaWni80c21ICRxUdayL2/KYxF3lSsZ5fN/xhpEItIcsiIYtHeQZXZItIy6
JQ4p9t3D8jE8RVQUN7BikJPQsxm6mjUCPYjvIsyhfYnXj6tN40P59SFZSc3mBnBN
mm2K3wwBDvLqw+JvP9d40vW0iNj0+UxtnmkfzbxAIKcpreJ23HmbNC4NnP2sfkyR
VF6Tw/fyOrkMoylAxNyFaDIkKUFhlVLDkOJEM4N0Au5KKlOpV8lQQ/2fJK8eJQT8
1thcTzGRbGH7BmpsEjmkaRVMrUx2HM24h2MmtdFfQmKQCCMq5uU5L+ChB+I+C/5t
VrJ2Rv4HTXMkCbNbcTXCRAnPvxEZr1UiYFB0Rftjl6HYRJe3J4GNlRSt/UNuRVsR
BLpYznLIDYWJEYUiic4MgGGJRidqV093I6zq8tAsG0Ue4X1QbKEhlGcPDMr7lNZL
hiF0t7htLZ5zEBY0F17seJ+TUBfTT2N6EgG6irt+nmuN66dqyvB8GE7ZRycv1xtB
Y7I/YIWNxvGTyI65FS3FqZxYPh7VkUG49BJgJomvuDat7lPpVZ0y/v6V9dU9kH1B
988NFmS48mSfGENn4HVKGFOyx1RaO3jF0xwPN0t/y3Q4Jw2ydTwbypKkiCwu+d6V
axveGYd9dOuTDdc1h9Xy5Xb4JjNIjdLKlHPmBdVg6EDTB8YIbQ9PH3OFDX+GBRO/
7DcUAVxpXib38aernQkvyvvdIn6llHvIrA9Yzc2L0h9eAdPL02rCVHMuFg0UT4Ir
3gN0Qu4SxgrIySj/VYE0yk9pnvefMpdPAzjT2ecrZrB3LXmEHypl+jhIR44kDpYH
CnOcofPrFSu46gFw8wa7/LttOeE1Vytc21EjDTAyCnxurPx8knnnuYxSSCC59IyT
+tTLxdN2sFZBGaVYyn3VXGodHHUuC69Cxl5bQiojBw+f1wsXaYlJ+0CSStaXJJw9
0yQx883VDXURvTJBGgDqH4zDsA8jziFnxsvfVJCZ4DdMs2bKJF+x+3Kk1BWGcgwV
+d4z77PtzuuuOB7MiEK60WMbVVvS9YR6vHJxSxO89j5ixpTAUXD7lzDmgoI4N+Ck
AExW2okLprnQb/nZy5Z8sk3YsQnuGkfBWU0CSBVQWBRSRlTYx8gHSGWgY+fv073S
8Oj2/JO02WbIq+jwcY8X9n562y7kzA/2AFxfKEcLFZA9ZwbKxd0Oal28W/Vkz1Fi
psD6yoM+3kpECIa9gOdjCxK/PLUqbXxqtGr86EXgcGB0PxbWnLhDAxc9WZAZNxg9
3edsbzyQP1NEfgAwRcbOww8PBto/xg0MU/P93c6fcQhUmnt9IAyx9aWsst/tbaMQ
rg1v63x81SiXU9z5lctTjIxavzZhVGH1H8mcQT1CNfr00qbbbvsdhIWDD7ckuZKN
EwrU5o2iC+N4R0znjFwVhIddW3fOqQDlcDXz/tQWQ20j1zLN9N89ogg4ixIrN1Xl
yPdnQB1x39loaxNcdHGRNMPpnFs+SxF3Ec7xhr1HGoYCgrrye2IItLDFhG9vX0MT
Jj42Db6vgnRTStgqEQLCLmWCQWBsKFeVpaCoZ1uQI+P+y3dVVLEqflnn+Z0o+IN9
qbb1vtwjW+ENMl/OR2iKJyGid0nd7hWRBwN59hAXvx7cSTUZvWauiWqe/LbILCbt
RcnVl84VkygqhIrmR/LpaKfm5fHMWhi6GMHM5GmZMwM3cL/wpnyTmRzhc73OIiwz
8S/SxIrwbv4OZ4dfqQY5sSgTLymyiu5l84aYwErMF9t9eIWh6ErwkEYkniI1pe21
zjgtXUdFsqwfWHq4sII//z+mFkYXJTS+BuJIoZMaCPxLj/mL9E7Jmq/jV7legAde
zahlZzsqODp6MdUUXXXAyfMelHvNbEhvyj4jHw9JnKmCQ3+MsRa1Jmug/lk4acdC
yarJSWohnsgd05qQnH4GG7mOok0x1OfwVRICepYbIcmov8ERpBvmaWLTNUiySPo9
IA9eTmHzz2raflU7FiWHx3CgH6ezuAg5ew+Y1PfTFX5qy9HRQ8lX+BdV+xIu77Qm
5ZigzNTjKbCJ0E6Ychxoy33oN2pUsJZWTQuZmonVH1zcdqQGE/FcV0LnNc2oVc9q
+jsYGwWh/xTcbBckPA7SiNxX945sFd/F4EnH3by6TP4eLMRGBep7ujliYOXme/mV
19FIanSCDxpqiMq8mw7dh4RPAfs1cNDAYqLfisB6ENF3Ii+Yk77GzyuxlsFRwlV9
ZrmNr9MplGLVYqXgTDOSb5GRlM2l3MZ2IfB1ZIqKlpo0azFEY8/2/cDxoZckO4X8
8yuZBygRbjcMNQqHOh+NIicMb18/1Oa3AmP1IN0piJk1LRqThK2EHjjhNplTWCwI
iZQHS+le8Ue0IPWi3HTfiBCrB2EZ00NXszFfvi6+Rc6TUXuaaKbFS23v4KXXuq5E
lyxfXrn370MKPmkVvn3LYDZdBFwFgNHZUS6YZQim8WWsy8wNuBG95s7wjnNugw8X
QIVH1aFvV9oDLJfBTvRqNH1THNVyevD+r9R4h/KsDpIO9HudqyR7UgJKK9YY6NrU
hqjuet+CtFzVUkU7PBFT6+WpyjGRk49gDZLLyxULznxr2JmnieHz11Tno/QVLpeo
XojVXFCIRSZ74aarz5mpGkXC92lmEfFxqixTqLUoHaZMcJooX2fTpVD6gzLNB7pB
ObXE955wwFwcjS2VA9wlQB3T5NrJuKq89hIHTKzQsOL6ckeewTZAKmetBVoEvOKL
D0byvc2sUuyTVA55KThHV2755rifxGrqVjHAk6EPFVue0BdKzNa2v9IvkZQsugMH
/OSOd1E6UjbmjmiOrmwGM20rwgJZKB/2e+jbtL81qjpMGXM3CppLKp0IV7LdxTpb
qov+lAYVaILyTNKFsAqXGQzS77jsJRNVYdLxj17H4QOeUNWvHESGOg5v+zeLQFbe
FxP8bqjKlEO7UKmMnX3sXKYQ7lU1o2vZ2PO0DojQXiglLanL5Y5vDzanJlxihFJL
ErhcW1QNdthsXrSuaI6DSl0jztScR6ChOGGZzOJz8sjKtVuLmgmBnUQ+Q16AnpWK
lU+ntvjMfy1lEE53OrY5Q+RxdJ7U8jUELvhQZGA5SyN21I0f6FSKv/cBvM4lDS/Z
x4NQkHrxcy34yu9adOxaaPUuj10I7HRJcS96uqReOT2ZQTqajvYH9/CSPD6baRZL
n9e6/xdcMMa4V2ajiDw47+9ajO0dCQgkFZasvnijovyeyaikt/UHkjTG8LeAyH6L
2LSoqMr+fUBPZm0qNgFuq/zrTfE6OY5fHpUlT8T+u8q9KrtSVsU+5H1OuAF2fySw
+dhvKPm1MJ+StOiDOXa/qNGVPtPKewlXiHZe2rw9acfZdRSSMfZtND9yseD/mMJr
9JxzWv27B/sDqixv2hrXLzVuV8tZjJkaEPiVXT6qUiP4rioexwgih3mC3u0zMHUP
9QS1l4QrMyBWtebCptn4c+U06KLecWzmvyyJDE4yRVOVmnxGJKYGrEvD2j6x73Kx
OAHdO/nTA3IdXKLONXYBHQweVw4U4KtNEbXY9KR1nmD53FgJgyWhrfQSVqDdsAIw
BBLSJpzGEqXypb0roerTbouYacDnhKa8FvSkIy+I1na9g7dIlXuE8qNMLBsFogpA
UgRAOz60rk6GHX6bhOaJkIqbaeL0lvfAElwiftf/HHEQADCKQ3nsBXKUjv/XYsiJ
P0AvG1wRkS4SkPjhnV2jaSl/wzLx2RCvgIHtsPJSuaEUjWC2exLe2xY+nI0uRi24
1b7GnJYH+CXp/PAzzZdizPic6OKEdXhH+yle0FFf4O4vNNYEfz0dfRdrC/6N62p1
NxB58fSlTHa7RESC9RSBVgxB7cpmsLO3MqTU+Omii3i76hnI/4KxmgB1eKElYIHx
g4m8QQHN/l8S5R8sRodJFsXGQDGBogd5fcxCc8SiuAao38QDXMAZz3xUEq+qL+ka
PbxiRQJZK12T7vFQUQUUmJS3IFUjixjGH8etAEUWvc+NofqX6LRdy0hlvpsh4KGB
D3uuwKu2tFslLPD8MamC02RIrGEnuGuzt4KKnVKSMIo3Z3CCt/sSJe1+TJ8mKzft
096ll3KJiR/pN5SgQu/Tg0DnDfRsCngnMWuwL+T44kC0sjQx9JLLeDGHuX27dxo6
KgmpuCeQxl3PHynmReae8QNCDPROIQx9gKWvckONc4sj/MvX63MbC2t9PxNa2nHa
XwXPq9ZYDCkWe+bIcGJTBYubzfXxOVaYN+7iPDgrsaGu1GkB5yFZ2I0VUfukfb3A
9EjMHg8PmP66CHgWopeq/eznEFDb5D4JTfEy7ss2A9x1Mx/MM4QEZDKMJXTPP4pS
b1dt5/tCJ2jD0hq93y9I2LBzZmxO1bvDK7VUwI2irC2vYef/2IYOOd0BqQzKOLzh
EO8Fn3tOB5Ui4MNiiwtwCYd/kdW9Ap9aCj21iB1qouaMvoTug3dbh+pkilbNdTwr
Y7mDCEIsP7Nos5hokofr0yc1eZdGJ9CDc9IHUmLUCYWY2laWuOKJQ7pOWbrrZ8O+
fQFWGkedA3XRsvg0O+JWo159MKR2c0T92gUQpIvSX1gMjGJz01LIyfHHcsHY6VUP
Bp3rArN4C31N3k2ddYKBo6ZonOkgZNFOmnwaaXnQ2g8YRXPdMJG/u1U+qZKzI0xg
6+8EPYNk700cAO+Eka0r2TVEnejPAg11fu4MYWjLXLucA+PZkc5E6HrrEnykJwnO
bPrQFYMcuxyG+BY+ZwKLwFJk8aveRwhajfNDZRu+zE8uF79W3of8qYza2M84ApYS
TRzzuF6ovNpITENWRioYDmvxK4ndn7jJNIjJYqdZpi1DcPeRNHIXNJXlbHsxY/f0
tqoi8VP2SeIkHt6PdZEfABDwXV8UvQq7zy+W9/iUa4OpiohH9TOcDS+aNhMzqGrg
8bW4bQJWwaQYBfpltROxwoXTxZ6PkYmk/93mhXRa4gknxVbZbi0l8SqHJrmjEY65
jnwHT29ocy8ReHBpstj8jk57V3Dfr6ZwAYd2S1zagJi9MIFl1DR4Xx/Fn//6Ik3Z
FQjOuBU75l6IjDkCMFFXi0a1W/0rMrX6siAKYBfCPUEiBNW1yVigkpfR1MsSI72d
ID1EGTjKTr+9d1MEqAN5bH2Alkug5bHoXVu5SFg1IPQ3wRglh0brwJYaLi++Geoh
sLbFmPnj0zNhl6LfkLlYEjj/8rNmD7l3BMT2+pgM6Ai8MTn5XbjxpyH19J6vQhJd
cimpboVLp7XdIZWQxF31FaxSllD7xJHqPWUX3IzJZ8DiX2+9J10qVen46zP9l/bb
NURilxwZtNdJKHBYlVRGX7N60AtHBCtfpd4nJRcqS7nkmhboUX2xtV0YWG8//QC0
ExsCpisIHYRt73pBmSHKiVMTrb++lRS6FX8tst36wuaR6AtsGWWRA92cg4ARAAm3
u7i2G6q7emZDBuYv7Q+E+G0d1K+xHCGwdOSbEb72BzAGl4p1mvTQD+Ht0RhBvSem
pgbOe+lzHVOvbnG6RxgAE0EhJXV0Qhfx+bQNalOznL0c4buWqyv0hVmSOEizJH4c
jtMDXv7PkHIkFc9ARFbMwSbUy1aV5/PDGXdktIzqajU60VKoNdMuz8sY+MJ/mwXs
/AiXNEyBMm5jEqDsQmonT7r21t9jytrmkde5e4NEncU/w6jm9+BdwVuoJsRn8lcn
DAWX/b2b4KacWgPU7OPkURqKjmDJ2VkB5xUi8qZokdg/9vepSGNaL9WA75h6erJ8
XRLSP/2UXwlvA29AigXQPrhGY3sKv2vr2yh4gNt9othzW9J7DssCDndC/qfyaeZN
3FV1MdCqMMbFIUi1NVctjRJMPF2h2OdCYQ3J+ewn9iJA0X3YCnJ6rHSToeyS+Odk
+uAX/O8dUz5/HI33HwRozVL5Ob5NUVxWOQKATaBKKNZ9W+f8ILaKaXSATmyVPEoV
kLIZVPrHu3Y22CDk180EeR0AJU0Z7AgFDvQ72ntV+2qcTgdK3m2heoWljM+BLZOG
wazh6B42oC/xIJhoGnUznq3jAzja0DvWE5cEyDqZOgNRWvrYFVBlHL+L366RSO7g
eeGYfbTdlswY2FVSquoOF4NE4jmBVIAI8C4l119hby5aE06bciMQA58TTBhbCHQg
NjLiXkCkJPJAGsToTZfeZNZ2LLl54LkrQrhKsdNgKUzwb+OyZ7/u1A08N8tr5+8F
LIXQMufV4Z3mcQrR3T7eBKGpS0lTVoOxhTO+RTD+T6kd3mDWkARGpSD+U7mfC4tM
M89wRnnkWqm7gbyr2NcflRDTluCFqFRJnfJ0x7nyc4jcjcxbXku3wSuVKnHSRbio
QpcAb7B2gxzPXorDswB/ylSJ+dToWcmwQtPjAMo8XrGBFCASHO0LCr0IHfNgOF9C
f0uaFKJyG3uYj+RHIoJ3RgLf+xF7U6PKLIA/XpzwlbPRY9tLSVXhp0+5VZd6ev0X
+QcqbCwQeYqMjiyMp+dOgja3wexSWdsuZL62RAt7TFbOuOZfnnAuC5XAaHLSm0zy
hamgiyJEfxOt1b5PTGxkvSK083INCcOb18WOLi/uAezdk9Iywf4YWJ0cbhWeBsOH
qYFYeZ5BSmU/ZhKkf0ex7sCT/rpc1GC7oLNj6PCakpZodq3mpgkGKozQInnxO5I2
DZzevF3sfqGn9HoQhGzejrFBGBSju6fcpvQ3ZlLkpZW68+zX64xV6ohQfe/jbgfH
fk8vYxL3+Hs7Q6H/UavzENyhrzq8X2AXKMTObVxHO/4BY7JWdrFaYX7QKEfywSwB
Uuh6gCRslEUDfNTHGX/Psxv7QiWbhL1S7WfTZm15St0DC8/lafQzy6gbXeWq/4mG
AakUCSNtSUC4o15ZupNzGPGBCK6lo+uuLQTpeSQ+Ky2BZM9gkK1IzLMflisF+omx
rfAiQ8ZWT3si1PVJsXzHMXZd7LPnCeB0UiqcAd43k0RIt3eor3MaG0DjhhMOaymm
7giufvMf5L7Le0yAo6bwhePsDBWLkzSXLzOxKg7PG/80d1LGwvzqm/pSUWisIwMy
7kd8zJ3+MhHY8C1usgbGMaR2xfhR2Z3e+QgsrOwY9NWuod8oStX8TC3se2UKWIOM
3eYITP0WR1kRSo8EkVv+obc+J741JJ0dThrIy47UVIX2JrA46G8iLg5Hu6+ku537
lQt9LfV1fiUl/IsEFls5ohhO5dAAMwMbzv73r920Fr6ZurbQmzhtvg8Ig8wCmnC7
ZXxpblLjJ1L43hvxT+A+beT3vhVD2vujUI/HMISTNiWaZeYGmTRMPXqGxGOqO41X
W0mv6cm7fFX0PIm34xRa0rUbFXht6RPOC1jgo49B3GPuZb8Jf0OPWSqK1Qjm78QY
TbsYEl5iVC+uleaDIh04C/riqfh9+wi/5qR6s/lTVpGiPXDnL8cmxZhrZY/TJerb
ivE1p2TFm8QgEgiEv8yS/WO9ZFZhTj3Ojs8qz08kyNfev986oSL/+/cpFcWpxTOo
DsSXUruCrVvw50CtWy/k284i8iKA7MitFkdxnIYS19qE7FP8aDRjM1LyBMCq6IBF
85LCkU305gSfobgYxl5ujY1h/425pm2Lam97aD1gQCMUNviThtHa+SpWm6Or//tm
rbfgWr8zrGoJCMXYiWiad6UavipQwa9E+DGz7NF4xBV+WbTlIctby0uF9wOCsG+p
bCuDCCQYQEMNKWqxotlzIVbJKByeezMAamKhhuI3danqqJRPIfHSKnQnfmRNWZPy
9LELIR5BrfWgTJgEuSvTWHPspsYPKNAVWI8OSW/5eoW4V+hBMl5DRdXsaJB1prfO
8oWAncjJv/1IVaSS2lU1ZciZtyYCo+tBbl0gVltDWF7QkdcZk8pNlC8toS327CMO
rfulhibKnEMZ/cL2fo59tXD73qXdRArdJvaMChUjhyXv1D88XBqhMZhDHs7NaIpI
FKIwdpJTza6gs9/rm3xpgFdqedtHs3KlxfTiYL+q8bPftu2WbI+GyFs+5prJoVzg
C+S2wPAg+w24HaITrxSkDZHFkv0FwtwoClaIn3Du2FnrfeQ2ikzm7+K7bkflA9YT
IB5WbRASeLKisOUa95VlLhLWujQKSK2xzLrn+917sj0b2LibnkJClzz0R5J5BU5i
xKTvspWN+CLA/x981YuLrrY/rnPdfNue+kfJvq4uJwpbcU9kyN7JrMkmaI3BvU0C
emby09c7AQKCg9Rtz7Yn+oqkcKOUVa1/Nvsqh1ZgfYFmoWSek+Z+Ljh1CtQ9Z/D2
LjS3x6nhIn4uOUSXlNQ68iZpBXD7JDYK4HV5hPFN3GBTnzGJf3Q4U3MTYqeLX9cT
QxIkP3SkoYjMd7ToD5g1kBJ2hHxdO8fxOhMeGUKEDu5ty3U0Qqgxss5J5Xv9RyN2
ABeYk51772J1OlA4tDpeB8+U8M6y8JH+t5UnIuS3IA4MbNYt9iMpoAt6qQRRxZaE
fVtB1EeSrqF5bVQ83CUzqw3tz7Q2fCabyfJk/RaqobB7DUPfZCsc23w9cgsIqcJ1
PDK+QLXeBCPM2LnZpooAl+m6CXezwBBhNnGGrIu8yH6/KGlk0Mk13K+7NLAKX5eS
fFgMknFFrnlOKzwegjx/knNyMCw3Hs2/cqcCzyNLrghRT83cZ4FmkSri9pVRazKV
LLVpNuyrE1t1aKq/gT6rsS8ueD3h4f+WwxEJrMPyqFlieIpqv7tHTadHqKrplIX/
JJvukpGB8R5BToEnvs+8WzSbKWkeGKS2vS1qGeK00bxC2r3lqsZO8+gToU+Jorhh
qO56YA1y2d25ATRhPgAOpmOK4JOoaQsdV9qiEcadOR6zAYsDrZTDQVSDVflwB6pK
4UFTG8bnWWBhsly6w/IOf3a0PEdaWbNEkVAAja3QNyj8KLedFi3YswnAC177AkzL
OhmfmFnvQrVdtNJ2qB6f97b13I8jKrU8a1QE5quEsEDZgvaTGyZ1sbZhZ/YSA3KS
K0nF93970I9mz4/nL1aDM6qf64biNnHi7sHkIUYsHZrrgy1M5yvdHYVTBsFa2qU9
A9HeSdnBRLQdiASCr681JhqHfBRJz2fz6ohXQk79aKZKfOCLjsKH6sh7AqLcz1Hp
bGgRE5oClaUDgtssarPVQzIByANDcCOeHqqVf5qTEpCPlnc+oW/J1CIbuPcdfBk4
ncwuAhfcr4EFs1itRp2XI6i2v0kBvxc+MW+TxGEmcKpLAiGezvVjCYHzOzbNHKCu
riAXddY9s8m2mYyq5Lh4oa1dpndy+mqOm//OKdYu+QaabtO2Yzm4pO4/El1+Zhc/
PUcbAVf1TG7+WLbb1htTxW5vysGvXrB6dBCGHtMRoEzPabQUgDcL3OHdpsHUa1qE
cZHpIwN8NdXsN3ISo3T2d9U+S3zYIT1gdZnpdvRAuqPFfXubPTHbX8mSjZErR4OR
q4FCVIyYoBudq//kJr8DVgC/voQvSMo2k5dSst9LqVxkE0ZmeX0Ocxqzg6we3lsI
cLH9N+l31pVoC25+scYmkiGoxvUf1IUgnYZ57XxLef0NAAMXiCl3ky4xi7T0tXDv
sj4pxj6pIhcyulv2h0aytVFDgyTGWPyAgcDyMfi2nJkK7HzAukR9S/KeoyvudlBS
m5vdtRbiY5WnAdbSw+eIJI6uEnSLSM1Zic4tTGR2R9Fq5e4BhUDH9YPuEFWzhpfC
25svuZg3x0/z9oLQy/KK2ljjRyWiDFKS1+ztu/7D8JBIcuq4Na4btpoZhpikNd6/
+MTh3Q7hkAwR/Q1fIo7JlF01NEZLcY4pCJM2YlcxwttZ2sYXCxEFhx12Yc4wqv+j
SZcIfAYnV8Bh9truJ75k70i22o5uFVP6hGyJlVQazYQdtu+DhVBMj5ae0Q0psDsk
T5l45cf1M31cNwP3dzIz33L4hmQ4NuNCySF0FSJJ9R8YKAXU3sDAnUR6OgxB0Skp
M+iNxq+gwsgLNjqC+ec6FQLDAurPLBQNuyqnYfvf9VG3X4QeTxcgvpjw0hoem1vS
vbR2hol1RJRSS5CCZqxQ5eFAnGAoyKe64Eoa0QZCpPVlM/qI2Gl5H55wUeUtylCc
JCqP0Vrqpq8+SrZdSV6L4D9oD8WzWJuaBH7tf6WVTvN4c62+Z+HZ66Wc+D44x40r
QkHeNi4Pgo7uxcKFo4tY2Y8B8uVHfjj4iMtBYq+f5O2KCw4zXJAZefsrk0Y/jDbb
cwf9PC0rlMSC9cWHzdcy7jq3bTyVQPfHQIRXP/UuZXCiEPqA1+ryadPuPOYlt2Fd
mV08ZaqchO5uzxcz8hqpOHM1+3fDZiI4wvsNMyzavQQatz9e3Fj3I6MdEzl9T6gi
Wtk8tNs2TPRHj5+LrtmyHByJXjGd+9N/wYoJ+lFaRAagPzGJf8KNI78Z5AqbtCoD
1TogZqktiwNiSkZSsDnLLAqDX2K3e9wBPLxI1lnNJJyp4g4GWinW/FQt9KqC7b7Q
WeoI9L8HXDvv4nhHgpk83EApJv2fFnxZQYzGS0qABI24OEpuxDrh4O7T2KEQprKq
CZKh0ZCmnx2oFUfC2fxCN1SMoe2jYZwdAOLmL4SxN1mEsvTlicjMV2DPWiN4SKdY
2uYhCfTEIjewlUq7DWKkXJVNTHCy9MABxWpcjewi2dT6hytq+L6YiaLczK8c28Rg
EnQ/AgFCBIIiK9vuHRtuQDPLChaIEjG0BZUbctf46vAvHTAQkQl6aBAfw9pdifFX
+SpZVaKpuv7FN5NjtJCd2AklbyFHPzrb5D54h78qyPI/UvGg827d4PA2MUp6LapC
Rx920VcdlvVyTCtnvEg/K5ST0/P5M5sa6FYGSESQUJo5cNobr12pNacMU9b3IzFV
vEOroRqUFo0CrGWbfJjPTQYM0LJldm3q366koOYUbifIupp0EvTXAmOwMqQ3gxTG
5cImPSmumVbnHybOJCyF0APahqr6RYDZP1+RcLpvlprJ/f7e4lhMBk6xnF2pA+Pq
BIz1ktlTn790pTICxAyAvztcTop5bs9HUEp1b63V4VREPfGDaA35BTmH2j/WnXrI
x0ymru0TKb/Q69BlXMEVMclyMlRgXVpk2i3rmctL8p3O1F1t4+rb5OQaX/4Dx9w/
N/tB9p7ixp7l4ukr5MewSsgxYEwxu0DSVfMi2CrQ1Q9b6KTb8rFAYTfDAum8exJh
1Lzkh+ijcv59jC1FcIaQXBuEKFf5+QryrvMQLppLoiHbNpy2tG67OPoMnTGvXsEA
v8lo1/qfab86bFY75x8dDUqGoSZuGQjcFJPIcSGeWCg6C8IdfxNISvv5Vn4GrtML
n5p8A/WNkopMb1rgbD0hEFIaBeq6PRcVc9MJS2FWl+1gALKTMChATOqQt/zSTXf5
KmIubwIeQ11jzCcBn+hBROBjnC9zJjasOBgrXnhRhFRTQUka3EglWAoQzbtAIMxu
qI8eQzWMF7w/dI7rHeQvd7TAecS2wvw/1DN3TODtCblJbAKPtjFMQpf+BsKZOqto
9aV6Up0LKwz7bbzNGXRzphrhK0EJWYBEMqENMve05eALSAQY/1ou5f2g6qSR9JfV
a7BeAofJRa+iZFUNBOkPktESNEvghj+Jvru8nUJBQ+h79/Wg4NG6dorz6YCio9GX
FR/6hMY9VD/9U9QnKHLROtyuOaJ7Qt0kr8pzMdIWwI7Hp2CQjm+FIWypuXMj5Dzz
akPKikUd5cwvW2WHB1wKZUcv2fEIzZRAI0I6erAdRprWiiM2LpqCMMMKJ6+tFAqY
aZ+DzjF3SkVlD9I/tVkUZ29pORyat5wKEmVeufkwL2Qv7kJMMG6quqhPmJJfTLAz
q+i0D/qlVLkvajYFnPU4Cu5BSK3JK+jQ8+NH4etLDXVwpYK728Gbt+NjWlcxrXK5
8pUTEL2seE3RuCbx2iMVapT+GDSSznRBS6v+lC4l1W8s0bDbsKbj8PCHXwAsD0zi
JKoiVW/cO4dDLfZlYIjBhBzmuSvaUouWT3Vz2C+hwGGh0Xh4kbD2Ugbxkyuoc2hG
VTFw0jabN7YXEh6U0+qTuI132lra3NilaDM26pEgvOF+AX8IfWvBFSQJ7Ua3SAFX
/cMEjflqMnfhNiaKPJyIVDz3npWW9uPD/1Y2O1eG5Cfn8AlpGp9NkpNkga+ZRWxE
1y7o7Vy4TbjbHECl3VLgmQjqU0N1+BrRnb86f6lrBFRUF8/Udz2dc/NcLof9an6S
JlcR32RUnnOmM+4KBphgdRQRaLAgygeR5MYPhETqUO4LnsMVVoC92AsgrhiLnYtz
cENvbLkUbHzmXSJRmpZZNZgXuiLAo+nXBo+DjaMwI1JCpXn/hzyBhqQmezOYrjUg
jiBdIHqaE2WTeo1K/GwKAP4y3Ps5dnRNO/4uZpVlNsvf2O6TSrR0C6kN/zGLuLyE
zArTTWuw7+vUzET2RBHRLKC4A5IJbwlyFoUQU2+cN6kDx0nntehbc+bh++X5J2yW
qqu7Exo1gWkHDUp5XMSM0+HNphuPgPKHfqt308WKcuuFffqBpRbE+kWk71tfSFas
zmz9T7Ffv6WdtnSxNLKCYXYD3HncPtA9bOcvdMtUhvRanTtgL5e0TIMiH//tBMaO
hC6m4acN4radD6Ea+WGK+erADs5XlyYIgVe+YBparg2AXooxJL9FCp7KGzj2ea8l
cJZGsbNNe8BV41yfrr8ITLubVD9jjsj1RaWPZDMXLaZalIp5iLXrfat+GtKtsgtq
/cdASqLi2M1XPfjDMgX0ZOWsZc9VFHmKP5zoM1xJRXVW7w0UIwtMb3JZHSZwl4QI
YsqQMR3RRU2h14KvVlSc6Km5CmpDp9rGXHvVQK7aD9u8TURNsXse62dWM96/mQFW
712ctvL1DCyZItNlO/AV9uMBycifpoV/QrpcBdcdqa5tzzA6Akp0ctQnmTUWKGLK
sdFqDEbnglAZ/QJ0pc4B/O6XZ27h5fnWqPMFWdiptnGG2rb/akZySXbg/yROd4dn
2PocYg2JC9bAu6pBErDlEMkwBpgwwh+mDgT98gt2aZh0TLNfazLovACqzCJdMyf7
M2I9x9KhlqNqv9IezNOVxUsrepQ8HZsemGhUBSTf0Z1N3/UMeneDa6/yI5Q3OS+6
h0yjKeIcjm3hSThS+HEqCwWZSol85aop+EJZfJKDbl2x/yUR2AVfj+NmhHcrOAV+
jVOvxGFzkbhiGsjffuTGRTXRQgx7tlQK2vpyABOnxL9SgMyN+c2XgcvChGeQCHPv
JRpHpK7+CHsnIVhoSeE7Ig83BBdcwTqznGBgS2xGPDoOJ2yxhjXlj+HCRPbEC8Ls
XoiqopBVUyGzH4DnUN41z1qzEEtrgMnn+EDWIxLtQH6X790QuNvbw+ZEwvc6USwv
EqpKDplqCZhw7OcDacJZLFD8lMvAAsDmNJYU61yknFVGKmS57DirD4QubQNmpbTj
lYi/PSnGBMUzrzhWCLWAC+tvyhDL/Rmb4fzSpA10Pp3AJOtBvdxJSsGJxqW4U87s
mPAy6IpfLDqOtU08E+8oX5/l0S7NHILxZvz5SIJXwm+02FBS7GHt+YOgSxZ+YvrS
frhcm9LhbAoG0usRzpeLIWZR4ifKSlS+28Z5cJFOUQnH9IixWd4prF/gG1SA1rzD
`pragma protect end_protected
