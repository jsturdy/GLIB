-------------------------------------------------------------------------------
--
--  Module      : mifgen_dec.vhd
--
--  Version     : 1.1
--
--  Last Update : 2008-10-31
--
--  Project     : 8b/10b Decoder
--
--  Description : Mif File Generator for 8b/10b Decoder.  Simulating this
--                code generates an output text file in .MIF format which
--                is used to initialize the block memory for the 8b/10b
--                Decoder.  The verbose "DEBUG_OUTPUT" can be used to
--                generate complete documentation on the inputs and outputs
--                of the Decoder.
--
--  Company     : Xilinx, Inc.
--
--  DISCLAIMER OF LIABILITY
--
--                This file contains proprietary and confidential information of
--                Xilinx, Inc. ("Xilinx"), that is distributed under a license
--                from Xilinx, and may be used, copied and/or disclosed only
--                pursuant to the terms of a valid license agreement with Xilinx.
--
--                XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION
--                ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER
--                EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT
--                LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,
--                MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx
--                does not warrant that functions included in the Materials will
--                meet the requirements of Licensee, or that the operation of the
--                Materials will be uninterrupted or error-free, or that defects
--                in the Materials will be corrected.  Furthermore, Xilinx does
--                not warrant or make any representations regarding use, or the
--                results of the use, of the Materials in terms of correctness,
--                accuracy, reliability or otherwise.
--
--                Xilinx products are not designed or intended to be fail-safe,
--                or for use in any application requiring fail-safe performance,
--                such as life-support or safety devices or systems, Class III
--                medical devices, nuclear facilities, applications related to
--                the deployment of airbags, or any other applications that could
--                lead to death, personal injury or severe property or
--                environmental damage (individually and collectively, "critical
--                applications").  Customer assumes the sole risk and liability
--                of any use of Xilinx products in critical applications,
--                subject only to applicable laws and regulations governing
--                limitations on product liability.
--
--                Copyright 2000, 2001, 2002, 2003, 2004, 2005, 2008 Xilinx, Inc.
--                All rights reserved.
--
--                This disclaimer and copyright notice must be retained as part
--                of this file at all times.
--
-------------------------------------------------------------------------------
--
--  History
--
--  Date        Version   Description
--
--  10/31/2008  1.1       Initial release
--
-------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_unsigned.ALL;

USE STD.textio.ALL;

LIBRARY decode_8b10b;
USE decode_8b10b.decode_8b10b_pkg.ALL;

-------------------------------------------------------------------------------
-- Entity Declaration
-------------------------------------------------------------------------------
ENTITY mifgen_dec IS

END mifgen_dec;

-------------------------------------------------------------------------------
-- Architecture
-------------------------------------------------------------------------------
ARCHITECTURE xilinx OF mifgen_dec IS

-------------------------------------------------------------------------------
-- Constant Declarations
-------------------------------------------------------------------------------
  CONSTANT DEBUG_OUTPUT : BOOLEAN := FALSE;
  CONSTANT MYOUTPUTFILE : STRING := "dec.mif";  --output .mif file

  CONSTANT CLK_PERIOD      : TIME      := 10 ns;
  CONSTANT HALF_CLK_PERIOD : TIME      := CLK_PERIOD/2;

  CONSTANT AJWIDTH  : INTEGER := 10;
  CONSTANT HAWIDTH  : INTEGER := 8;
  CONSTANT MEMDEPTH : INTEGER := 536;

-------------------------------------------------------------------------------
-- Signal Declarations
-------------------------------------------------------------------------------
--Decoder Inputs
  SIGNAL in_din       : STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
  SIGNAL in_disp_in   : STD_LOGIC                    := '0';
  SIGNAL in_disp_in_b : STD_LOGIC                    := '1';
  SIGNAL in_sinit     : STD_LOGIC                    := '0';
  SIGNAL in_sinit_b   : STD_LOGIC                    := '0';
  SIGNAL in_ce        : STD_LOGIC                    := '1';
  SIGNAL in_ce_b      : STD_LOGIC                    := '1';
  SIGNAL clk          : STD_LOGIC                    := '0';

--Decoder Outputs
  SIGNAL out_dout     : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL out_kout     : STD_LOGIC;
  SIGNAL out_sym_disp : STD_LOGIC_VECTOR(1 DOWNTO 0);
  SIGNAL out_run_disp : STD_LOGIC;
  SIGNAL out_code_err : STD_LOGIC;
  SIGNAL out_disp_err : STD_LOGIC;
  SIGNAL out_nd       : STD_LOGIC;

--B Decoder Outputs
  SIGNAL out_dout_b     : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL out_kout_b     : STD_LOGIC;
  SIGNAL out_sym_disp_b : STD_LOGIC_VECTOR(1 DOWNTO 0);
  SIGNAL out_run_disp_b : STD_LOGIC;
  SIGNAL out_code_err_b : STD_LOGIC;
  SIGNAL out_disp_err_b : STD_LOGIC;
  SIGNAL out_nd_b       : STD_LOGIC;


--Internal Signals for Testbench
  SIGNAL stimulating : BOOLEAN := TRUE;
  SIGNAL dlay_din    : STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";


  -- compare the generated mif contents against these golden arrays
  TYPE t_golden_aj IS ARRAY (1 TO MEMDEPTH) OF STD_LOGIC_VECTOR(AJWIDTH-1
                                                                DOWNTO 0);
  TYPE t_golden_rd IS ARRAY (1 TO MEMDEPTH) OF STD_LOGIC;
  TYPE t_golden_ha IS ARRAY (1 TO MEMDEPTH) OF STD_LOGIC_VECTOR(HAWIDTH-1
                                                                DOWNTO 0);
  TYPE t_golden_k IS ARRAY (1 TO MEMDEPTH) OF STD_LOGIC;

  SIGNAL golden_aj : t_golden_aj := (
    "1001110100",
    "0111010100",
    "1011010100",
    "1100011011",
    "1101010100",
    "1010011011",
    "0110011011",
    "1110001011",
    "1110010100",
    "1001011011",
    "0101011011",
    "1101001011",
    "0011011011",
    "1011001011",
    "0111001011",
    "0101110100",
    "0110110100",
    "1000111011",
    "0100111011",
    "1100101011",
    "0010111011",
    "1010101011",
    "0110101011",
    "1110100100",
    "1100110100",
    "1001101011",
    "0101101011",
    "1101100100",
    "0011101011",
    "1011100100",
    "0111100100",
    "1010110100",
    "1001111001",
    "0111011001",
    "1011011001",
    "1100011001",
    "1101011001",
    "1010011001",
    "0110011001",
    "1110001001",
    "1110011001",
    "1001011001",
    "0101011001",
    "1101001001",
    "0011011001",
    "1011001001",
    "0111001001",
    "0101111001",
    "0110111001",
    "1000111001",
    "0100111001",
    "1100101001",
    "0010111001",
    "1010101001",
    "0110101001",
    "1110101001",
    "1100111001",
    "1001101001",
    "0101101001",
    "1101101001",
    "0011101001",
    "1011101001",
    "0111101001",
    "1010111001",
    "1001110101",
    "0111010101",
    "1011010101",
    "1100010101",
    "1101010101",
    "1010010101",
    "0110010101",
    "1110000101",
    "1110010101",
    "1001010101",
    "0101010101",
    "1101000101",
    "0011010101",
    "1011000101",
    "0111000101",
    "0101110101",
    "0110110101",
    "1000110101",
    "0100110101",
    "1100100101",
    "0010110101",
    "1010100101",
    "0110100101",
    "1110100101",
    "1100110101",
    "1001100101",
    "0101100101",
    "1101100101",
    "0011100101",
    "1011100101",
    "0111100101",
    "1010110101",
    "1001110011",
    "0111010011",
    "1011010011",
    "1100011100",
    "1101010011",
    "1010011100",
    "0110011100",
    "1110001100",
    "1110010011",
    "1001011100",
    "0101011100",
    "1101001100",
    "0011011100",
    "1011001100",
    "0111001100",
    "0101110011",
    "0110110011",
    "1000111100",
    "0100111100",
    "1100101100",
    "0010111100",
    "1010101100",
    "0110101100",
    "1110100011",
    "1100110011",
    "1001101100",
    "0101101100",
    "1101100011",
    "0011101100",
    "1011100011",
    "0111100011",
    "1010110011",
    "1001110010",
    "0111010010",
    "1011010010",
    "1100011101",
    "1101010010",
    "1010011101",
    "0110011101",
    "1110001101",
    "1110010010",
    "1001011101",
    "0101011101",
    "1101001101",
    "0011011101",
    "1011001101",
    "0111001101",
    "0101110010",
    "0110110010",
    "1000111101",
    "0100111101",
    "1100101101",
    "0010111101",
    "1010101101",
    "0110101101",
    "1110100010",
    "1100110010",
    "1001101101",
    "0101101101",
    "1101100010",
    "0011101101",
    "1011100010",
    "0111100010",
    "1010110010",
    "1001111010",
    "0111011010",
    "1011011010",
    "1100011010",
    "1101011010",
    "1010011010",
    "0110011010",
    "1110001010",
    "1110011010",
    "1001011010",
    "0101011010",
    "1101001010",
    "0011011010",
    "1011001010",
    "0111001010",
    "0101111010",
    "0110111010",
    "1000111010",
    "0100111010",
    "1100101010",
    "0010111010",
    "1010101010",
    "0110101010",
    "1110101010",
    "1100111010",
    "1001101010",
    "0101101010",
    "1101101010",
    "0011101010",
    "1011101010",
    "0111101010",
    "1010111010",
    "1001110110",
    "0111010110",
    "1011010110",
    "1100010110",
    "1101010110",
    "1010010110",
    "0110010110",
    "1110000110",
    "1110010110",
    "1001010110",
    "0101010110",
    "1101000110",
    "0011010110",
    "1011000110",
    "0111000110",
    "0101110110",
    "0110110110",
    "1000110110",
    "0100110110",
    "1100100110",
    "0010110110",
    "1010100110",
    "0110100110",
    "1110100110",
    "1100110110",
    "1001100110",
    "0101100110",
    "1101100110",
    "0011100110",
    "1011100110",
    "0111100110",
    "1010110110",
    "1001110001",
    "0111010001",
    "1011010001",
    "1100011110",
    "1101010001",
    "1010011110",
    "0110011110",
    "1110001110",
    "1110010001",
    "1001011110",
    "0101011110",
    "1101001110",
    "0011011110",
    "1011001110",
    "0111001110",
    "0101110001",
    "0110110001",
    "1000110111",
    "0100110111",
    "1100101110",
    "0010110111",
    "1010101110",
    "0110101110",
    "1110100001",
    "1100110001",
    "1001101110",
    "0101101110",
    "1101100001",
    "0011101110",
    "1011100001",
    "0111100001",
    "1010110001",
    "0011110100",
    "0011111001",
    "0011110101",
    "0011110011",
    "0011110010",
    "0011111010",
    "0011110110",
    "0011111000",
    "1110101000",
    "1101101000",
    "1011101000",
    "0111101000",
    "0110001011",
    "1000101011",
    "0100101011",
    "1100010100",
    "0010101011",
    "1010010100",
    "0110010100",
    "0001110100",
    "0001101011",
    "1001010100",
    "0101010100",
    "1101000100",
    "0011010100",
    "1011000100",
    "0111000100",
    "1010001011",
    "1001001011",
    "1000110100",
    "0100110100",
    "1100100100",
    "0010110100",
    "1010100100",
    "0110100100",
    "0001011011",
    "0011001011",
    "1001100100",
    "0101100100",
    "0010011011",
    "0011100100",
    "0100011011",
    "1000011011",
    "0101001011",
    "0110001001",
    "1000101001",
    "0100101001",
    "1100011001",
    "0010101001",
    "1010011001",
    "0110011001",
    "0001111001",
    "0001101001",
    "1001011001",
    "0101011001",
    "1101001001",
    "0011011001",
    "1011001001",
    "0111001001",
    "1010001001",
    "1001001001",
    "1000111001",
    "0100111001",
    "1100101001",
    "0010111001",
    "1010101001",
    "0110101001",
    "0001011001",
    "0011001001",
    "1001101001",
    "0101101001",
    "0010011001",
    "0011101001",
    "0100011001",
    "1000011001",
    "0101001001",
    "0110000101",
    "1000100101",
    "0100100101",
    "1100010101",
    "0010100101",
    "1010010101",
    "0110010101",
    "0001110101",
    "0001100101",
    "1001010101",
    "0101010101",
    "1101000101",
    "0011010101",
    "1011000101",
    "0111000101",
    "1010000101",
    "1001000101",
    "1000110101",
    "0100110101",
    "1100100101",
    "0010110101",
    "1010100101",
    "0110100101",
    "0001010101",
    "0011000101",
    "1001100101",
    "0101100101",
    "0010010101",
    "0011100101",
    "0100010101",
    "1000010101",
    "0101000101",
    "0110001100",
    "1000101100",
    "0100101100",
    "1100010011",
    "0010101100",
    "1010010011",
    "0110010011",
    "0001110011",
    "0001101100",
    "1001010011",
    "0101010011",
    "1101000011",
    "0011010011",
    "1011000011",
    "0111000011",
    "1010001100",
    "1001001100",
    "1000110011",
    "0100110011",
    "1100100011",
    "0010110011",
    "1010100011",
    "0110100011",
    "0001011100",
    "0011001100",
    "1001100011",
    "0101100011",
    "0010011100",
    "0011100011",
    "0100011100",
    "1000011100",
    "0101001100",
    "0110001101",
    "1000101101",
    "0100101101",
    "1100010010",
    "0010101101",
    "1010010010",
    "0110010010",
    "0001110010",
    "0001101101",
    "1001010010",
    "0101010010",
    "1101000010",
    "0011010010",
    "1011000010",
    "0111000010",
    "1010001101",
    "1001001101",
    "1000110010",
    "0100110010",
    "1100100010",
    "0010110010",
    "1010100010",
    "0110100010",
    "0001011101",
    "0011001101",
    "1001100010",
    "0101100010",
    "0010011101",
    "0011100010",
    "0100011101",
    "1000011101",
    "0101001101",
    "0110001010",
    "1000101010",
    "0100101010",
    "1100011010",
    "0010101010",
    "1010011010",
    "0110011010",
    "0001111010",
    "0001101010",
    "1001011010",
    "0101011010",
    "1101001010",
    "0011011010",
    "1011001010",
    "0111001010",
    "1010001010",
    "1001001010",
    "1000111010",
    "0100111010",
    "1100101010",
    "0010111010",
    "1010101010",
    "0110101010",
    "0001011010",
    "0011001010",
    "1001101010",
    "0101101010",
    "0010011010",
    "0011101010",
    "0100011010",
    "1000011010",
    "0101001010",
    "0110000110",
    "1000100110",
    "0100100110",
    "1100010110",
    "0010100110",
    "1010010110",
    "0110010110",
    "0001110110",
    "0001100110",
    "1001010110",
    "0101010110",
    "1101000110",
    "0011010110",
    "1011000110",
    "0111000110",
    "1010000110",
    "1001000110",
    "1000110110",
    "0100110110",
    "1100100110",
    "0010110110",
    "1010100110",
    "0110100110",
    "0001010110",
    "0011000110",
    "1001100110",
    "0101100110",
    "0010010110",
    "0011100110",
    "0100010110",
    "1000010110",
    "0101000110",
    "0110001110",
    "1000101110",
    "0100101110",
    "1100010001",
    "0010101110",
    "1010010001",
    "0110010001",
    "0001110001",
    "0001101110",
    "1001010001",
    "0101010001",
    "1101001000",
    "0011010001",
    "1011001000",
    "0111001000",
    "1010001110",
    "1001001110",
    "1000110001",
    "0100110001",
    "1100100001",
    "0010110001",
    "1010100001",
    "0110100001",
    "0001011110",
    "0011001110",
    "1001100001",
    "0101100001",
    "0010011110",
    "0011100001",
    "0100011110",
    "1000011110",
    "0101001110",
    "1100001011",
    "1100000110",
    "1100001010",
    "1100001100",
    "1100001101",
    "1100000101",
    "1100001001",
    "1100000111",
    "0001010111",
    "0010010111",
    "0100010111",
    "1000010111"
    );

  SIGNAL golden_ha : t_golden_ha := (
    "00000000",
    "00000001",
    "00000010",
    "00000011",
    "00000100",
    "00000101",
    "00000110",
    "00000111",
    "00001000",
    "00001001",
    "00001010",
    "00001011",
    "00001100",
    "00001101",
    "00001110",
    "00001111",
    "00010000",
    "00010001",
    "00010010",
    "00010011",
    "00010100",
    "00010101",
    "00010110",
    "00010111",
    "00011000",
    "00011001",
    "00011010",
    "00011011",
    "00011100",
    "00011101",
    "00011110",
    "00011111",
    "00100000",
    "00100001",
    "00100010",
    "00100011",
    "00100100",
    "00100101",
    "00100110",
    "00100111",
    "00101000",
    "00101001",
    "00101010",
    "00101011",
    "00101100",
    "00101101",
    "00101110",
    "00101111",
    "00110000",
    "00110001",
    "00110010",
    "00110011",
    "00110100",
    "00110101",
    "00110110",
    "00110111",
    "00111000",
    "00111001",
    "00111010",
    "00111011",
    "00111100",
    "00111101",
    "00111110",
    "00111111",
    "01000000",
    "01000001",
    "01000010",
    "01000011",
    "01000100",
    "01000101",
    "01000110",
    "01000111",
    "01001000",
    "01001001",
    "01001010",
    "01001011",
    "01001100",
    "01001101",
    "01001110",
    "01001111",
    "01010000",
    "01010001",
    "01010010",
    "01010011",
    "01010100",
    "01010101",
    "01010110",
    "01010111",
    "01011000",
    "01011001",
    "01011010",
    "01011011",
    "01011100",
    "01011101",
    "01011110",
    "01011111",
    "01100000",
    "01100001",
    "01100010",
    "01100011",
    "01100100",
    "01100101",
    "01100110",
    "01100111",
    "01101000",
    "01101001",
    "01101010",
    "01101011",
    "01101100",
    "01101101",
    "01101110",
    "01101111",
    "01110000",
    "01110001",
    "01110010",
    "01110011",
    "01110100",
    "01110101",
    "01110110",
    "01110111",
    "01111000",
    "01111001",
    "01111010",
    "01111011",
    "01111100",
    "01111101",
    "01111110",
    "01111111",
    "10000000",
    "10000001",
    "10000010",
    "10000011",
    "10000100",
    "10000101",
    "10000110",
    "10000111",
    "10001000",
    "10001001",
    "10001010",
    "10001011",
    "10001100",
    "10001101",
    "10001110",
    "10001111",
    "10010000",
    "10010001",
    "10010010",
    "10010011",
    "10010100",
    "10010101",
    "10010110",
    "10010111",
    "10011000",
    "10011001",
    "10011010",
    "10011011",
    "10011100",
    "10011101",
    "10011110",
    "10011111",
    "10100000",
    "10100001",
    "10100010",
    "10100011",
    "10100100",
    "10100101",
    "10100110",
    "10100111",
    "10101000",
    "10101001",
    "10101010",
    "10101011",
    "10101100",
    "10101101",
    "10101110",
    "10101111",
    "10110000",
    "10110001",
    "10110010",
    "10110011",
    "10110100",
    "10110101",
    "10110110",
    "10110111",
    "10111000",
    "10111001",
    "10111010",
    "10111011",
    "10111100",
    "10111101",
    "10111110",
    "10111111",
    "11000000",
    "11000001",
    "11000010",
    "11000011",
    "11000100",
    "11000101",
    "11000110",
    "11000111",
    "11001000",
    "11001001",
    "11001010",
    "11001011",
    "11001100",
    "11001101",
    "11001110",
    "11001111",
    "11010000",
    "11010001",
    "11010010",
    "11010011",
    "11010100",
    "11010101",
    "11010110",
    "11010111",
    "11011000",
    "11011001",
    "11011010",
    "11011011",
    "11011100",
    "11011101",
    "11011110",
    "11011111",
    "11100000",
    "11100001",
    "11100010",
    "11100011",
    "11100100",
    "11100101",
    "11100110",
    "11100111",
    "11101000",
    "11101001",
    "11101010",
    "11101011",
    "11101100",
    "11101101",
    "11101110",
    "11101111",
    "11110000",
    "11110001",
    "11110010",
    "11110011",
    "11110100",
    "11110101",
    "11110110",
    "11110111",
    "11111000",
    "11111001",
    "11111010",
    "11111011",
    "11111100",
    "11111101",
    "11111110",
    "11111111",
    "00011100",
    "00111100",
    "01011100",
    "01111100",
    "10011100",
    "10111100",
    "11011100",
    "11111100",
    "11110111",
    "11111011",
    "11111101",
    "11111110",
    "00000000",
    "00000001",
    "00000010",
    "00000011",
    "00000100",
    "00000101",
    "00000110",
    "00000111",
    "00001000",
    "00001001",
    "00001010",
    "00001011",
    "00001100",
    "00001101",
    "00001110",
    "00001111",
    "00010000",
    "00010001",
    "00010010",
    "00010011",
    "00010100",
    "00010101",
    "00010110",
    "00010111",
    "00011000",
    "00011001",
    "00011010",
    "00011011",
    "00011100",
    "00011101",
    "00011110",
    "00011111",
    "00100000",
    "00100001",
    "00100010",
    "00100011",
    "00100100",
    "00100101",
    "00100110",
    "00100111",
    "00101000",
    "00101001",
    "00101010",
    "00101011",
    "00101100",
    "00101101",
    "00101110",
    "00101111",
    "00110000",
    "00110001",
    "00110010",
    "00110011",
    "00110100",
    "00110101",
    "00110110",
    "00110111",
    "00111000",
    "00111001",
    "00111010",
    "00111011",
    "00111100",
    "00111101",
    "00111110",
    "00111111",
    "01000000",
    "01000001",
    "01000010",
    "01000011",
    "01000100",
    "01000101",
    "01000110",
    "01000111",
    "01001000",
    "01001001",
    "01001010",
    "01001011",
    "01001100",
    "01001101",
    "01001110",
    "01001111",
    "01010000",
    "01010001",
    "01010010",
    "01010011",
    "01010100",
    "01010101",
    "01010110",
    "01010111",
    "01011000",
    "01011001",
    "01011010",
    "01011011",
    "01011100",
    "01011101",
    "01011110",
    "01011111",
    "01100000",
    "01100001",
    "01100010",
    "01100011",
    "01100100",
    "01100101",
    "01100110",
    "01100111",
    "01101000",
    "01101001",
    "01101010",
    "01101011",
    "01101100",
    "01101101",
    "01101110",
    "01101111",
    "01110000",
    "01110001",
    "01110010",
    "01110011",
    "01110100",
    "01110101",
    "01110110",
    "01110111",
    "01111000",
    "01111001",
    "01111010",
    "01111011",
    "01111100",
    "01111101",
    "01111110",
    "01111111",
    "10000000",
    "10000001",
    "10000010",
    "10000011",
    "10000100",
    "10000101",
    "10000110",
    "10000111",
    "10001000",
    "10001001",
    "10001010",
    "10001011",
    "10001100",
    "10001101",
    "10001110",
    "10001111",
    "10010000",
    "10010001",
    "10010010",
    "10010011",
    "10010100",
    "10010101",
    "10010110",
    "10010111",
    "10011000",
    "10011001",
    "10011010",
    "10011011",
    "10011100",
    "10011101",
    "10011110",
    "10011111",
    "10100000",
    "10100001",
    "10100010",
    "10100011",
    "10100100",
    "10100101",
    "10100110",
    "10100111",
    "10101000",
    "10101001",
    "10101010",
    "10101011",
    "10101100",
    "10101101",
    "10101110",
    "10101111",
    "10110000",
    "10110001",
    "10110010",
    "10110011",
    "10110100",
    "10110101",
    "10110110",
    "10110111",
    "10111000",
    "10111001",
    "10111010",
    "10111011",
    "10111100",
    "10111101",
    "10111110",
    "10111111",
    "11000000",
    "11000001",
    "11000010",
    "11000011",
    "11000100",
    "11000101",
    "11000110",
    "11000111",
    "11001000",
    "11001001",
    "11001010",
    "11001011",
    "11001100",
    "11001101",
    "11001110",
    "11001111",
    "11010000",
    "11010001",
    "11010010",
    "11010011",
    "11010100",
    "11010101",
    "11010110",
    "11010111",
    "11011000",
    "11011001",
    "11011010",
    "11011011",
    "11011100",
    "11011101",
    "11011110",
    "11011111",
    "11100000",
    "11100001",
    "11100010",
    "11100011",
    "11100100",
    "11100101",
    "11100110",
    "11100111",
    "11101000",
    "11101001",
    "11101010",
    "11101011",
    "11101100",
    "11101101",
    "11101110",
    "11101111",
    "11110000",
    "11110001",
    "11110010",
    "11110011",
    "11110100",
    "11110101",
    "11110110",
    "11110111",
    "11111000",
    "11111001",
    "11111010",
    "11111011",
    "11111100",
    "11111101",
    "11111110",
    "11111111",
    "00011100",
    "00111100",
    "01011100",
    "01111100",
    "10011100",
    "10111100",
    "11011100",
    "11111100",
    "11110111",
    "11111011",
    "11111101",
    "11111110"
    );

  SIGNAL golden_rd : t_golden_rd := (
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1'
    );

  SIGNAL golden_k : t_golden_k := (
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1',
    '1'
    );

-------------------------------------------------------------------------------
--Function Declarations
-------------------------------------------------------------------------------

  -- convert 4-bit slv to 1-char hex
  FUNCTION std_logic_vector4_2_hex(v : STD_LOGIC_VECTOR(3 DOWNTO 0))
    RETURN CHARACTER IS
    VARIABLE str                     : CHARACTER;
  BEGIN
    CASE v IS
      WHEN "0000" => str := '0';
      WHEN "0001" => str := '1';
      WHEN "0010" => str := '2';
      WHEN "0011" => str := '3';
      WHEN "0100" => str := '4';
      WHEN "0101" => str := '5';
      WHEN "0110" => str := '6';
      WHEN "0111" => str := '7';
      WHEN "1000" => str := '8';
      WHEN "1001" => str := '9';
      WHEN "1010" => str := 'A';
      WHEN "1011" => str := 'B';
      WHEN "1100" => str := 'C';
      WHEN "1101" => str := 'D';
      WHEN "1110" => str := 'E';
      WHEN "1111" => str := 'F';
      WHEN "00U0" => str := '0';
      WHEN "00U1" => str := '1';
      WHEN OTHERS => str := 'x';
    END CASE;

    RETURN str;
  END std_logic_vector4_2_hex;

  -- convert 8-bit slv to 2-char hex string
  FUNCTION std_logic_vector8_2_hex(v : STD_LOGIC_VECTOR(7 DOWNTO 0))
    RETURN STRING IS
    VARIABLE str                     : STRING(1 TO 2);
  BEGIN
    str := std_logic_vector4_2_hex(v(7 DOWNTO 4)) &
           std_logic_vector4_2_hex(v(3 DOWNTO 0));
    RETURN str;
  END std_logic_vector8_2_hex;

  -- convert 10-bit slv to 3-char hex string
  FUNCTION std_logic_vector10_2_hex(v : STD_LOGIC_VECTOR(9 DOWNTO 0))
    RETURN STRING IS
    VARIABLE str                      : STRING(1 TO 3);
  BEGIN
    str := std_logic_vector4_2_hex("00" & v(9 DOWNTO 8)) &
           std_logic_vector4_2_hex(v(7 DOWNTO 4)) &
           std_logic_vector4_2_hex(v(3 DOWNTO 0));
    RETURN str;
  END std_logic_vector10_2_hex;

  -- search for value to be decoded; return its index
  FUNCTION find_aj_index(inaj : t_golden_aj;
                         findval : STD_LOGIC_VECTOR(AJWIDTH-1 DOWNTO 0))
    RETURN INTEGER IS
    VARIABLE tmp : INTEGER := 0;
  BEGIN
    FOR i IN MEMDEPTH DOWNTO 1 LOOP
      IF (inaj(i) = findval) THEN
        tmp := i;
      END IF;
    END LOOP;
    RETURN tmp;
  END FUNCTION;

  -- search for value to be decoded; return its index
  FUNCTION find_aj_index2(inaj : t_golden_aj;
                          findval : STD_LOGIC_VECTOR(AJWIDTH-1 DOWNTO 0))
    RETURN INTEGER IS
    VARIABLE tmp : INTEGER := 0;
  BEGIN
    FOR i IN 1 TO MEMDEPTH LOOP
      IF (inaj(i) = findval) THEN
        tmp := i;
      END IF;
    END LOOP;
    RETURN tmp;
  END FUNCTION;

  -- verify validity of decoded byte
  FUNCTION check_valid(golden_aj : t_golden_aj;
                       golden_rd : t_golden_rd;
                       golden_ha : t_golden_ha;
                       golden_k  : t_golden_k;
                       myaj : STD_LOGIC_VECTOR(AJWIDTH-1 DOWNTO 0);
                       myrd : STD_LOGIC;
                       myha : STD_LOGIC_VECTOR(HAWIDTH-1 DOWNTO 0);
                       myk  : STD_LOGIC)
    RETURN BOOLEAN IS
    VARIABLE tmpidx  : INTEGER;
    VARIABLE tmpidx2 : INTEGER;
    VARIABLE retval  : BOOLEAN := TRUE;
  BEGIN
    --Look up the value to be decoded     (it could occur twice)
    tmpidx  := find_aj_index(golden_aj, myaj);
    tmpidx2 := find_aj_index2(golden_aj, myaj);

    --Was it found?
    IF (tmpidx > 0) THEN
      --Report on current test
      IF (myk='1') THEN
        IF (myrd='1') THEN
          ASSERT FALSE REPORT "Verifying Valid Code...HA=" &
            std_logic_vector8_2_hex(myha) & " aj=" &
            std_logic_vector10_2_hex(myaj) & " K=1 RD=1" SEVERITY NOTE;
        ELSE
          ASSERT FALSE REPORT "Verifying Valid Code...HA=" &
            std_logic_vector8_2_hex(myha) & " aj=" &
            std_logic_vector10_2_hex(myaj) & " K=1 RD=0" SEVERITY NOTE;
        END IF;
      ELSE
        IF (myrd='1') THEN
          ASSERT FALSE REPORT "Verifying Valid Code...HA=" &
            std_logic_vector8_2_hex(myha) & " aj=" &
            std_logic_vector10_2_hex(myaj) & " K=0 RD=1" SEVERITY NOTE;
        ELSE
          ASSERT FALSE REPORT "Verifying Valid Code...HA=" &
            std_logic_vector8_2_hex(myha) & " aj=" &
            std_logic_vector10_2_hex(myaj) & " K=0 RD=0" SEVERITY NOTE;
        END IF;
      END IF;


      --Check that the code has been correctly decoded
      IF (golden_ha(tmpidx) /= myha) THEN
        ASSERT FALSE REPORT " ***Decoding Error_a1 myHA=" &
          std_logic_vector8_2_hex(myha) & " gHA=" &
          std_logic_vector8_2_hex(golden_ha(tmpidx)) SEVERITY WARNING;
        retval := FALSE;
      END IF;

      IF (golden_ha(tmpidx2) /= myha) THEN
        ASSERT FALSE REPORT " ***Decoding Error_a2 myHA=" &
          std_logic_vector8_2_hex(myha) & " gHA=" &
          std_logic_vector8_2_hex(golden_ha(tmpidx2))  SEVERITY WARNING;
        retval := FALSE;
      END IF;

      --Check that it's properly identified the K code status
      IF (golden_k(tmpidx) /= myk) THEN
        ASSERT FALSE REPORT " ***K Code Error_a1" SEVERITY WARNING;
        retval := FALSE;
      END IF;

      IF (golden_k(tmpidx2) /= myk) THEN
        ASSERT FALSE REPORT " ***K Code Error_a2" SEVERITY WARNING;
        retval := FALSE;
      END IF;

      -------------------------------------------------------------------------
      --  ** Commenting out the Disparity check for mif file generation **
      --  It is irrelevant to check the running disparity when we are forcing
      --  the disp_in pin throughout the stimulus to generate the complete
      --  decoding table for the mif file.
      -------------------------------------------------------------------------
      --  --Check that it's the right code in this disparity context
      --IF (tmpidx/=tmpidx2) THEN
      --  --We have two instances of this 10-bit code, which means that it must be
      --  -- the same for both running disparities (therefore it is okay)
      --ELSE
      --  --The code is only valid for one disparity case, so check it.
      --  IF (golden_rd(tmpidx) /= myrd) THEN
      --    ASSERT false REPORT " Run Disparity Error" SEVERITY warning;
      --    retval := false;
      --  END IF;
      --END IF;
      -------------------------------------------------------------------------

    ELSE --tmpidx = 0
      --10-bit code was not found in the valid code list
      --assert false report "CODE NOT FOUND... aj=" &
      --std_logic_vector10_2_hex(myaj) severity note;
      retval := FALSE;
    END IF;

    RETURN retval;
  END FUNCTION;

-------------------------------------------------------------------------------
-- BEGIN ARCHITECTURE
-------------------------------------------------------------------------------
BEGIN

-------------------------------------------------------------------------------
--Object Instantiation
-------------------------------------------------------------------------------
  decmodel : ENTITY decode_8b10b.decode_8b10b_lut
    GENERIC MAP(
      C_HAS_BPORTS     => 1,              -- 0 one decoder, 1 two decoders
      C_HAS_DISP_IN    => 1,              -- 1 if DISP_IN port present
      C_HAS_DISP_IN_B  => 1,              -- 1 if DISP_IN_B port present
      C_HAS_DISP_ERR   => 1,              -- 1 if DISP_ERR port present
      C_HAS_DISP_ERR_B => 1,              -- 1 if DISP_ERR_B port present
      C_HAS_CODE_ERR   => 1,              -- 1 if CODE_ERR port present
      C_HAS_CODE_ERR_B => 1,              -- 1 if CODE_ERR_B port present
      C_HAS_RUN_DISP   => 1,              -- 1 if RUN_DISP port present
      C_HAS_RUN_DISP_B => 1,              -- 1 if RUN_DISP_B port present
      C_HAS_SYM_DISP   => 1,              -- 1 if SYM_DISP port present
      C_HAS_SYM_DISP_B => 1,              -- 1 if SYM_DISP_B port present
      C_HAS_ND         => 1,              -- 1 if ND port present
      C_HAS_ND_B       => 1,              -- 1 if ND_B port present

      -- DOUT val when SINIT active
      C_SINIT_DOUT       => "00100011",   -- DOUT value when SINIT active
      C_SINIT_KOUT       => 0,            -- KOUT value when SINIT active
      C_SINIT_RUN_DISP   => 0,            -- Init value of RUN_DISP (0=neg,1=pos)
      C_SINIT_DOUT_B     => "00100011",   -- DOUT_B value when SINITT_B active
      C_SINIT_KOUT_B     => 0,            -- KOUT_B value when SINIT_B active
      C_SINIT_RUN_DISP_B => 0             -- Init value of RUN_DISP_B (0=neg,1=pos)
      )
    PORT MAP(
      --Mandatory Decoder Pins
      DIN   => in_din,                    -- Data input (10-bit encoded symbol)
      CLK   => clk,                       -- Clock input
      DOUT  => out_dout,                  -- Decoded byte
      KOUT  => out_kout,                  -- Command symbol indicator

      --Optional Decoder Pins
      CE         => in_ce,                -- Clock Enable
      CE_B       => in_ce_b,              -- Clock Enable B
      DIN_B      => in_din,               -- Data input B (10-bit encoded symbol)
      DISP_IN    => in_disp_in,           -- Running disp input (0=neg,1=pos)
      DISP_IN_B  => in_disp_in_b,         -- Running disp B input (0=neg,1=pos)
      SINIT      => in_sinit,             -- Sync init for decoder
      SINIT_B    => in_sinit_b,           -- Sync init for decoder B
      CLK_B      => clk,                  -- Clock input B
      DOUT_B     => out_dout_b,           -- Decoded byte B
      KOUT_B     => out_kout_b,           -- Command symbol indicator B
      CODE_ERR   => out_code_err,         -- Indicates not valid code
      CODE_ERR_B => out_code_err_b,       -- Indicates not valid code B
      SYM_DISP   => out_sym_disp,         -- 2-bit symbol disparity
      SYM_DISP_B => out_sym_disp_b,       -- 2-bit symbol disparity B
      RUN_DISP   => out_run_disp,         -- Tracks running disp
      RUN_DISP_B => out_run_disp_b,       -- Tracks running disp B
      DISP_ERR   => out_disp_err,         -- Active if disp rules violated
      DISP_ERR_B => out_disp_err_b,       -- Active if disp rules violated B
      ND         => out_nd,               -- New Data
      ND_B       => out_nd_b              -- New Data B
      );


  --Clock stimulation
  stimulate_clk : PROCESS
  BEGIN
    clk   <= '0';
    WHILE stimulating LOOP
      WAIT FOR HALF_CLK_PERIOD;
      clk <= NOT clk;
    END LOOP;

    --pulse the clock a few more times before exiting, to insure that all
    -- delayed signals get through.
    WAIT FOR HALF_CLK_PERIOD;
    clk <= NOT clk;
    WAIT FOR HALF_CLK_PERIOD;
    clk <= NOT clk;
    WAIT FOR HALF_CLK_PERIOD;
    clk <= NOT clk;

    --suspend clock stimulation process at exit
    WAIT;
  END PROCESS stimulate_clk;


  -- stimulate decoder data input with all possible code points
  -- store generated outputs to .mif file
  -- compare result to the golden arrays
  generate_mif_dec : PROCESS (clk)
    --for file io
    VARIABLE decM         : LINE;
    FILE decmiffile       : TEXT OPEN WRITE_MODE IS MYOUTPUTFILE;
    VARIABLE decout       : STD_LOGIC_VECTOR(13 DOWNTO 0) := "00000000000000";
    VARIABLE first_pass   : BOOLEAN                       := TRUE;
    VARIABLE any_err      : STD_LOGIC;
    VARIABLE any_err_b    : STD_LOGIC;
    VARIABLE new_sym_disp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    VARIABLE test_aj      : STD_LOGIC_VECTOR(9 DOWNTO 0);
    VARIABLE specmatcha   : BOOLEAN;
    VARIABLE specmatchb   : BOOLEAN;

  BEGIN
    IF (clk'event AND clk = '1') THEN

      --for debug output only
      dlay_din <= in_din;

      --check to see if we've reached the end yet
      IF (in_din = "1111111111") THEN
        in_ce <= '0';                   --stop the decoder
        stimulating <= FALSE;           --stop stimulating clock
      END IF;

      in_din <= in_din + 1;

      any_err   := out_code_err OR out_disp_err;
      any_err_b := out_code_err_b OR out_disp_err_b;
      decout    := out_sym_disp_b(1) & out_sym_disp_b(0) & out_sym_disp(1) &
                   out_sym_disp(0) & out_code_err & out_kout & out_dout;

      --Do a sanity check - cross-check results against valid code table from
      --IEEE spec (golden arrays)
      FOR t IN 0 TO 9 LOOP
        test_aj(t) := dlay_din(9-t);
      END LOOP;
      specmatcha := check_valid(golden_aj, golden_rd, golden_ha, golden_k,
                                test_aj, '0', out_dout, out_kout);
      specmatchb := check_valid(golden_aj, golden_rd, golden_ha, golden_k,
                                test_aj, '1', out_dout_b, out_kout_b);

      IF out_nd = '1' THEN
        --for debug output only
        IF (DEBUG_OUTPUT) THEN
          IF (first_pass) THEN
            WRITE(decM, STRING'("DIN(binja) DIN(int) | SYM_DISP CODE_ERR KOUT "));
            WRITE(decM, STRING'("DOUT(bin) DOUT(int) DISP_ERR ANY_ERR | "));
            WRITE(decM, STRING'("SYM_DISP_B CODE_ERR_B KOUT_B DOUT_B(bin) "));
            WRITE(decM, STRING'("DOUT_B(int) DISP_ERR_B ANY_ERR_B | "));
            WRITE(decM, STRING'("NEW_SYM_DISP"));
            WRITELINE(decmiffile, decM);
            first_pass := FALSE;
          END IF;

          --Inputs
          WRITE(decM, BIT_VECTOR'(TO_BITVECTOR(dlay_din)));
          WRITE(decM, ' ');
          WRITE(decM, CONV_INTEGER(dlay_din), justified => RIGHT, field => 8);

          --A Outputs
          WRITE(decM, STRING'("         "));
          WRITE(decM, BIT_VECTOR'(TO_BITVECTOR(out_sym_disp)));
          WRITE(decM, STRING'("        "));
          WRITE(decM, BIT'(TO_BIT(out_code_err)));
          WRITE(decM, STRING'("    "));
          WRITE(decM, BIT'(TO_BIT(out_kout)));
          WRITE(decM, ' ');
          WRITE(decM, BIT_VECTOR'(TO_BITVECTOR(out_dout)));
          WRITE(decM, ' ');
          WRITE(decM, CONV_INTEGER(out_dout), justified => RIGHT, field => 8);
          WRITE(decM, STRING'("          "));
          WRITE(decM, BIT'(TO_BIT(out_disp_err)));
          WRITE(decM, STRING'("        "));
          WRITE(decM, BIT'(TO_BIT(any_err)));

          --B Outputs
          WRITE(decM, STRING'("           "));
          WRITE(decM, BIT_VECTOR'(TO_BITVECTOR(out_sym_disp_b)));
          WRITE(decM, STRING'("          "));
          WRITE(decM, BIT'(TO_BIT(out_code_err_b)));
          WRITE(decM, STRING'("      "));
          WRITE(decM, BIT'(TO_BIT(out_kout_b)));
          WRITE(decM, ' ');
          WRITE(decM, BIT_VECTOR'(TO_BITVECTOR(out_dout_b)));
          WRITE(decM, ' ');
          WRITE(decM, CONV_INTEGER(out_dout_b), justified => RIGHT, field => 10);
          WRITE(decM, STRING'("              "));
          WRITE(decM, BIT'(TO_BIT(out_disp_err_b)));
          WRITE(decM, STRING'("         "));
          WRITE(decM, BIT'(TO_BIT(any_err_b)));

          WRITE(decM, STRING'("           "));
          WRITE(decM, BIT_VECTOR'(TO_BITVECTOR(new_sym_disp)));

          WRITE(decM, STRING'("    "));
          IF (specmatcha) THEN
            WRITE(decM, STRING'("VALID-   "));
          ELSE
            WRITE(decM, string'("INVALID- "));
          END IF;

          IF (specmatchb) THEN
            WRITE(decM, STRING'("VALID+   "));
          else
            WRITE(decM, STRING'("INVALID+ "));
          END IF;

          WRITELINE(decmiffile, decM);

        ELSE
          --mif file output
          WRITE(decM, BIT_VECTOR'(TO_BITVECTOR(decout)));
          WRITELINE(decmiffile, decM);
        END IF;

      END IF;


    END IF;

  END PROCESS generate_mif_dec;


END xilinx;


