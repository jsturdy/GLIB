// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W0flajLaJv9GlILwd5pCPzG1FGpDRVzmm9oKsK1FNShKngYDG/D8rQLhHzbcAQhr
09kfobf2u3UAnZNeLaP9k5iyd7Gfgr4HEuuR91scjEqehWBDn0VDJNDycdrVlbk3
6S3N4xStu2PDp8rVQXI6qxhlXpgQ/D19+m2tNSrrink=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22496)
nBr7S+LjYe9894gn79O7jmJ4JO0YSAyeSANwdGocv9FA8w5mH70l8AE33oDtVPtN
03WYYAEzS+pgQr16NQQWwSz/kjEFqYRhEK3/BFaF5MIsWJQrip99drUthrOrLU2h
JFAw5l36IaUi0dP/nJ6ni9hFzhkVqqDYwLKpkgyKiLpBU9F6ZDHK3ZER6gZcCC+v
ZtaBUlVnkyQ9Xf5UEQb7gABwOZqJjn9pFOsBNiOJqKZYSE+h4O1mOpjhmIUgKaKs
vns+aQc8pAQ0zty8Vll9TqL3y1TaNUlkj+QEhskSlV5vOij9VS5VjtarPnvelyCu
/ePr3H/5OfW/Ynn7bRPU7f16syxEdFFRleMPLvFUOSTd3NI257HWWBWk4wuROdaE
D7n3++/yFrGKlqbYVV6LeuUiaKoVmULWkGrHv5ml4pS1Ef0TRrQ5IsW5sw0dJ8Uj
WldQB98/e5/+g49+ACbYod+b6+NSrUlEUWJwVBH7H9OtswspoyfDMvgv/3uC1oDb
GBTDrMVksrKneEAV1nJiEhpjm3urGhVeXDQDQgY7ve9vcaTxXEGl5+97/tBB27wK
/yBKx2le3PtOpK2VINhVhk7zKxKLwknqPXIaMQ5kPHnysnabX10mmnJA0gnn+Dzy
BsCDgLXmb4oFmsIwnHuTQmrs+Uy8+F/bhF5aHQJstsMlgN063gCfjNfhj0JyE3Ba
18razoCiA6aYAOio0YtpzC4LTJ7ms1JItS/ObM1ntcTMbPO2ekMGC0qRrGTqc4+3
B78kkpWvTC8fmYV32Wto/bTG1mJ2jYd9dGhK6oeCLb7tZudvmg6vBCawORdrQvEt
FjviykANnv6YITpOkPRDUzQCUWqDz9wXJ6HD2P+Nd9P6xciHIxk7+8HtcwpYoIsp
HOv5hqtjY54yliTMLbGivfSuN6jDNTFRHCHntKensjDo2JH0vzpdduN1OqO7TW8J
U9cieTxDDtY33ageXuiTSRv78lnFBwLRybJ3adkqBuy4s8dGvbYVptLMJXbfKGmo
7Rpo5v4WX3YpQP/0ADOU0gFoZfPrBdpRb8U2613MeAgynAbM2VHZiRNBO49/ZqgU
wW+lYEi4bSFqboFhQvk0braPwrmK6mQrrYqoTik7LSPSC48hA/4HNR398Ad/P/IY
YpuL75dMgK7LKkG126hrniWQfq6l/Wj7qHNnhRY7NBilvh5f11Iacbtz2rnawDxa
9pT942EB5kqOie9MIXv87HmcjbaQPyuFisoXQBJM89A5s2ZACeX48N6UEtPdlGiB
16RQfSkA7KSunEAHjDNYWan6SseY/t5I9n91Khqhp3bcuV1Hpo7oULY1dImlpS6X
1MdZ6VDmW9v6RnCSl6c3z+q8P/1s9Ks4nrttlMrKDiL+iAZlkTtNEO2AZTmox+O4
Cb811l2qMj0eJvC0+F0pFofaaRnivPBw/l+vLO5hn1/MwWlRZh1wLnqfr5aciiKd
vTN1oRD215aZUVjHtdukNSTwngRTpTGrDH4nYRsgatxyBkZBSR6TqPpagUSM/YXN
LWwX0gCsKllnG7qNI49X7cZlVbhCDREj6kbrRrOTmykSYjCSdmFfPAjSovGB3zGD
vyGSfiX3jGl9FZbQAxKGZHycbKS4BOHWgZi7hQAc0gfaGf6+W3u2RFsadS9CzvPB
b9Y/C9PBBJwO8eYqgMRAEx52BSUnTKaxQVIsMTlnAemSaOB8EVJYIkLFPtH8GWf1
bszlV45hcW/dtjvjxnXSDB8w0ZWp5sjhMUi/Cm+13zMtUH+2Pt0wa3W6gxtHF93M
+I3MwDP+kmkVeJCkx+bLF1aH3KEDxc1Xm1SXgdDpLIsX/5bO+sLHdUvDnToxTglt
LuPw6tsdxd++kTbRhbYiSYZqamzd/Pfiw+wTj3qhBivys/n/r09kl29Yq0TOLgop
WZbSz2wp/pS2EuHfDYv2hDX3wajx2Uym8qiUe/MR/nTvBOJasbmAWBquiKBmt/uY
t32iOKn1sQIopbhdt/uJVmDF2bw+LLoaS5cpSUde6wflOqxasm64SN/WwkYmtiMu
lTF8Xineimpw8MYSZ9bhkD/YjNARSwMBkCnvhhKgWFrzPdQt1CBNKFKVSvP5t1VC
O9S23KlSax01S5tdzOBNyXQ+EUXIPTQeTanlzAigawv/zivNLhq1xE/rZZ/yYnT8
iwXk6ZUk1VTUQEqjOgVsMxpq0GysY1atv54quaE23DfPsfdBRnrdvUESmwP3BUmg
6d/knZ1/RD/6tHPXXAF8tFhMNgUgMfTx3BqhNGM7ZyZ5PyLqXjwO72hBCqug0Am7
tKKvvqjov5DSxSjGUfRNmjS4bWDnmPvWjuuo0zJFwa4qCGWjWfOP8w8sEblRIwyi
QEWcSixgzRNkgv5+/tUERdGtD99bqFm5tj6gmLB4SJ1SNJgVYaSQUk+xG3oiMb3f
HcJfj1hahgZd+NJIZLOp9xygomYoINTEQMRpOFVTz///DF46QXiYrCFp2KppmtuF
clvu7hdNOPKxCaZQOvPn8qMkK9IfqNppiYPRyzNWV9SxwozPtD3pLwrJc7dZfnRY
l0QPuFscYjGw5Yikvel+ABqvKZ1StXsr+uSBSf3IyVmXAFGW/Y4+zvo0P+RyGLMo
KRhrRkBTV7XIKAsP4RGuluAA5p87FVrP0cptAkliox/GeakIt/shN/dkj5CkfW6q
OBr8qlz34Vo7+U6/coY/Q0IBK/MJlWHw0B8IF0dOMePDosaVi/VJu0l7v4g6d1+R
OLhU5ZkzByOrql95rtzLTdBTo2qWMm39x6mIAXYyqe06q5H+GoPfEAK0cBIBXtRE
KdyI+bPsvCenw4Chu0alIP/2Barke2zP5NUmiQVCXnCGlbzGannOUF9zoobpahZv
sOFWFPHvpU1bd3hSUncUMjd/QQ05Aexlw6zIq61Oc8v+95nk8Pk5mffVJE/+jx9Q
8PmyYA7bgwFJJRseMXWRNf0GCEO3fpL0dvVC1ezI571mTreRgeQpG3AKuJWI/jrQ
IbKEvvsrj3o5+SKyicYgkB5ihIsJTac4HMyJoL+VfpQHdIqtyAp5o1g4/Ap3qWG3
cYdwP47smSAWhHtTBDpj3H0w3pV6dpDx2kWcA85v0QOV691Wv99f7CpI4X6Bcdrm
L3eYUDuDJwkL1xjJVICmswnvSgAUg3Sh0buf5GHWql7b6zVtDBQq6jOeaESE7U3p
V9+I1r4PVVHwDWo2lPoc2wtmJ25c4FyTLfI/7szpuwvAOMgPqfnPy8wNDohzE0qi
QwruBE04uMnNO+jGRmQKOQdntndPyBL/12XCKiaagfLnS0rF2TDGpeJrL5QRRu/i
7H/m6/ZOn25j0G7I17pTMCm4y5Z3MJjmTCAidByzdendVEWDEwsgRpXjfEufIHNc
N63MY+PwCIQ0zMjvS3r9wcXCB+OUZUrfXQa7M1pInFKTm9DsjkBTVXkHdE1pcuqG
gUnvZ6WS7gDiYpS9Gy/vdtNIZ32WpDznaCnWWo6dWWBgDkcAn+7f5Yazfa3P+LUc
z1cx23LrhYEyOBwyqpfGjWQU4FoSIwPdpTx/rVvU8kCV9WtYD4vVTsUp5rsSmbtE
J2+cmmpdoGVMpjEptrMOZtPVsoaphzjr4gAx/koGFi8y7dP0HCraxaTI3n17I+Va
Ahod6YI35qmqH2qCLC5MA9G2euazAdj6fjLJidygPYbx9IpsdlvzySWlnABTaZhQ
xiir/tPk5x0TQjBuBw+gYzHsC1Ox9Rfiws5jH+BTtpW+ZLIITDwglS2HN7qSkxwh
S25mFHm/LVa8cYXiD1kECdFTxLblQ3JzAjeBLjGLB6Pl41J06M/uXoxx6shMe6nY
fW3zBuh7FpI5Iz06d4ZjyNKPrE4HwzUJ58dCZ2XIKbCR9owlib5oSDbDl5reLVtX
E9POiZHoqoE+8u5A/A5XiUixXXg8IkkPgAl/PHXzH64zhAlj6uC5Icn7+PowTUBx
mW6/m+EgzVm2IdF45P2kMXRsTacU9H3MGKcKc9YEE7IyvbwPoVSXUS5lhDtJkZQw
kzvNXd05c796SinXw3dtodBF6Y8XICAf9SRBde79+6aaxBhyFhRVLHIHyp+ahh3I
uhtQ4bw+/pSQi4JHhiOYRzLgLgvXdQ+Q3PumwNGxIo4iIP9eqXKXeMxnDxi9elU2
EES1LwnpEVRstVU6Xp/3LqdeYLg9cqOTeEZm8j+PO1x1KycofrMXcRI7Rtg5pIF9
RmAF9dD9JPStYVysIz4gFYkuHjF0XLgW94yIUBzLq4HRYVWeCWHhMTU6rCsyc3r4
nECXl9QDDfvEuygKkbsmAD0smPMF2nGuQApkYulCbjv9RVemvkQ6BqqhmEz7n4ku
c8NQTmJC58/k6gaitagKaFUb1UxZJLms+sv6hB8udhXnV7vX/6B95YBQ6/8tOnoM
Jiaqr9IXCFfv2VuYYuUquDkB5shJZsHnl/OdnNeDavs1uogagENRGU0zSPtF0RsQ
RjsAcg6sLY8ONAid6YYkXTuGsxyW02QCXi8WlL0Q5s81UgL6WND5iIRFbCzkM4Jr
ZVJYrwh/AaJng8tsNRz0/K1VQs4gQieE9FnUq2M3icxzzjwvdvz4Ae9kNot7cdXl
8C8G/RUbjpS7dDTiN/qsUh65YN2LWgZZC2N7OQyvo+bvEzLwfJhuNVevLMt7f5pA
fS3VzkMYKWsfj70ogLz1LBwx2WJ0SlCbsgRsV4LraArXQJMwf+1w01lvnimgnnHl
pN4a3454FT6XHp8juPShGode8oB1t/XOIB0o7vj5Fup5aEnpG3DiOrsiWawFz//M
V7vEwED4ZkxapyuF8UFiA9vWZMiMCX2lE3I+IvlNxsAzM9MBvRL812Xv59d/VPUy
AVM4YATwVoDAGZXT9XrplfOgeOb8vJh4qB3ZkyhcM4Oz8n1jXVWWiBed4QaDLXsY
vgkQpOTt47ORcwDLRzjRbGwaTHb1GAgkro4i/hACMegs4qK5BntJBk3rkmL1YbpC
uhpw7MCqat7I2eQnZGIxdXG5kn8r6nkSGmgfDpTcSuOAIS9UW8aKvxioJt/tqoZy
aXPZsPmJdJ/a1PXLbROBOcFU0+GfKq5zwkUu5F75zNu/J1y95cellI7i4vsQHM6+
/MuCbFWC/+qcWjyN1x2TKPPwMxAaeFPNdID3o7Kmb5xEUplMaqsrmXJWBA5sJKKe
ad7l1nHPBdP1ff7cDBufR04D5+UA2M8JvP3xNoTb6+BIlgR45VQTSWOtDYG4Lr2k
GyrHdzKUqGBO+lA9ysluzTnvba83Yj/cSP3FEzCPZET0DZ5S7MHM3fkdZX+Mxeqy
ihR1JZrhpHxPzZQiydoZw9c3+4oGqAIa6965pwx7PoPNOXG3XnoTA+GPdYmJ5oFm
YVQY8L0VmttXeFYK1cHv92rU39vBhOmKhkmbocLXaudS14LUSjI+QZbiu+XzRVWQ
PBOdwJOcr1k2L1eno9uHzAvuhkdhJp7O5z0UCdSs6xFhrgQvJ3YtAlNvzQvOK+8H
UxtB+FYLPJahhx7Maltbm13gA4FOf3ayjR6TIE0cAaZ5gQXuoHNjvpqVht9H5+3q
hHIt9DRLd/MAzVHhPWH0cO42cLyrwKuRPWXca/njzKan108iKZeDEGeDKmpFQE3G
ve6ZOM2K3C/gTsbAMGIOvP5Uew+Viz4GphQgMK+vby+B0BC5kKqTcL1VfsvUeVmr
4EJUzcv9WNB1sgM1Qn2bxgtAKW9/UoIQRBpYItoAXp+/UyRd9LjFhrLsA6W+z3JH
Z7DbapqL1BMjaSmiS1v045ihOWqqev+4V5hDeM2lfp5vgpZu1yqvrp/RdjOzgiE/
3HVESYLq+DPxvqBhoyWyXMEQWHcQCiiAefoubOuZ8eu52mXZNy58v/giYPhBf2Tw
2XvbcoczCmWob8H552uxX8RAqS5evv4ypVNjiJjRPN1kpl+sGcI/RPEE7jfs7taU
iZh7EDdyr9n7Ew6KmsKaR5bgl3BMqtQ9yMDrhOF9lhRw4ozV6N6UlgXXbqAczK3i
4d+IDmSYcWCg2pUeIf2BG1QYglYe8nXtMlUCf0jLHt0SzcIpL22VLIPZ5ns4Cbxh
gECi0qy2U8+rDdltAaTzBRimLQnQef7cdNLHtrbthyPe0MdRCOvjtdxQF8klmIMj
dJ6MPNFa4fU9GU3pQ+WOkfLh0eceXMILNDr5TNpL135dEcWIk4WxjLiAVb2oY4Bu
WL0AYKfUsrUyMNlbKHsLFPw3E7+M2c7owCUkfav2YjaSNS5Ad0oFJPqZYjJ0qF5b
it2ba19nV2z/95f6fVGrDLw5/Olvi5iSutmTqdWxzMLCj8HczoWQXzDh0MPNr5D5
qwIM0iqvO6Fnpz23qq53a88x8Aq2RtxJe0FlxoACPonCPNvsyGo3sKfMJDxASznG
C/MQEMneYKhq9Qbo2zGf4qLj6xC0NOIgHnG0GqlDbuNp4gux+bpjcNEntj/5lfEI
ANQ9RJB6zFLpgYgFA1QSxrXuUXEBwua5yKnNLt/UbwJ8p24wOuGcOr912l5+iRdA
1Iw7EEcVchQG3OgOVIGRU+82lK/had/f1xRFYk2jEeQP04J7xSnLdETIIbYOLcGB
ST3VAHkB6wK00bDv3qbvZviswb52btWP9bL06ilZam6C/7MEHeQEUg2WazvYuNCV
FRRvThpd4Mk5PPD5axDYr7L6SZVFzni9G+Lmitvo5lRO2UA4av79E9ASlF2i83WV
CfTZe/mwk055glUyp1Vvm6ZaJQXB2KBDy63OZUZYyitPDL57jmSIwATMFeEZE9xb
ADq5wUgDLLGJQix+Dta4NrWwZKjVHnylM7CkTn1N0d1tEbQWqOiepXz26e/2DscW
PKtwXujrk7S0nk4J8m3sEyxJog6VJLsXKNZAxQv5odZmoPwl7JXXEbp4C7bX52RZ
2rHUHkXgUxxQKuc/ulttHUSgBn7LwTnhN74fk1Rcxwy+NDVD1N/EswWNFYmodGRk
ifyhTSjqsXlIySyqaHezK2SyBZsZ8iOjZ++ul+EBNh0x39t8RGHUIcK43hKqXw0r
qTLnL74VjIpWoswr23HXg67HNoDAt2V+pcH37Bl1+LkAmuvWh/zwvzOEkQCrUYmu
0Y13Gi1p1E6n55gbYDbAcGXtLBVAkJWQc+I0KWA/E32rkAXvH3Q0zbsj8TQ8w1R2
60avSOg14ZkkURc7CaiCGkkbHjiwR3PxEIamfZQ9FC/zSkjyVpM3uAci47zhn0HW
xGcElvSpvFUcHDBOLcVgWGNHi4mDZ04B9dfE4MpOu0coRr1wdXPt2e14R+6qu2oJ
QfPV6KdnhpQ7Csf55N2zdKpxW8rtD+Zu99m0YZ+/1aqW2fPLq8o/upRLOaNsUjI+
rHQ/jUEgywKThHB2nUFTbPC0CGipBAfmTA5HvpPd1rU93If/6oa+YweRbOzI4ptC
p8/f/f03GhsDXiuItrybw06vTCNT1+dy723kR5JZh7njWS4Jlj1/thGSkxpBKmVh
JN5kwQeSs5MwQVMUyGXzSPUSsttuZ+dLbet6RvYPWFeM7K3E87m4WfOqKKysMrYo
5VPg6KqkbnPxyzj/49Vah47BMTt23IhgIGMYq9oXKafdGjkWc0VnSF7rH7QXJ1jY
gWYwtEm6cVTBrXVC/L7HLazeJ61XcmtGoes6/42UOqYmQiz9ujLT5RNvMCj3rgNX
ZHbUMUTHH7xbUkreQQZWLSDmocqLG/aqcm8gycj/k5ZpqXSVrhFGMgydMQeVQ5kv
tyVmswemaPvMfivut4+0Qj+t+IKezsFr2lzVmogu32CobO+z7uwym2v0f4T2HYOR
SvMKBK63cVUB60GOBMMGwNg0Wl6W3voJIjgOBzQYqtFIMD7DQsKdnTtvG6daY5Yv
iO5oI+Cxz9kmebA2BaWxHwKtQLW0NX0xIIKUMN5O/M0EskHREYXWir/w5Jv7rvJk
ECJwCiUJn2N5oTmHfZf3ojPQ2oioV4919s8Ma2/QUniaN8wEZ9vNKWnXItqTIUit
OudqKrFni0mYiszsoH+399GVLyitiIh2c4S+CdnBf9J0xBRqWHZVBgJhNP+cCEUo
P7NMMyAB12ah/a7bbO1GtRJQ64vDyqVxdTKNiELPCtQpY+ZYUoGsWn9fcm8hAVk0
CYRtc6P096e3SaEhDzA+FX7K6j2Xe0wr5WoRR6EciJhV8m5DLbPQTLyUKp1LlMY7
admQJCFtMOHEsgFsulF14KWj6vyCliD8kBgGy9TUsg2b/PWZ9pCjk3ARxARN0j2Y
KuQ+OK8kIoI8CJiqp1g4vxQ408l9nxTKmj6jcr4P6clF+mX60kK6BdpIN38O2Qnx
MzcQA7xgCrUp2yaSADy5q2XMqR1nsqYOA/UTwWrXT28ipTxdkQQZzR78SlnAbaD4
St9xL+kLcTrrxfwhZueanQSHxlOnJhQL2pK2cG3iyEfqjBtP5XqHmdtT6AC/Druq
CRUScVqbPKvj2QxdJWna19DHsuEmCdfNgwg9qv0F37M80coyHz0qWwBuhEJdy1Sd
7BPhnjtZ/TTu+WDO6JVPpI/Qdjw9XcapmkmBwHfFRmOB9k+SjTqag4dekXgxRlxN
VzWkfAYG64W6f34v3GUrH4R4pPoGEkgchQ01oC6GsXpkiHioT3Ma6OgZ7Okdsn48
vy2hdh/DE7RBJkvZWnnMaZFF/VRoDTvhIPMJ1Otif2KAXreXCgetP81SrzI6K13D
vLrBv2FFlItbPHMmmcWMz2EeC9YgxBju+M5KJgdE/q8CW+xe3jNXrJ77sybv1lxU
961Vlq6KsgCnytzEnMJ9m1T4w0Y9ZUbekP50c+ze3mShQNeBHyoa4O0YCPm/+jY0
5/HdrFrUYdyRQQ7OcvbUntkTEJF+xZ7G5TVGx89+WVCCoxQlGOcHJCnkwVUHq5Vs
f2TTvatqBH8hv3t7KYoDWGw6eJOqx0vaoOAi+fys2C5sQ/A58DNNByYKYFLJdcuO
HF1cXljk8lAmPgDFyypVCGVygiXCa7cx/70IDQb+h9CtW/o71hVJv0N0nz0kIwul
8YnBKiApHIO98ldZgAMB8qijnN6Bi0oTStYsoDC6+vuW7CFJWOmeFQhZdDIWpHFl
FKRnD0+KiJCBuMzYMsDvbi4yUhwRNZ8rxzZEKjnxGED6tkVAlj91Nh3aqj98NoyU
84IDiWLVRIvTr0UwakDpDZilEOp5sB/PXGu7xNuWBk+ExDB3Ed2o8TFVAxcjpS0Q
4ByQj0jqDh6TTdKHyeJKoeWQLu2CO9sGTluyycC6KOxBhn276nUzDU2I2BrgT4P+
l1NxcT9U+hRuYFRbn113P7fpPN1sx8ok2D09QCh/MAtjqeOUTagfHMK/pgE8dPk8
p3kDgd6OGEuxR+NglTUHffIcOdmWFTjwaCSIRRhO4VnpDlqeTP8atFgjMDvduB4l
DVEM1BSgvNsqWdgJAO5ZjvlC4yRbgPLg0Gfo6EAWmHCgpAn/JCbavwfi85v7oINK
tJHTVBcYFJiICY/9qpXqk42t3haKG1HV8FLrE1TBIXRYJC+zUfiC0gZc/YQcx2Y5
YQFf16oyXQ8mkzQHvon/sk7VZ35kQ4XjrbG2OOfkcwWYbKGU5OKylcUSBhOLXwM+
Zv4ljKFlY0lG63RdOh82AKBlqPe0h8jW6kOze4FJzDJaawZSSfGGv97wqk0aqyUG
xyy7jF3T8dyLiphKV51TBN1ByREvYkMaKBXLRGPL3lrsEtif9AeoKKYT54UbRZa3
CxvrwcyxiO7ELUmjQbqGyxMJ43up9BJYiTO6U+nbSm+91bd5Y/cVzzwpTRt9pS3w
dNnpXoRv0+AWTVkco2uWEMBNZxDe5kc8HN+qlFyIOIDViPgeMuWXuGlFhGyGOsJO
51Gg49FQ3CSLq2Dar4EhkppY/ctqawYvKGujCQsKhorXc5PImJvJO9ilFff8UYVp
dJlgYh0eAKGG1oaL7HxlQaFyMnDI9HU5fot7vcKpIpFrnNkwjRCfzoAWlZcSSs0u
FaiuU8Z88GVXplT6eKKWrwsEqeVUaIvE6mmwmsLK+lNbY82kJUYXeOqPAHPye2R7
Sj2lGmppPbFsDToDstAaVDtz1CEoeYolwVa2UxxS3dMxaQwfVnleK4Ibw0IMmmqW
mq6jR+590//D+G3YuUtida5+0eb6eEDfPgympX+cjUDpFvzDWFwYuo/mj+qgud9t
PR1hJQl3UdahQuPZhlTNCov6tUkwGoOM0qgv/zxBzlSq/orH3CgFvJqLHv66nWhe
bi+eIBcamNHFRL9apV44uEa2x9mWOz84WA3WJ0vuOFlV6U77yEij/amrbBsC2MZt
ZEl4mJHE9TdX1717tEfGj80ikQRi6ijGHZmmOp3RTLTRoS9zYYtZdFKtewz86rut
bHJylBDvCh/6AGLYCDYooMof3OYCAcd3aCGuYppWeXLlO3NZNMNfSJywI+P0Y0Ca
zCuaSrRSNEIKTxYqEk2+XMIuloMwv2n3/sYcXIwx9xlWJi/VG2gdFiEwYbYG1QvB
ApnP3xnz/DlToDPxAsuvKJalk3+8T+PbVm7o9dyEEgPzifSXfifLB8SJgriwMBDN
xb4X3UOD/RB/wA4ZDF7kC+RZuflzL9WQZC/eFK4vIcSOfIGbRBAYp1HHxC8rblNj
J8SRS9VLiub0jCJJlediIwBNi5Z5IV0EDL1A1mVKC0TIp1BdZC2buoXC9LlhhmQH
vWPhVTki/vUBKZrRYr1ZL+ezfpFToq8CpLBat+q4lGiUZw+D9aCvbgEbU9A6GKfw
+o04Qnp9IUt5vBL8SHqUkOmeFrW7zFJyZzYcyfvNprtGY9+75iNi5e7bZEPydHYc
kS/H4EPbzNyOj2dSXTqfc/GaOw0nX+r39E4VyCuthJIVMcY8RwzcJ1IBkeNp9cCv
77zXTa4LtgioEJ9iQx23Ju3Z/t6TbeevaZmuKG1bbpUNWNhZMlHjFJAkBCEEXy4t
V/KURULA6vonKYrgc5mxrOZq0P9mlpU2Dfztkcpb3dUuqdA7AdaJnkx4XXnf6YAT
pOivlbxhcHANsVoVT+DDeVVu6EqCF8+D2nKdbkZOv5tdJjGR05o5DBg8lRd6dJBF
VdqtE5jz63A+vpcALszzCJ0Edl/7s3/LwFFXRIRJHHPApcXdC5KUn0k5vwGC9Qv1
dyLO2DHKmvCLa8RALofr20nD7faBsP0Cgwc08T5gQ+9ijY5tzddPrbmxYy4fSEfI
rhYdAt9K/8vbgdtoB0lrVQMk50bLIwFoyjH6r1THFfDDPEdK54vxWJ2vuLt1v+Dz
tpKSkGjXE/WTZIQTSUnqk5Tw+L4DOzqaXTsrJeXkHOIsOS55dcmflDkDJmAM01CJ
2FFGOx4TvDmnBty5e6ECc4HQ1RSbzU7XuVXImkHovEudU1J+HCMLLLyRGs1BMG9E
SN0o9h5hrSDHARzOxNHHdlIu4ynn2MVTG/pOJ6+qHFV/qoeGHq+SxXuP3Fc16QEM
grzxlrNCyExa/LY8MKSD7ZqvkaIVg8k2xheiLjvGXXwRaGA+POLj9P8z0XLs9Rff
WudfPrjPt7sbF10HI+nF/ifC8larjynG4Ex4rDosIlpZjLdSM3zRgWs371o7bD0v
8Gi2AGwaOybBvW+qQXJ+dR/adgLybZOB5IiAKN48ql2O8GsdvoFbTT0S8zEStqAV
I9sYEWR5W2W/Zc+/vHZMtO/Bh40zrXOOZ4g/CHjcnsbCEULOhiGODLXLegz6OdDu
YB20aLPIkpMopckkWaKvpL+3pv8f1xL9R+5cBpfsfNjOYM+3+BL15NAhYEmPnqVF
wcUsXE69mQNm0qsLgozqrrrDwZ+sAu0c8z86dW2qBbJFfr9OHTTVo4fv3ityhgsX
K0m6fyPfoDjexjDslIc+/RwB5f96sRhMD6cUr4T1VAcPRauOjwZwW2HbgISbpfgp
WhD/g4A/gg8FvI7sXSusTNzGKuVo3I/MlG3UntQvY3EDePopjeKsZIwMoadNA/Av
HwDbEr5aH0YmJ4Ifoi6ylCBWQWeDslT8cGM5U22RKnJ4gHojOBmcrZQDxy4E+X9T
W72LmR3rVeoCIbRXlKUvQai/jOryZ8+4JGfX+YLub1uC8/EFnGoVzxxLzNaqLIDv
qj5JgMP7WGWca98h7sqFzodz2/5Bj4vCRkEv1gRv4vw5UXiKLOtQI2J1/rjM5L/5
Co+zxV2xVWvyz53rJ7ZJ9RwR908UNJo3eFvFk9zfj2ypvhfTuB7sPYwB9hU1RrPd
5RsCH6D4awRPENs+3B5xh3OjuMLGxh5x2SwJ4lW1UgxfkJtABP9Nu5Yurro5lbv3
H/y7cZoJkBWOPcuG9Sy0VmNpi4v2LYGC08jgM/AANAfBnx699DttT4tzIHOaB+sX
m+R62xQn18LyysRqXVq63VtEtZ2Njr0RoKXTkrwfSlD5Kn90Zsws/usO2o5uozJF
OTl0dU4LbqVBY1Xk4afci4lSYA33QsjI9JiqGGE3mFUgbuQes7KXm56d/vPasH0L
ADrWQsgE/N+1YDLBrX7AhdBGJDmEssDh1n+BRQUC3eEX3yb+KeGZO5uKl1haydZB
F+59UW8P1StUQkIHt5V45WcS8egv5ShDxE4Z8NBlaEo9sCsioJFi7ARKmmxqBXBb
MtER3n8BVs7WbQSqdpnWhqqhOizEQ/hHiFitLK+5HpD4xQzAuw40DgxvM2WrDmUl
uZ/0++kZePXd+fVRnVjidfqSK5zMWjU9qyrsXK2mMdodI7fn7tVcJ5i+DqwZo4/E
0GqtX7PScafL9fj7kcE+dSDXu6Ndbr4EoN5iqvbBR17+KpQaPNq8KCGxAu9U8SVW
+k4EAzmIoW+A/Rx1BhNLl6BN0JhPgXXw2QRkGAgicLtALOZDlwuTdzJzFsjkSfPF
eiMH6Bx7gPlN4Jh5rmIzsgw2HWJyWyxo7IuTW/oRoToljuVIL8BrDEy8C72r28Bj
z7Pd5dITOOCb2Xbju7rXGM/xiCyzKZETN2X7DoXt4JW2dWs6xd1/mnWNcmYAKnPl
E1pOuQurPiQf4oCbQKZxvVylVzQ/76eKr3ewa1Zg9SWpcG16kllOTgggoONzE5Ps
EsEy9BUQ00Bh+zJ86zY8qW8/maNId8BD/omz5e++2B6wzOse4zrYEqlaCC1o0ng4
MXrrInWihZJM0BwOxHNvl0veTQGM+ifojDKZinxjV+IKquDVeZ/INbo5EzsxpA1S
YqHPEQ4OaYuNFaRFV1XzL7AAwDLiKQUEqSlLD4D+keRytcneJjpFa7gcOm+A2PbH
pwH2oA6E090tx0GLAM57ldVfRXtDOtnBddU6+BiId/ZijcG45loAEth+IWdGxh9v
3nYCqDFqs/4gvIW5r89MkWuKTeA8ArG2gVEkZKBLkeOZ9JyefbRwcj4xwJ7Wv3ee
BBUGIHxNHkg0XWOSphM4AEHqY5G4oXlOpN8z0KxumfM7pZ4zx2L+NrIkxfh5uobQ
+qChOiHpAVsFSqbWUAaSRFkEexnWS84L+2El2BVgNnLgmAWYWU1HxzMoifYhwDKW
XEBVaVtveNoIdrmjItnP1iBTueOmm66E4nqN6tCUY46BnADuFAJmyfAx/cqJh87D
8f0RSbcap1pvidlDJrxXUQlGhb0xGR/AKVpyc1XtKEUGo6sP7EkLf0uijCh+HUEr
RqK2HVL6SNp2Qw61/xkiSl6WQaY8BLSXhv4MEqxl9UhndS5ZBHEVOqf+b+CWXURg
CzU7kyNpugdgIUUeFMD5q01JxRpePW2AlEZyxG5+rkhsacw7+Hwo0y/BY4AKihvw
93CoufDPPjDvuC0EDerzr1bJyv/JBtcZq3mcnjb7o7BYfUhPj/zI1FHOTSiIUNEL
/2g64Tzhiu+jISPOavxBbuUMlPaOc3IHXNyLTCkJLruJQs4V+BVUUhrag3Eb1Fjv
mL0RjCsiqleNW3ANDNJhZ7r2Q95gxeKcUq6b+37uhEduzDNvK0Ixcf3N2HzLsSFA
e8sERZN1xUaa9EVlI4kgTwRSIf2oOaiPhd6sYDMEYJ07tiEHv0in5XAGkSGdrzUK
QD28QFvRDZLL/p1dvejc3d9caAYqDy4mWb+ZgSlVQWyE1B8GcZFE7hfGmaPIdatG
I8ixPoER274ATwAzLwF/Tf/LC1n8TsccbPoAPwvPdaxjP/eJnWTYxid2mraf5TD8
JCY3C4JmOCCvmKxG4veUgv2bwMJ4pNTYWAWYKOlKP4WIuTgRXcLyhXK1xA2inT0/
shpotmnGF8uTD66t5KqJVnr7Omq7012uOZOtk1ZQtnTdTgz7P4IyE64oPPiv+BKk
ZFc6f5SRlD2pqw8NeGdJwOigfkhw92BhB2vykBPpPvaUs35OyJ4CSAkaR/cYkUhh
wpTPV30YYXRAzG9GmaW6msT2vZe26T8olVIRhzXJLzHZ7NEksJz9DN/PRI4SjCdw
3FUEVlUUBZDE9/YbNAsK/nhx8SXQPX7eveUifObYQZv87iWxNiJjkEFNNeSMADqY
ZSTvogQGfclHs75BuayQiniPGoKwrslFCmxysSnFNhncXVZq6yLlPpcQGUmGKilV
WpMYdt3+oAeR/RN+COzKemIeTFuk3dF4oS7sCJumZ2l2YnL5zfbT/5eCQNPo3H2S
C469jkSDv8XyM+baK+qhMJxVeGUH7hKUNVtffKtjp6FjoOY/47Tc0LpwAoE0LZ7D
CixCsJf7gfiZktUYKtjgg3N4L7+1cFxfNO1E77nwcTLDcFLdfdY1FRGe/g6SvoWv
SO2u5w7F23KCx8vWoa65yr0pqV9k125JuyvkjsANq+R/1ctXerimDxYBL84yWwaL
wGPZOa320BnNjowZCRc66SP1cfwrReTYdrcYc1kJrJ+XJiOkOmcvbrfjMp78Zuqd
W1CHi7T8uc0JNa/PC75lqyZUrKvZD3gBAnSFG06DM82Wfn26/Z0qkTHHCEKwh0eo
dgrjURMsi9a8LBNiDQQ2rHsLx0xu+1C74HQscHkFlk7yoeCBARAXfZtQruGNcO6N
8Jifho09e7XTd5xxqfQA6FxA709yRydTHjaswJzIPfBuU20bD6d0UBR2NJ9MaOI7
U+9Q3ykKFFhoL9yb0q5DK+TtmEuIge292BnjR5dGHRv/gKbUwjAPkEE97pj5DRD1
6r9ZFtyFx0Z6I1WvL89HVwHvIuQE7SU/FiBeouk1I9YRiSCbFCHJ51aaAg0x7oDw
8yMHhUCXcY/SejQZ50HBZedIODiHz8E1aM8iR5ls0SyCK38KhcsABgZKAnSoDT4Z
V0LRZmy++dtW/gh3vPdN1DNcSK8KqEamRJpUNqcGXzEiwAHejpsXRbIQj+1E6nvz
id2yGysnEPTpBAZ+JV7X69id+RqJmbgwLdnPeSqDrU2Os2JzgoC1N/5W5Rhjj1ZN
6vmBOXchjMseWOy+BwDUbhIkqKNZCuo67FUB/fouWuoNO+MgOtTEcGc/52zN0TUl
6gfsM0dfxK9NsSL/INjqNSO5NYAHezc3b5m13MokPOmCPxAT/RZzmHSDPVxzZWqb
NggZxE6vhDI40E2SjLNd3kNNuQ5hK3t1De6N6+84jNn86ZZuA3pXobwYwUjMGe4U
tQWTVgv3XOXDHqR2wsxbfJoo1N4Fl2Gx2Deicpg2DfcpZDEuTvrhBG9j2tMJbrEf
o2V7HYSiSqTUUeBI5/EnA+Yi3wvilnYf+AQAbnLh3Hn95m88mx235Vnjj3waaExD
aex3m2GjceRyqJPu0fhuexFgrvvFpN/B9yGwREl8AUtaK+XtVqO/0ziwRSgy6K4V
blaWDj1lcT0gOyeQauliujj+9v3IIRRf+UQj5b04a4j7GD1VyxVHFrSYBJPo4wXO
Oapm7DbaaL8j6TET07HPdd4DHYX4WkKa8pP+zV9cpAjn5n6BKgEZ7DM/5+yFKevR
KmYZWmdsHLXOPT//mj07oYkC94DCF1axi9fUmnwUbnj6P0q3g5Y5YXlvzsfNbJBT
coNHJzVumrmXG7ETf/tp7RrsFGIxWAAxWaOaBSAZ2o7nAYWVvnFAXi9nzHvBQZ2T
8yU2wlPUWUyZi5o9qnm2NtxXPMTDjIcjZuNjXyPfIJNZ0MqUqDMhoUW23Ek4+/kX
WGNCMaJBWKPod0JmC6iNKxd49thBnhIuReOHPyOn0WLW5z7QVtPQI/Lnz88reGfX
4IusOEfEPlev5d6dsEX+/t4o/0NFhayApZv8LBoZ8RD/cjb4cFxy6KFkEI9daWrh
TpmJSqDhLCjgLFt/mVmcHlleTsR9JQFAkGN7Cp/VVqwYplsFP8n3bcH1IcoLmS7i
IFJZpRk+1OmbOVoa0xTXcYUUdHb3wLfYHwx4wheFhIssJWxOHcC0X66dhSeDIShj
lt0/rM/SXITsLiZ+sKv3g/Dj8uM78bmHSSpOd8brbM7+ZpsNvkjEgbHB+SZe0F+9
x7eVMSUBqea0H3zREuUk0ilDKcE+yfaSvYpefVSNtIQ2sBbD6v+NZ7BQIfi9DfZz
f6C3Ok+axQVnygkUI0Qst+Owg37JAY0rJvH77dGD6wL7/nUYuOqakBoa4D5ff+mG
WW8dPl2R64bhDfcMePxVa1/tUyHvU8OJ1B5+HjoIZn5Qm9McVsj3A9pE9Xzo2QtJ
tj6h+oqm9vIQhlnF1hc6pEXi4C9Vmn3Dmq9wyDp5Fz4434U30x1mHv8clQuSuCYq
pDtGCle+KfrvtxcIYA3rOeFiAy3Nm4Rk/0U5gAB3HlJjVdrMqQIDiRJctxs9bhlu
9sMwYB89FAgfWq1hzGsP02IXM76YrXeBA5Q3ix79vnucRDo+gIfWYe0dx1fqZWLL
2eueo62X30QhmC4dpwoetx3mZcISYr3GKdXORvtwCSpp/s2fR/cPMFpCDBUDhQeI
OA9yX/gvjaScm+4KdSYHXJVp6mZsssVRWEkvVeuQkUFJIgnieigcWQzeEOyo9J+7
hJeYH+h+KH1IKLGraMt7js49QjewMPS9Vya/BYOrU1qoiF076Cns4AAnA8Ua0oS3
uTw90HC/ndJxv6qwS9Nd9zOzwhTH4LAF37gJbYO2sl2qzwOyd46kBULmI+oSuNHo
etFLbtkdPvldLaAfR+WHVuj5slrGEtarxolsgISXruhKzqmQwmzj1d8jGLrld8tn
S3Ik0CpAVEhatP2uf4AW7VR/bzR5pS6A/EE88QEkSjiHogeWfq6v7OAEBce/URTK
rXJmcM2G52Qa5/NdH7EOJUOUyC6dGkeir4+OpDDECU8NIsUVH7/UB0K5yf7ns7dn
TgyVc3Dyq1SBgOWJODFc2RXRJIKIRDbS9C/K5VS841E9M67pJssUpzpeaSylVBgf
PGGojWJV5ppjz6XHBzb7OxoV+nqIK0ock0Bag0mEFMki8FlSe3OW7OjVD2oFkCWp
rD4EDJBe7egvQzNjpm6up3dSLL99TadrSgXVHNTu3O/B2lM9QSZ7HcdSjdvYmsOc
sCmx4yKquX87s7NonZNde7Y00e2qfqnkv0MoLRoRLwHtqQhkx2IrBBqVVfi9NDbR
q2cldvyNr9TM29yFVmL+nRSPvFeRmuzsmEGm3FbG5wX+ZbjiWJPHYvqAQAkAcefC
f4kKq3FcdFMzYa925OvLe3Z0teD4vc+S2lDszRuyKto2XCCiIUN+vaDG9Ozymlph
FEA8FDeh+AhEBt+9NYhBkd+isbaDYsAIiTfvf3JEjvJ2hpXZGrAjJkH8pMrZeps4
hGWRaJkliALlNR28DHjzB+kSZ/p1cyL0rIQ5ZbEEC7sYOjZwtj5HFLnx7/Zw6kq6
dSnQkch0GnOlxkyk7YINX1am909FbkUDivSTu6zKe3zf2UjnnRj6TL9z17Z0lp2q
o/4bo2PgtSAUDQ3EdM1Rk5qmxCJ6pbAdawLMBoh5abwO8Tl0LV+UFaejiO8A0/2H
xpfGJGGYEL8iojAlLHFVWGuU4zZ0ItosU9AC52cHINTwEykZERNloOZkPeuOHSkH
cyVtcpUJp9IZNlrHMIBqVasdEqn427ZFFrDgxrv5Ak8n63kelrIb8MU4qrhM98/I
OvoVKeisnZEYrlRrGPnWn5ECR4EkOPIeWA/hREb1J96/i3trROUw6rw3bNY0y0S6
FAG9PNbAa0fkpobEMPeZ/Kqmn+IA9IH47UAGjFTJkt2GVGYQK/ZW4WUKsdJv/pCv
8P4Ub4PbzRP/dwBxixIHkEzDGAVOT5ERJ4yDFt4okBB/eObIvkvNyzA7ThL4OJET
ALjeICKYYlXNxqxC5vvL2OGc/Lv7eIsJgOztU29CrmsNwewLBJO8uwVLmLLij1Wg
GtokoJq3VMYoQwbuIWRnuGZDOGxtQvOXFAh34sVVQWFYa/PGVYBZBHbG72fYq5jy
IxeaiuZLbCHQimig+gef+2FossBwzcDN2sQztYotxeuVgFQVlylqYF5zRYLnW6Eb
v7L95NUrM0iwJchHxw5ylOL3nSDBR7GtP7YuQJOQXXl1kuN2NEAnXKaVrKdllmjm
GI1COKxESIDqTIPWitsDKSkAvzaKmCutFp4qgp7iTp11MF7jhaXAa2PYKN3F0VuU
FCFUh0EfVzW6tLbRBINczHo1lUIwn8ux2LqNsJ+YROf1TO/ziTdkD3zra4J2kyFf
JKTDvKlCruJxnuZHHTs+7ohnaMnQhyuapkt3Fk1ulOHXibgf7nWjlKmmQGRuV4zM
fx7XCYoCkcias4Xsmro0ZnpW5EpkT8D3IOkqkIxtuKdMyPQhXXKDyBYjd81xI1Y9
UKiaJ+ABrysdWIYXj+in7MoL55XGG6gtBF6yt3bBRm0C+NXIYnCM3JqyF0ijPYNh
HtPvqME6gPrJ+9J8w6/5iCOKdLXul1Lrp32/teNioJdCHIrYEEJSGKXCSU1RmOYw
Gyne8RTTBjdIgoovZGbjLpVO8SZVTfHRz3nj6MV/ISmBURb7WkctrGU78IzsEQEk
rt0LYxDyLh3MuKr4jl1eYxHAXo23fqGBTke6WZW7QsOy347DmSqekPsRrZQecPvK
Nwbenh6xj+zFu9BdEAvGrvW3LmU90XakoRt8JSZ2Rwv2f/75gNQqmYN8finvRG5A
0hn3WDABOa/Dkwwj4KpQXeUmtBmWolxygk+eBMV+U84dxKTm/EII4fFkFsQ81cAT
fv9DZwuMzgpIsGuVfD8kOWIUznDUEJSkprzTDJNqrCI1PZyquo9wD7GA1BNpq4Zb
OyE7xQ0WNPts9HALZOixfGuAnZjPo/PGY8TGBa1njgfcq1AWictJ0vwshXQqUk+0
ql8T3rLaFZ9R4cQuwnOAsYOweLmFKMSx+MDq8JRayHBrWq+rH5fPzpyBdD2hlLTR
Ea+zLlHlryR85uJlgVOUJt10d/M9TKPgpcGEgdNVjdgTP+fsmWqfDEqpQdCKVtXP
bZQ0salbsSBGUbd2RcV82mhi4Pro0ejh+cwSuWPRT7W9Suqmpk02gCAmbXZ4qh5s
uswtF829p6cNcBlr0gKNpb8Lds9XysoUBlK7g9OlY2DDLq/8wMKU1Ujlk6UB9hjh
uP3S9D7qTARUcRNBV5UZeMPRz6xpm7a8sCREoUuSb+j9yF/9XXkJnDRlWNbmf7ba
qWUe+kNzpgveglWoJb0IIZ6+Hv9BsLus953scyj6S2Rj4hriesihA6ICyU+IsQq5
6veZzyZBNcZw2ZMA6FlKA/rSSJPYALflPirfE202udawHdDJjrk226Dhqmu9TsRI
MqTEiuhOUkNCUztTTqxyctrzlAobRWb5p6grxyKDUkLIcWucohjeUC43zYr94VqE
M6veysFSiX58SWhx83i9kWLCDYnHkool+FMRrHB1d8mtjqmT88UKkv7pGcfgUpY7
cdDk14CtxB6o46tqER/ipnqWUn5Hwg41cU6QBc3x6WxKjMJ9lqsHsN4FU0ota+zu
TDXb6WaStcZrhvLoYC32A8+5pdpACgLrNujqeCbqpoAX3h4Gtnds80NU330plc5e
XFjE2OTpoJMsn5X8Bh8Vx/lo+g9n2ZbizHvsCRN6mStJSHMH1cqIVB6XiT2eb8Ru
u0Gt1vqoDtBsn+RdF/gYFiF4ftiLxpMze+U9daPY0MzOn8ej+o3+aN5/YtuxOKYn
Kwk1VPIop3+7ZTaoULB6nRWYOzrSKPaP9wMcqg8IZa8DjZuwdhk8zMK4xECmhW3z
2Khu88TjJpG1TTTXgIMlNBeEaVQlSoUJS6xa1q/p7/ggWzyJa1rZ96GRcPTShGaY
7VX/UHgSiRw4AjSd+0FAS5oQA7PutyQmdRdL8jB2kQxJSiaFH1YVOSqsmZaWaBdR
/KSQtD00xYEhJh3PGevZzwNg6m+6Ds2JgV91BhtZGLheagIowywQrBtFwf0lw7p0
4JyF/P1VjT8JXcEnYxiOa9+fPZPEijMk6KNme2BAQcZvpPPC3xVOssYVsRfh0XVG
0GOZP0VJqYFdrXar6BTFdMFE0o/mMB1GtjvJqY7mV62Qpb+k6bRMgVhVFEkkgBCD
FCAc4ZNa4YJX8BYyK8Iqy06GpBhxClnyKTT8wWD/jyGlSuZFqvkH6qRR7LMj3oNw
rQ//BtG7JrvXZjAypF/emBixcotR/+fSqN4RgnoWjfalqR6IEGwzhRbuUfQIGvWo
6BG9eljl9d91lHBMSGhOANVGN1gCHNLKp5Gvf8/AfnqMdZK1EFeHDVLc1xfKsMNR
5yvBd+Wxy3XaQkbKKJauLdvH93D6RgfRa8QaKHOhcQ/eIQbGVPzkzxefOGfXkaIy
XzUoSQxgfPGAQVms9yk+CHG2TZKhrb5RNo1HI0iDW/AYaJNtwtcRKKFGqfpIK6cw
skkSag2DiPc+J+clFVK4eu25UO21AA7YfjWcEf/GXjb5ufVP/v/9DYAd8nVn9Fib
cd/tHe+7StJXSJWxAYgwPRjGNer2uULGrCye0plgflkIHg0FkJjzmxsmVJNu8kE/
K+ogjGxywWa9JCYJkq3WDa2FhpmqRiet4H1hkg3d0hlO6agruNEyA+QCK7ha4sp9
siaIvCatvgTVfp9xgC3ZjBvdWWTkAJB1t5y9rwUqw8aeetJZYJ6ZAcpm0C12wWF6
onbE96t7OpO7UQ65TNO4Jcd2nh6IO+Z0ucgFHFhFH25pTLc5jo2I8zM7DF+2XGMU
Dvlip/b0TcEO5OzkVxHvCCjyykbC7AcooCoQbnEt5fXxZ8SCFNPm948pLP6rMcK1
9RiU4VIqb2uIgPjkNo3qN16PE8OOO8dinoiqmAsWOYpdaHple6mI+OL1ZYfZPS42
4upZKq8THn3OkVKWxHfj+cHZRUv+qI9EETBAwzV86dfDhTYhKCDnfrwd5RzUK67r
jO5WwavBMBfl5X2pBGSKTQl/LsckImjm7ud77A0eWzCwYuDMOM+mfMnxI6P6Wty3
n3BECZiepNxEe0OJE4S1Vsh8xx19wtZtfdnDEJqFFtLXWOqIaHFbHaGgpzX8o5XM
ZeqBj0u6Fg4XiDviljRjkwdMwCxn/0ugsMNx9764EJqtN5HtUf4Ohi6ENJPAoT+b
TlH77lzNco+ALI+8f2xe7qKOtAB4zc2DzU1odDtPOWnOZInzkVTR9+GW3h1BGw6o
SIsV5+8uM0LmrXkRCqlBLsgTrxk62gaOysnltHD7yw75CCIyQfqavjy++GWZBIq8
llKWJqgYMVteO9IAC5uUc/wfLD59ig/Jm2pdslomgt/A/BhaXmXrpsHswslmgHak
YpuL4q8LSfVqShz+k0Wt86gZw1EUe0i6hJwyV7++uFQYxDonrHjEdJRL6v3vUH2g
b9auXsQ/BIfApmr0NaezFndIVUxSXKNM7MpHu6GAZdorqhBfXCbPjPK6vqybmOzV
J0Uv+PrcleryAkAgqtHg7yIxwGbnubVd1rrfozHN0o54mcqjdb3uGYMAa4UHG0TA
34xiK1+8PDwNqiOCCtHZwVNmweIKR3mXn6j8Q2CTC1bRrqu07GGoJ6+ouub1BYWz
ilDHkng775G68LvRDAbri3r9sf6QVXQ4ImCfF2iVzAo/gzTHTxvwhjPsyDnFB22J
S9aPucIbOZs6gn/RlKCMeuern87BFQBr/l2kVxhar76nhRa3UlbRdZPItpga1IGG
kEy5KAgztTXWhav3G2/2dY8uQxIGf99R87UGKd7FexKGQZoMTMxynSAaj3vYd7nC
71C3GARQ4JjqaNuW4dyRAp2BPnVPdvSmTsbE8CyL35xNnPy0E0pWWe+DjtFJfRjI
Y31pTlDoZJwQRIZj9cKAfs0xwXhYyB8uha1RaK61fkYCOjtqE09DX/+XLOljxvTv
JiC7e9wQozZY7eePM6zeguIbjmBu7CdYrMHtX+mbye8pHk4KzXjF0r1mR1C5Cy42
3xPDqyrm1xhLh2Tz8Z+mnGZ0nCa9U0f7FrcFM+x1Bw/6MvJ5Zl+A/jBQjSLYtlmm
SNMais1mbFLllMAETWF0UmByanmiTcjDKk8vJzCqJyrV6GM2s9ro2ppVd0U+cVFp
T3inN8bHQJ8h7NyKqcDe77AKApxg9BJtCAHZkO4l/DwqD5tC6cs5TaViJGAxbus2
gvNv50yg5395yFIm6y3CrR4AeLsOhlGicdxpUGkVtM9hnt5Z70e3We9kTjb80/5y
EDg1umVhw/qNbJVIWEnor7dblCMsyJc96jcgKJ11OwhhWf7rIHGAyT5H5Z65qI5o
QVldG2CA2Xp20WJUD5h90wwnZiSJ+4yCcgLE+JRaoyEkdw7W50yRce6ulxem6ZCp
qJl6GgyBzX2DgNq73UG4u7YCes0mWtUOrKIrIFmEK/4qrnoEaSRMLC4KhyvnmBbG
qSijtf/G2txKZLP4j6oTB+9hD2Z0Xpl7wiu5k23cID1+5VwYrpCGJjpykethxjTe
wHGf+f1/tzVCvmFAA6kxTjz0gHkUPgwEJyLJ1mtoDmwo0q6QcIixG+xNBDdVQCqO
RK9yr4LWwvbLgxIg5xV/r0s0VaZz3GFw0Tf4YGqOrpInNoAF/rftLCMC4+Od2Vm3
Z8pSAULYjhZKMiu2OuiyYLGm9q1s2y7CgJBgFzW7c7b9Y0rMuDqeOivXpj6h4NDE
LXlBbd//lLUSEx49kONJ0YDGKp8ptc+h0JTxN5iWeNYaw9OwegPRiVd/CFU9/jE6
dxeYNX90OkC3ufcs+O1iRo9bz4wMnIlopo3dm8x1UsJ8bX6rLxfMECR96z1QQqPI
hxEAKpRScUksSd+7ZDMzm4pU1OBXWzdS0KlZ8+nNcr9/vEQgxweRCFkT+Rq9pwGL
2dj59A9Yyu7MpZJ4y6mDAqniedEIujqlS7UQ0u7Byjin5a+8z85q4dHYsld0I0OJ
ijjF2pOYE9P+qGF4xkxbWUQj8dGjPx8x4+hL85KkidcBKiNqmKxtH4xqaVIML60s
JHogLL5dfP19Oy6IQj9hTIkds6EVj3KzSMbvQV2y26+0b3wbKCIggVV8g3PLiKaj
P1qXIy8teHlr/8DLvXJYONyuqKWTDpAfeRs/au3Hbli7NXqsOHdfx9ly8ZKfDOVL
XYGyRWiCTkO+nT4ZkhPIQhEGI/XBDQmouOPBJ8fS3e8SXmKjC3rhnyUf1OZ1TKF9
FW8E2GOijU+vaCscRCqmVQPL8z6rwyCPsPMR8SZoS5FLgISKGs6m1W/1X4+Zm5Ug
Ew6GZ/9ZZ5cJT0kAIwazdWJBwwapakG+eSNdZO+Czi8lRDGPe56oJU0wjguVElL8
ET+g67iWdVU+FK0MMqDvYhS6gkV091A3Fo4Wc5SQK6s9aDlMy0uW5Mln9mWOMYGH
xkNugOCinn4nONABx/iCduoSWs08IHwpDwAoeBoMyNxhDzHidIe02Zj3VfXERf6H
6WBEofiGRoBAhCJ15yHb8M+3hm74ApkrnY/oquuxKV+IpNpjRX6J/ZcSqFP0FpQE
ouPh0bfyK8O3pWlaNeUXjURm/dFXQfsdzoXGNk6NgXDpV8f4OYIoK1j0m0uZ9kL1
FcKKVA5pw/7QnDK87G93Ma6+SdJRKQhxA28r3PFneomN7Eb+rBkZcD+XjsOyP6fp
JJtdi5d0BNjwXHuSPSCTAUSeOAskGMy6Fw76jqprxk9Fpq3Ufc3+Nwwr+JTGV50N
kK2kyD/D23nYBqsQ9ZThLVT6wv++SS1vikuRQ7ueq7v/vXCDubez6TGi7VUjHHGL
s++4eRr/MAtB5dinNWoJamhItfNWDzRkXKHcl9S/2aRD3NSwHKWnD/4SN/Zookr2
0XVxTikvLxiLxtcvjMmYY1cGCQGvX2jPTbl32yJ6V+DLjZ+hKSqBqf3Sz7t9mykM
6MQ9UOeUm3CNimjTSDhIgKLVZxe5qrro3IJx2eJOgeJanryglNGXTD4Gww9Fl3em
YBLOcknMBQ9NZjbRFXHwlBDfFe4wdMxv5Q4Rb+AbDBzROvNKm0vbmPx3SDocwl0u
SBrMaKa1dxeETmOYPNWKSklfhKoM9Dn2ovIqQuEJvSyyoTxkGuzhVC+hPP2opfLk
qVkA4esj8diBXNEyEYSYAf8lG34fyK2VHyS9T8/jZ6SLQhqge9DZH0lBUCmSaE+v
hw2h7Rhg9sroSZq0zhFQOPAcr93Cqe3VC2PXfae1EdgqJIZjBNEhdj4tA1l/OI1d
x7KySC1gSdih2DdibG5y9Cpb4Whz9MFI+dN7dglNt9hElZxgwn479YvdBwlx+/ai
jqmj1HyKAE6vje2p/CrT3PYz516cw/c+DPaIc6ZZG5JebuWGE/cljMbXQfG0Af5p
JCtZ4ekiw470ug9snKGJwtFPmleKwQFwgV628qJx6dFs1+BwO2ZYJ8HFNNw1gls/
iCkIYD59ya9Wq7z2vil/wOTdAg6ds8B9lwmptw39tIuK2CdHqZFrJSU8nje7WW6W
JdMMZ03nGWK8NyxyTZr5xUa+qUJ6Z08gYGyk2LB+M5Uj98NiqIvlxNzL7/D59KEg
mC9QJY7KvtkYFx+jM5GYaZAhbQro448KHFoOKrFX1YqxL/r4q/eh+DdZG3rsC8+A
BBljT7gjLoDimspaD2f/4Q1zCXH+Bot3yW2okNz8KayUi2/+Ly4UWN/oM9L2NJos
60dzbVxGWIan+DO+yEk3c10Jq38KWQqr/j0X6R4OkgvgVg+V7mEZ46DAIDsgs2Vb
Ca/5GAl6OJdRkG6QD7bQmajUEHUJjwHPVUprMuy15Pez8ltq6lXfQ1SuM7DYLjm9
kVzz30yOO92vtjFS7i58UQIqlaTRtZjbhVTdTSeCox6hUqQZTN8OMV5skZlP73qT
lqhZWpk5Tc/8apF7vRo2ChgWgHvEALiXFIp/2Rq2fHZGm5gB+7TtZ4Y/Cckv6I/O
mQIG5F5BYDBdGVbsKGM6jtxvUzyiTk9+BF3+SGbRZcUuOeN1Ao0HdfrmvMb3p5Fe
JiREbqbkzvW2K08kPIVe+h9shBuXws4o7rWxIceBlBQZsjmhvUj7uEtfW3nDIuG/
20W1QDwCObJlPReEGjcaf41q9Y0rLyEP8PXMKX3ZJxAsof2G5uPP+9g7YVCEcCGY
VTAlxn9n8cyYOL5wGgWMNjd8DQ8rkw0auKX1UPPZQnhLillzEk5wbBmxOwgSkzLj
nUF5wwK6s/ogRc3q2YsWYiZghLUtd5egJUSb5y6knQcCyR6ZKVQfxmUoS2Vxp0pR
Ke9rtDhskHhOQ4i9AZEYvbJdNO8mZ5ANZjLWcNEI7BrPZ9GO5bfEcRMK3ZXi91qV
kc3dTw7DD8ItztCKy2I+gZ1LRDlw/DTyRrlyVElD8VyU1/k0LrxLQsfrWL0/hmeE
/cfdyrYZeVlgMmJp1XPStkKiKiYpYOSBZwX2c2pwUhMZwrwjHS3AZ3O9Z9y6UGWk
+EIyTC+ho/BPM8mqGUfVzOQKem3PohTW2GWjnDuLHDeBuqmlrluueBA0k9xedX0u
MsXI6ixkECA2DZBzDzAB8oeOcyUOIZC1DdvqLIr+NyH/lbjDS31EdTag6jZXNhHX
IsQvkCMAnuypAppzksNGfyzZhRJclrsk/F4z/YNisBIRyl74qn0ajiSnKOqKKk8z
uO5pbCgDwdaPEks+1UseOuKlQhjcqSSlYMdYNVy9Elou3AxLRCp4S3zYbX/uK8KZ
pGIjBJRkuKwcEIXcTvsSomTwVFckcNXn6phGR5tb/U4dP5yINCR7CboY7Dr3Mz5g
Ify2EHPWYqTpTnwr5Pyv0/51XcbszcDwDo04Ddkn+HsfPuOUF5jMx0qK5x+O4ijL
lCCXrlczLG91PhNHYHN3mMG4ZxrQu7KSGdFOUxcguCFCngT5E+kRWmihEzPVvtjh
DmGAa1uANqUGNa4kqdxdb5lZJK4Z6aP0vq9QLJG1xUwNofuIFJ9MulZG7gHfsgSg
arwn4/eYAeYV5ALN9IZLTadZCPfU4Ezh2uTfbFXyfCXL0wB+oXRdpA8giYwsm7T8
Lct5rpP4mFAwPCnOkVYvrUgFyYrPwt/BlU9DaYfI0GXfKuoGhNFLVbzN6ra82lbQ
Xhq5zwCVDiVRCx4FlV2mJO+Uh9DC+4oRoZFdCg9rV5UikE2dmof59uIVFeJ5dKEY
CZHrW3hLzKQPsLvbgpLHHKtS9Kg5sP3UQ0jU4xBOJkeGR0HnBlWTUNKlKEzLPMqr
QCGC636wePXlTWLfKw3JN85xS33dzTF0SbBiQf5GrqohSmr3iri+1WxhWVq/a4tN
dfZWMtbxMMpmu9Hv4s4WnyXV2WYA1HfKt8YXwuih9DBdGS6K+QZw8vWOwVzX2A2h
s2wORQ5zLRpVXl1I4iNy+MdGZrH0BL/dUwFGOGa78UG4vWTbY8Q1H8GZCMmAPEry
3mODSvKkTkca6WpcaNXO8LD9Fn33L24Ia25fr3WiiWTjJQRCQVjjBQaxYsCzBO5O
hT6zXF4uvY9LdYiPKCRvyw9be9fChNxjmpvOjfkGPJJgB8Agqrp+YjLLO3ITHtfE
q3lKvBA05FcMMGl4KwXOITzTaqTi5eTL7YcmNuf3OhKz1K6glzbindCwzIXBBxRa
kbv2oGzKXhp3IBKX6phe0koTKnntgylbl/SB3h0caU2SrfRVWwL89vixmdI/RkRj
TsNyvGmQtOkLFHs5DakrMhEZr3yZUafdnKV3nPtUiScWMO/ahrfT3+OwUUr1P/ED
rEXb7obwEsNX5gRwtAXCa0K1jGJlvMxQprKyPitEv7RFhTJBvEEcvY3ILhk551Ht
J03Bh/VU6zSGRCSVRUa0RJQPDJ4yXXYqwKmbkeqaKA9iUhxWrII/8IQQF+208skw
vwEsr1PUJoJ8+DMNh1oqNLYmPDsoJysONHUoPY9mBOERzp7JShASLVFZT0Vm3+oJ
R2HHhVJ8g6Ng1/Q0ypZNkI0YYPamwxS1BZ6yUPYQCtilK5fKJUl6YNgfYL5uDG5x
Q8RjhZvjAyEwC+HbeIZVLB7216LVmW04WV+o5WI/s/6RqLgdyJ9hquiLnPAZT+TZ
mAXreBp4C81ixVefUEFFDvWiAlXViWhvckOy18edA7swMcwtj7KdrqmmPkES8yBb
kGZPMBq/jsKTYdc/HYpc97TKqqxy0S/lpqIWe2DMfQw871k/N4qR0UOytXzl0owE
bkXDOabgeRUAIhjkvNrzyqGuDkpKLQpD2js5q51qY7RK3cGJWDUy679mZJQivgv0
B1hlU6b4cQEEp1UVfL1YL4j6cIIK/lpX59af2V2twibw6+7pmT0GVjmA4wwgAUl7
vITlMh751P+zCyPzquft/kc9xdFzvuGyz7Uf2Ig7tKmsoT0JyUTIuNo6ZjE5enfW
6BY1hAwCMSBfRAuqNquEwtYKy07XiZ5XMtfgweXTWNupQzFPD0C0hK5FmlOlJskP
66Y01Xf+S+Fa1FVU8QcxXtkxV5RacHXmV7R+0ZNVsdfzhVAvLoSQfhCgcitkNL9f
xcRQTOQnmZrpiby0Bib9DY+nXTmawimxqpJfT9DAe+kvjxc7FcsAh3Sj36wK9Xfx
v0Dr1VjyyTf2QlxDXFZd0n7rgHJtsiDevayIWZw6ia0PJqK1n8RdDS48jCDBEKN1
aMaxPGkyQcLu1NuXjkjWQlEwTOjU/ZKKwRku5k2eDXGoRvuQS4l7/9kz4vVibCIK
ixVyqJjeIWSBHHIEcrKk1Kz86ZXkmvDEqBmrCGjMuN48Qv4BiMHPlwYimMX3iTTW
4fG6A10p+VazbtqDRAr4/9NpZEWmJZ5semPjVBXnM6GkW0E4OsJM8xh8SfSnB5M4
+nWQp8NTHpDKY+qhXcNWjbb9a17cVepmmIMmnDueMYQvHspJ0qbFa4vxAOgF3joQ
vYgInK2oAqI0hC9F2/DJhav2uniYOCNJvAdjjsPjGpJvvM3XkuFVptQUnmFyBHFp
J8R9gppC5vmal7TD/Jsug4dbmpITl7d6IQtHaiDOYfpJfp6IduUNaqR5wk2stiIy
GIy2PVK5Dwfd41OKm7NSyTYAjMQyV/5KPufB2zvm/JDs4gUAqz3NoUt+QOPkPmkJ
63dt4sCdGyLov1ficUdi4zHYOiuy+7Hv7DmBiX36zDA5U52+VCzpOghIwOcvIkP1
x+MEwK4v6tFLJkiMz6oucC/3wdm9/ik38lxrgeJqsAWYk/T4uzU8xzLJ5+qKdNrd
ZzANbk0Bp2lENMcTj2XgzMYfvjkhwNwrEKHGWuVVJylESQwEeVg0S9t9JYQYXnHg
iyAlpKahaFLtMDsYM/5ZJJyt63WAJsestPtvrYz2VSEVWSPSsF8N4gUEdN4GXizT
0W2I1wTkeuRDfrGWfNcr04SWd25Rf6mBDPBbf7MNsFIb716gNzS5kw4Ha00/tEoF
iPSTwrwW2IwU9VUJtdaxY41cA6soS48LJ5YlQAFAxECDKJ/VQSZJkvvUJ1P/7PEw
SsdbGNy3soWLRymYVizTqtH+CssAmV2Hjc5GNeHsxTpbXwkB4yOZSur0Rwce67bN
f+diSMD9CZ5ZulIXE5gEaRt3573EuEGBImta1+qKagifVEzyzT5pycE5y75l0tMD
nr7kKm2UcvHvKJnZjasQIA72J22w6fELvFcuUzbRb5QzroZC4lqD0l8r24G5tEz7
Ovmlj9+CBytRp9sh2AjskEQapsnpk2IlcOZ1lipVZPcW0X8KADYjI60aBNI1D4dL
yPGqzBuSxOnT5TUxbz8t76NVkCDlEVJS1EEJu71zLhYKyaf2fb5PH+5K86cMdba7
ruqVnZO68ZTeXZhU6prM1fYg9hNXLvHx+TEOYpjkcTnzZU8bVsJI/uHSX69ryM+3
GirPpASUDncrm0q96RLssphJuXlQI8EDO3zco5PzHVsAO/1QDa78b5rIbQ4f9rTL
kA36mJAhYt3CI/1e6AZK+apiJtkrq3WOhK1CPRPIExzx94k2E+JI1Qd5aRxPFqyy
sm3fczVdtKiIySrIgn6+k6Mo/0Tw065umf9ni6Xz7hu23Sf+poa+Xg2EfvuVsV6y
cZb0Z3pZBOBSw7gPOLT2lJL2j+adih52xi0kQkDNxfA9+J2JVvuh4TnQac9yN2dl
TljzT1yp/cMJjRaHz1EJ5DlBeCUpqm8sE0Sok1SuCK76rGxsnt9KhIt/RD+P4MpQ
Y0FzLriu7MTTELn/RZPkAcdYsJJzUGJ2dNauSCBkpVNXRElHnY+OD1Bom+R8wC+E
XNjrKRPbiTyEjhzz3vw04hRn86vg96rmg970R7eB9PpJWJXsh7GD+4G0fXLcDO8V
OSjhMUiUTZS64VhzAe1zUwHma/2VLkRwBL/K0PLBCk5YHJBotSnd6Lr1ItsA0QhU
/JiUe2eci2FWAv+rfyFE1O1JOAJEHIDo1M2YuuXxWbMJuw44+E2M599LSiS99OpT
l8ZrxET6/RKUYg22CtT6+B4PyMvwTj1nB2HfgiVhsT2DIRiKZnLuToRvwkltzq8P
6t0RJ6j0e8p8HKJ4mtFAuyC3pQjIcz5lDSs3PuGPKFnI+5M+pqRjzgKLOP06aGub
vA3uxtsrnsYzn/qR1YEM0QpQe3nmjUuRLhHZ5NMTaWtHDvxpd0pJt+lVJ8aZffzQ
dLYEn2yXwNm7R4L36dS2Pr3t9YakBcENEsHlDPpLDmZyruODdG3YbIoJ8apwA+da
THlSk3OZ81Q8IgjwXOAYL+ubxrP1O5qbuekMdWofEI8=
`pragma protect end_protected
