// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
khDaetTkwZVl59YJG+zqNb9/B8U/nT82DkG3EORyTOyN926e3IObYbFRpM19nzTi
j9zSEuAR+JUwzXh/MtIXz7dY2BqDvNI2AoV2emfcJ9wZXRRueUA8kWoqQzeOUa6L
Tn9nUBKXY8am3nLk4WXtziQzLBlgfN2nZ4wcbn4l40o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20768)
PKOp/0FM5tXbHudNplr0Ux92acBN0D0glu0BOVhL+XVrmg+chXQl8gBAJh0WECs4
jEzHsK834j5dPDtB+ZdJ1a0bwv6ZVUpzHHaN5CsDQtgZqe/9D5crkustQbJpv5t2
RAM6sl0VZvQSkAbzP7M7/yGw2EwUlK/C+Y0lHpDeiUytjsREEv+4CGnIFVFNR9AL
0GOVA+0qa3RZIKybinvLXYyMprd7+BpvvVp3PdcUe0T1srP/YzV4SF5kQ/q09zMK
pJo/3bStixnh85Rb+V/RhiIOiwixjsvpKv1mQzFiDrh8kkDLjENT8by8nbwOtpkE
aSGDGMDvL5r+xa0X9Wb5bP3m/3GDZVrCSxbKUKJSqCEkRn3uMrAZ96UGPzYHzDYP
84zKPGZte0ljdXWaV7mwC3hLNk05RGSirgrjnKvXpRV3boKVNJTyotwZBtdjMAQ+
Q1JHGklr/ln9biE3o1oJBxyfsE+PfgFI2rhHH6ETznPd9TZuMEL1yP629NqFTmK2
1D921DhGGRp0Op3/hiMSjpbBwlnaPWRnXGpM502vjDh7Qi4f3PiFpwbOADWrxPXj
CRhjd992SQPgN2VkQEPrKf8Pza27tplL4fxBhhnGl3v4ETh5HTjrC5m1rHl4YSf7
pQee8dyttbMqPHuntBcdqu4A3cOCjgQk1rMqNnyPhg+Bh9iSm3eAunoEjqAOAMuW
ovEXGL2YdcVbWnvuBWM2/l6gtE53bDQAvK2TWtbYkutspebmmORa3+rmjWeq+m73
nCnclK2NU3LCpFVysF/j6i9/rtcJYin2XrBEkkshjfJYgj7xbEnnj7JjrH7D/R3/
JsoEjYp9RQYVINQSaS6FWUSF3Dfg87/Sh1y0ELhBTbyRUZLOE3aPisO5qYs+q9fG
aBxZh/A/ubAEAH9LkIj6mhAlgiWiXHbQGAkfEfLsvrgEyLmJg15iAKYjUMd7JQyZ
Z/5d28IsVSEugUHnbBsAhFxN3dpbt2yG03hlOkyc+RgTe5imLG0VMgO5gfbuPxGG
wqsmj656yb0Cq9/efVYNUj3fp3OSi/iGKnRJm5JPk8GXQP5EuzP2lKimtSGmffzQ
kJvgFfI5xyVYJAg5Zt7WXGroSvJFlPLslhk7LToEkfsRpxzFUAqUr7NoRKHxXRKC
iabRWHfVlDsTWRi7RX15wCWXAv1I8X7KP/qvJCDhR7KQOiHKAj8SV4QDQ1YWIhfo
NOoa1YVoZU/XoLOPENJkYawRttC9SngEr3LEZIy0tCec9f0i4Z3wWXnP4XcLViur
34CLmol/mbAabQrXZ12oAZV0WqM0fNBhdhwxCpdHKjGPcAdyLl+FJg+MjVvxx/Bp
Az5GFoVpiHmN996uPYmBc/hpdStMdrhZMNnA350e7GhRv/QgWqN7DKnEirwtsbli
+YDE76CKjAB3q5z3Vd0K3v2E1aS4+7p22zyYdMkDxWCIHtz7QoJJbucx0CRtUUpo
8FjO7BMCNPaf3lK0RgD30YIcXfqPz/rrF4yqRJthcDPG6DMYeOAQ3j2D8dhnML1M
JxNCZ95VoYOoFjQUkUIEJMc1Zhsd8VgQ3c/zNFixumPUWra1aINm1LgihDrXc/+d
jtNZOZh0IXKhY3Lv/lYkBxzgBpHeuVwQT5Rk/F53YtKBnuI3FSsWOwlYyneBlfDo
ZQikMTCvGE25dtIGFaGxGx91Aw5eAezWNrireBz5+Ks9UBv2OqsIk7Rqu2CTViqY
nouueS8WYF1VlOrjhSSh4itlqAUdLGRxjqhSpIr9CtkMjM3JA5eTzbzMqiJECJc4
Bgj2GWkcSC4rp6aG5y0XQotF/nvJIMEwF2r0j4Cyv7Nbg7scrAJWC4Eb3G2vPSy8
HXIgp5/72ffnzlYzw8J6csl54bEzUVq8eSSy3uqPjQXxyDPB8j/l5ZRLp4SO5ZTl
4LhE0E/FN0DZYADRKpUQTvBZfrrT2g5GdfyAB3cTjz9OJ4v8/34spIzBo8QPvB59
lJaL1XhcsIK71FMTFxoerJ6kbPitooof34u08GG2F2xfJyS7+c2zW/kcKs3miFSa
XosF7OeoFK0ekEb2wyqD1qZchAme0+F3JpEp9lYT++N+bGVCwex/uFjE7B2gan/P
CvJvUEnT3TMqE/Abo9NM9Ey4D4Z4UaxbrqfantNSd9BO64EP2mWbfns4Ei64JHBU
8FaUSaL5pjRVa1O9/lOM9jTAHKpxmq6EfOVcvHDl+3joeIP8QI4wDJ29tyDJXclY
gl5mamRCEB4K6KHiW80/zq/A1G/ih9QxoKPs5lStxSim8NvotzcnUoKVn3srsPqO
j/xLrJ0o/2p77UbbK9rxbXklerI0hm6+Yhgl53NP6bo+RLRQHl4A0vhkc+ToI8i5
QeFCi8HkI3lNGoFSHI92sQQ9wm6BhABWSY7JbmdzZMMfUephBAGOTMj5u4Mn/dP3
W3gvqHynsL8QdtEDKM+Akzp2Ri/+Et0JQxzNH0xJQMFnrVLVy0rFwZKTN4WyZPfF
ITvMnmv02NywWSnac4lrcYlYKXOGUzbSUSU2CSLP/WmHBEQnB/IszHqUgCBM8VrW
JJKz4FLju5y++G3HH5OKsgzcnSgzbf5EIOKXds87zkGSa78zfDRstEcmM3HkhnOx
LZX2jb5mJJtl5AMMPJzcCs3irCtegBMuRU4o1Mp/244h//D4TjHdskYUM6HhI31Z
Qpk+dy/em2cpW6FiwUlHTM7nQ4L3k/EvZGPlYkoOd8Q/P0E4WSdpbafZV0rGMq8T
//LMiZAaPdUbEBEv6/l6os6YYY3IYgoVmp0pM+DQwVdk49Xr5ZjR4+5swDKNjTJG
U2m2OGtdCk/6e1stUGI+uP+8KnVNzc5mIDqIvojxfC7NYtAR/AgMpLMxpLF2x13w
gk3zJXcNW1AJHS3rDTTb7fVELXq2VK+3K6aw18x4KwGyZxXV80200eCKYZ8abe4W
IuMts+A8zch0aUNaCUFmN7XN3Hke+0BR4SEMfcc6TTDWskjRxjIQ0eorpx3t4zkz
HfyQn0JomnKNxfmIsovLPmDBRjugW4oVhvs6RkF8E6HPww4FSAJK3mR1CKXhK+tR
C75cJiAZEL4hcJrbrZrhj5o6Vh4eu7ZCVDiTF3PFTyKQAPfz1umzcAZxGU2xE/A3
nz7ySmD0ck1CR4Qq8XUIMfNipGIvpq4Dh/OKtEtZAsf9GQClME2IbDG49naozH7P
6uLB76kOB3Ko2Q2Rd2OMV0DNjN5E8tZqOr1cQs78yKq6vGW4lUX4CQ9sGqfLNWuv
sbnT9S+4Ea91xjcvMfIREgtX4o2wZR1WgwgrAf+EiUWXBGUbypO8ouBWEnfaNGK8
Sx4NCv0hD2dEkDP8We6Xofwy/a8Z2Xwh6+UjObcJzM7m5DFBXMdA6k0MKUC+zkhp
TWQKIutqYk+ZKaONtoVwQZv0I73YWn/znRrxLpqYYQZTqzfVPCxmiBWdiKKPOp8q
4DlgdiGbJPE5/3IepbaKxdsSwvyVO3IEzCgOM1nUUuoJveRfnIO5hsdshHmQ9WmC
TszyQ/67a6fdfHXtyqSeg0B7T+LffDQ1+ZP70Tsclu8wUZNegulV8AVIMksIr5NB
+lNruiJLH/ZKzXHWIoNQq7WVZLKUtJpB6vaAG/lCyFWDsqd6K96UYXdyon1SymfD
mDe8JTSu1ukWFuBfEbxQyy+NCvaG7PoPv/lPnwD2g0D0K7vlYXPHLSOhI+Nqas9m
aiBIYTTaYwvaul5Au8meHvgPBdjJ1RolWf5NkVlo7ZsmJOzOtwvYEotQfEqdAg9l
LP52DSMTsfA/evZTpGZbM71b+vc5nvgkVaLrA1Jt5JTWhI+kAp4H7c9+MLcgQG5i
oU/RfoalpUcWPKGXZpN3r0ji9F7HzA0LbDIeokSy3dPNTguJb+q4ND8y9ZH4osj1
URc7Qowb64J9qDO34XgUk2aN6FwTVtejtu9cOQMTMpMfTjXbhXwxar8X9mbhOjIp
4JOp2mN9rFOWVA7hoaSO9Zy/SwvzI9xCwwFSGjkcjsrqA/+gg8cO1ojLcx7/0u4P
AHmhxo430snXzV6y4alveFqdvK2XEha9tJ7+3uSqK9hYqp0eYD0Q0p69YHQ1BVwS
LKxEAKWHdEsIbJUY60j096rCGBwoFT0+hLx/ChRExws4fGGtgfW0RxGkKspuGik9
gz9KAc3Pa2sGScRYHJB/TYwES8NDjltJl5tQVT9zYlw2+ua20u99j3gDA35Th4pF
XsRUWb0KmfupBAe38+Sa9OD3GKcqM2RO5u4lspWz8bC3hILcUWrAPawnzg+Osv59
biwW9TP+D3TydgoZ4fO8QaErhH6por1kqv8lIy8x7Ul4Mjrkb1f/L+XbAG0IF2bN
D0+YEIynbfTc8W3DMjuXn8J27qkbm5rbbHRTLxBct2r9DOVsgOfyWMFlFZdWj7Zt
CyyvnPQZn8ZM78RtOk05gwYtQmerFG2aK9whQ30N4HI5jxccKg0+P5DN7cmzVD4i
MshUUs7cq/UHfk5AmqdKmbFFXwe0pvA5U+BDxs49MOyOEjnBykA6ZC5431La7A0O
uQCwn7MRSERMekpX37H3KcrIbpeF7sIFYaUdrutCFlUXVXKAc4oA7/CDGcguQbpf
ibb0BrmOaZmHsm75D3vINx6oRF1OlLKhjuVs6fyH7yUHc9lRgmZVLxE1SCZvKu1T
MjMx5SMW5mUISQYKbxMFIguKveM0x9WZ7xpQ7xxarCGDuDy/UDs+OGT4sjFp70vG
rSt7ejgzV6nGbmSJFpppTE6IG3L0Zh8XD0W0If8MGFdecWI1ObDY/cMEALWdjPaf
90t1v9pgry2iFltg1VcgC++PJ2dDnU4VLVzgxLSqUPXR6IkIsVw8vkZbAao1H+YH
uJXMQO/HVto1gHWQd49wbihoa5ClEUd9OMd3aHjYT8dKonUkXzPoiBktG82djlGm
t8Y8PbGXfS+snFqjaYsV3R0uIGJkU/UDmKZljCCCRSbV0u4LuYHip8Dj5Ec+fDuS
NXQborUFmbdCEE2KTaLyKTKinj/mW0Ih+dDXPEmPwnSm5JD2/HhubyNDkecHYTIG
EtwYmWDjVWyQakxs0ISaBhEmh0tYFKUEUhyfq7b8TU0PJussabZ0Ma7KQyXHdnm4
eFO3Mjun3MWa8E1UA22nMqbtJMTwg3HciZnQ66SHljDT2ozHzZPn49+0vfc0gZqP
svX4VCpEuiE0fgFZu/PIcMX6zjFuCNwQVt8A2w9A1BN1BDvZFYRpgeNGSINOG7CN
sq1y31YPmcR90JMxwcyihoiI8U12Q/hfwTaxdbhFOkagbVjt6oQzWlCVq6+VhIhn
sLNNwoxGYbZITfnvbARj0rnL2x1mrB5lg0hX8xiXbdAVHnVBnh15/zAx10DlvHhc
l2/uK3i9wLUg9p9VfXAqAwyHju5oUi03dS7Ocjlajhzt5bmgbIDQVIdbeaO5i1rL
UYt0sjArKZkb3dqQiq6NsmXRVB6DNHqrX5YBjogtehSgVztvKBTKfFm02g14iwv8
qUkZAMCPxEqOUQid7SkkgoBzBesuWLa9PAR6TuwkvAGdvJRXBehR0DCGQ5HQ8Xu8
81Tk+LO/5pK9G8GC4zsi42h7vUhKXUF/WS4paZMcSFMFVyujrY3/uxs7BJ0WWGoU
gCkMmhWsRRWbv8qfamq+9d/8UATj1lGhZFi29a3yoGorMcMgMVYV0Bp/iMxwW2w8
O0Utx380lsogCIIqOoMpaq/1fPXstK1odhQFAVUE8oUbI9dsBDLFMFoxxXMQcYWP
N5iSoH1qKZxWZAgkM63AGOyZys+208icwgR/DYCkea52OncIHmXckEiKe4RKnGuF
Btj0mFS9eldynusaN3gm4hQXPbtmh1SkddaVAYv6tF4nCA2hwHcwDNi0Eym9f0Eb
NGcbvuD82nt7++ywr6xqUVwhJCZkMddes5gSFXGZI3JaeSrbKhydnA141K8QEw5R
30SS9W2h/J3MFCoA7C8aAFjJHRroACNDR47XUAMhetwOJVj3XVj8MyQZisO82hJ0
zGXureTXHl7yDzCYBrgumecSY4CTaaGOwftbG8R65OpJ7d440hFJf+MeDx1KPTNg
Xr5YaiXm/4LbulMRjm+uIOEGzaQ8JGI0X4lagPQ4Ehs4cEcbhrmROxv04v0yJHdx
NdAxwQjyVGUcBuH+Ht/r6EN33WvxYp0KpO0oGBnGGmA6NtSpjhw2ct/LbKxSbQh5
8d/1pQ5XqvOwAPKlPvbO4cRSOH5thCRjSE5fxZ38Rq+wMPy9YDjmFc/D7/yA7EXk
UME8P5fJwFUGWOJPBaHzYl+6C6FogDjO5j/x3AQg08K0anazasxOFMYPJd5K3TQG
I1D1LXV6bK0j/DdASdYGp4VCx9AjenH7ykbkmLzQFvpn2w4KyooOFTMTwcY5yQOG
YL/AHVbIn1LAD4g4yPPJ9UtmgYSIgWuuCBntU2yCDrJHec8kS2dBo+4giSsQljdB
xddx9S+Ut781p2XcqmxeOg1Ve1kuxJB7BODqiRqWc6l72J+WTeHEbzwEhXU5Ny/9
ymRlbullFVxMiXqDmeOfrHCrzdngCMh0nzsmRxTMzm3UIYFnzT0Neh9/AiCWGgnc
4L28i8W6VYyf0ZmCLe3xqrUWzFnZsvGrz+eb80V+6dm+jZN5TIK5Mond1NJr/4n+
QtxOZZdPvbEQgH8immkwLlEd4NIFUUqzwDz6+aDItuzxoqT7CC7sFk4cf5uw4vpU
q5n/XFA/VTEk9oOPyJGGeCB6UYT4C2Y1En9CbMhAX3vlFd6fZRbLzxBlJrfqQViz
aHBuP+gVuZ/Ujr+tac3hDj9rU5PZVFkmHc1cClSwBlU7e2fD7qGzYfyhfWyh3kKV
Z2UG/VIlNNCSYI/umRf2D+uOpOMSXhykMNgzB7QUqu6O4jdOmeKL/1XJ76oAB/eW
jJ+9UttSF/whCa/AuY0T7N9Bbjd9yRlculckCtePC89O68aZ+wvEA+JEX3uI3L9P
2TL3QwSXN0vshK7Ux9jVIWsk2UWoyoSj5+P5TvaZs4HXoVu9ylynIxfWveJ+iMMq
SVIKjGvTui5vpLXHQ/2DMoAMVrXq6OZ7xHZI+T8BT02cPaOKD8sK+LK/psTsOP/+
y0WwEZIJwjMswCWU2dBGzRZdI1cbyj9BE7y9rv+oRA2NBdV90OJx/3s4Dh/b5iPV
fA1irCFHoKbIoql9VVQDGOWnIfyRzuzQC3MtXOIOAyucs89XQcmA8KIQnVINgTBL
N+v5Cjd2J5+tdQq+r4IvfgZ+Rx+mElZ2a0KDVY7Cp6k9Rl+3GnHe/yj0SKu1sZU/
XBRnBeGo1Rq11iQAU1bLl8Uzh7PPQPkmAPXLn2K8fSNyFaaD/A0y6YuQvbvptvzX
q871shltMK7kZxE1ffkz8Fa7p62DTf3uaTs40crM9qv6FwKLnG9+D8Xbh1e7TzDI
EF5vX30KB8y2TI5jfilJVDlTxOzrjq604XJvXl7iGc+ofl+iHmrj7vvD3bNr7sx5
GiPWEKUNgOtOgLQBqxIRj5wgE3hTUPLwqCEW9x6FBeZwQqqv/g7qbRscrIveDa4f
26C1IXQ5Kc7NMnQbGZbR1Llf9ntpv9OybgydPvvZTIig+O+Lw8eEQHcUtIFnoY3R
UTAMc4rF0u3lJgkdQAqtgSr1uBJ9MIoGmWiVRuzmtHxC4JN9lxNldoRAM8thr4M3
iER5lvcq2QakRjwSh50vPqp6AcR4SW12TXY8PjeeNhONg2NKdzHWfEzmvXsFG0RZ
ByxETkHjk13rYY+CK0cu8OdvVgu3LKXVAKfhxXdh/itpNEQTjg191om9NuvfaoWa
/caJFGXlgkE3QZ/r6FbJI83LoFsjVeWqwkYOS3Qlcik+UUmthKSezYzfiJbNPubF
qnuUTolXjXe91Zfxt3kHqc41plqidaGYGtaDlnS5uaZf2+drhc3fujjASFhHTkpL
zp2oXCe1eEkq5CVf6yPNtuuSypGj1WbsSOsVRTpIAwUZtQmfM0WuhSfzPK+RlbMA
boA4va2rh5AffbOwf4FxitgQvBg7r6zVvI7vISfT9qWyeLDXFUz3xrwx5EKRRq45
WNEedzcQYXbVUifqTqcTMDc/raMvEJ73qw9J36Tgjh4UPNESBy0X8oIiDardIkop
lgA+uI6bu8U6y1Hf9lkPVVz9meHbcPpDU1hxe6BjDqpY6Dyx5erzhVU88LG1QRuS
y5ivtEPWvVG6G5icGLnUTfSjPr17wtYq0BnuUmld0Flao07M4Dn6hz7AWi4tBFfb
oCOFgy3ffTxe2/woF2sosHQcJykwKVZS1bE8VO3rru7JViCRKGOg1wBPmd2oB5R4
P8FzdhjVlrmaic9hJDfOhdDgM8aRmwVr+OJUUS26QHcKKAyHnhYObLwnjX4GCzSb
vbo8RaiK9H/tRSdovOnMuTro7XWL3SFDlCdd9i4nF1YTqvif6fqQzIN7Bi6IYnY6
cfBZ0jQOkGoWwTfXYp+oN47C9R1W38P+q5u977HJNtAS/X7Pf5m/4J6RWJP7S9/A
dq2TthApjfpY1VTqJS6UYcPx7w2Z8NijBYrOHw3Vd7NHxS1G7KGAu9cla7TwzF7a
TMQnKIwSSCZfqxxRR7Krr/55FMEHRbguATrk427PshRDhsNPxaG/zaA22VJ51eSk
yA/WnHUmQZp3X/kofOn2jbK/1ESPsO9zdgtvXmkf5NTfCTfHKy5rEL7mceFlRfSx
+9FlSixcn2fTfIg1imUpSbYpq7k72nBvxftdPWBAv8slXqsp8CrCLPybidfSc3dV
bsOivzoIUa1Puy+o3g3NUVSAhzVMtxymhPJDrP+5l5kmxvqYdcpet6OCKqjm7oWj
jXtHjYN/zFl1CN1U/PQsHOCn9rvX/2LPco0RhcZlblFJo3xPvN1da0fMNgpjfv/E
qntAETTDZVoFpx9fs6YF6MxA3I4UGFrSvBDN6gYYNs1ysWnycEz8InJjk1k4nwMP
Ee9NIFjHQ6NU9teC/St92mZuFoBMrylZOz91A6tQ53PBXqGKxgYDDOPth6rcGpYj
o3MEzHY34y4jizc9jctWS3gwQViytOP41LaHMTdyuSE1LqxEHWID6Nl2PVeZFhlj
07ytCOEUPC5xSZHN5ZHamxwi379mXdx8NMeK4UqnhsJHbEBNcFallSoRv8ajbhtA
a34gtBtwNcjX2QSzZ4QG8W7Ev7WmX8inDMHaumUl2NeeCKzv8BxxS5W4YrZhXNh8
LL324Wqemj8BtSMiCOL7VMi7xCpluIMu/64UJOQo12JBazfrszY7WygKilFLwUiH
D7zanUwnbA4/Kmqw+W+t0AbqGONZiA7Ld+vFgyUnQbjOYc969f1+kErUEFDEsURM
BNiS0J9kHYbRW214jOI8hj7M4btHtZxFdtdZ8Uw4MQme72fCdnWXBAcJXn+pIhTF
3ndu0HqvgFbnVCOwYbf8PH977z3hGNzTwZK47fitZc8MWvWuPanUWP8sFarbmtFg
is7GzbWnrR58LRV3rynD0Qj9RTvUDg58wNwQJ4sXq4LNFwJe+eh0a2ZJ4PuMZl9h
lfvu6bbn8ic2Mj1z3nladBjRcJo40Pl84mGkviuBUzfGK+k3jJbV6ZI7DF5ADKN6
PGBJ1f73UYofXGqxbvFWUyMKcZJuYHD0ddjvEjCKORQIYHU50DWPQEq/v/KZHQK0
NTx0t+rFmG1UlbXiSzsaw+0B/96+hB/ZipeQ/vwvrqFS3uxemT2d2pvPKPKMTBmz
mtGwC6koAhAwfU5j9xe1X22Ad6m1A6FBNFPEH1u5NCScOHuMrOW2YVz2vWVAmkxD
FhLpyfSGgauCxB4s73w0KFCfFOOmsg1soYbjE6+nXX9Zi/SRYmMzoBH1ZgHgPABY
S2qEu136NvpVyExPcbPiZty8gFPbO5zrFgrccridpPrODuC+J3QKwvIhbaH3nbZ5
cqMSnUbuiBNpdJobe1Cv6TwGxD/GWm5ah/uJ6S5y88IXXzr7oaBEU3xm871d6P4Y
duEt8csbAvt8Y/XbkK/eC4pj9haYMelVFrue/uknVs0wbtPiSRCpq/ZMSsUEVyrM
81rl4vjjFKVWHg9sRwuNcSn/5Yx/dZIaDMrT+Zc+bV1ZQo+MP5eenzAUTVLxKBIq
qFAOpBNNDkE+/uCGjWthPvSVe5p+h8WunXYyAuvrkiBqc5FE0Zyb7rlip6NALqAr
Mkv7gu4qAEJ8fc/jxbffhstpxctweKozG3IpggMg26b8BqEmkfc9repK7/usf7bY
Ge8NZFwt92wR66On7GVFGOLRWiIcitvY/k0IDeNKwEHenLaL38Wvl9Vlq2kXL/Wg
A3iKNHAnJ/GsY8bXODpwd0vGKvTWoE604Umhf68rDt9bxv5xDP3H86RgeLgAXO1o
6QCIB3DQM/RPmUpIRe8qo0/2vgjx946RA0tEkhdyrlC0eXvJJRO3S+vS7BUl1Eq5
RgDsmG/aZ8n6tz4zX9gNIGrMvb+oR3Dmq526GaQc1OALMblg9vczhC3DivRSrURE
iqHUVx6ObEOFVNc034QNf2Km/UuPloPLjnZ7B7NTMRgqI0jBh5Dt74/7Qg3nkObr
b8iy75JqROvxtrTU1Oy1nLXdl2kICeH0+ZRYupmaIDodvDzMD8qqXmmP/mvdfdD6
LsggufLooOZ7UOdZS8I7krGIpxmEN6x/ufy/vDomVaakIHQx0zax4LiWkz7CgZq2
tIOqk9xs3HoBqJcMBjlZDhHYKNeFBcuA6a6fSY5Ia0+c93z2WAfjk3aLuVMDnlEy
LFZWHsBuZx3sb1NtSH7oUJoFcq9wKDoj99g4CUDbqkgqpMeQU+/sffduIxgqt0fY
T1pG5mWcSlOdG6hZzobpxeCyvyzty82VKXf+CfbSSbGbqVfu39w1IIfkWKHRqpp4
UGB9plq+02dorylal0/k+TX1CHak5MxNpfMUnkYV+XtrU5U8mcZBpswMsaFB6gqk
IXp3zSWDH05I239xshIiFsPzjihBLZwuTalxvJbLPDPmIBRtO1TTBb2lsCEMR/n/
hn4fN87ron6/wKARQeY9athy/nYSY99WmYk0OyZ9TNw0AeSRq/HUjRdRaccuFkCH
LkvetU7y/PHBDvuZPWba1OznNhZwX9S8UhiJOhypi5IWE8YLSjAs2lJy4J0xDzwO
UE+dAc1mFIvuBWLdvpnYZVBwuSRXTfsCrrARU/kEyC4QHf1Ihhrf9K2SssemTbVb
hJjxy6yxMpCdtKGsLd5FX08MyCIRcRtEypy4E8KP6Gosezjqaa7coJSu4z9uD2RA
Lx/TDAGCjRiJKOlON/nai/zkFnTbc2CMdqaj99g7m9Wcr7JPKCFxxuTitMvW9EBl
jENE/FmwuD5aTtJrc7cfFmEyl6Y93Q/AWdpLfiDINhJqYCXjZEDYKdufRomTmdlq
8ax7uhKqQLgfLpC0DzAhfuW+gZgyDm72xMl/WRBUesWfJ3t9SJbOG0AvGlC5bq+3
zYDIlWI8KR7dnPmhLuO9GVw22Leysu9v8MhHUuSa5YzjvhkvRaXW6Fl3sITh+bTd
083wY4PbWOgZYYFCfEfxs4IG5O+Ee+9jtqLSXc/zwrHV2JQDeLUNBTf+MfZ720sn
SqxPb9zMGrLZU+hp3s1LP/F7NJJEdhb18wnT0tl5XNuqO7MXkPRTmDarwTX8CU14
xWc2er7oGWt5Xg0+679aD2SW1/hvS+Ulo5kXXPkWKoFjZk0xz10VscjNEptKx50I
f+NpwM66Abd635SOa64Ra4EiDxx2Pcm9aelpSaOl1QMb2ngj+6WBVvSL41vq16Gq
X6GCWhDyLuaJeMk/JUxvpDGWcMWLSW6sOv1uTYKUhDW1HcBQQPFuWRirSp1Ige4Z
QBVZNOuWs9ZMCEB9rcRTMVnoC9Vj/F7wD5AxAYIAqQVDRELIuy79/sYjlTgi+jN7
keT2MN4T/6jLNGOggaHQBtTVGMoSIXQ2+v/o5VIjfaO1hOzOXa0eDTvQz1+9wn7d
qyWnYniYcmfcDwjd8p3JmMtgXgNjmr5a647qeV575sx7KtaB1xOtM3VcgQKcRjUc
rseYNCwDzVpQP25jj4bKuIcZoM9/NNLztNdnlrk38l9iPpTajENkaqNI+8w/i9Ls
bqiB58jitQpPlQhRcJRgUwLCKm6hpNyjzfzH5rTbcer1CXnFErAGaqLP26+4hPgh
tiXiRmjEtDzsu9afKkeH0ECzWDfuP4V9N1f6NCAggjLl+WuUk1Aye4NB1QKPeY9N
18DBNiGi026VwLRHXQtvbpONlraLOXYI0IaYG90m3PY5ilpLm7V8KdNmdQBn4bjc
PSIlnuf3S/ZrOf/OU0iQm1mfyniKzrvTIXkquLsL4HYqXXNCWVlcuR+ZfSwHTpKl
16cresjne36I3b1xi1D0iFGI1t06jfsRvXE83wnc2BntCNujZP1+pqUu+h7PloBb
ZsxlCDNNmhVaQofQ3PU+WCon6xFNlmTYWeWUtmMX3rxYvh3T36Ly7eQQ1s4M80BG
A9Y5J1mBgbo60LHxPuWWBo/ajwCkAZUjupttXPfjmR44qxNXxg8ZcGE6YVBRj/k0
RH6ckKSFeJGGXZ3GpsHmEhVxpFCDoCH6ucvvstgU92l7kkS52MDBYII9yyjR4nqu
2Sm5G7rSq48OUufoQ8jDd//RqjLczWs/UHIoXBa8PA2Flt4c0DY+xeqBWEkuLiCp
sRdWkxYee1JbA3j3TNc/HFFnGZ0BqG5KRl8/DOQ/nO5MeIK4yrWqCyMHhkrkfh3a
QXSHFwIeN+geJJjSkIqiOHWya+p1zTUmYq9ykSviLZp3RHWkOJvz1JnTq9A6D3GO
mT8XNSFuiscV19yoHvlzx0QssbYy8NqH3QRgsIIVBus4TOtjSTFKGxHDvJn8zRB3
OUez49ADuHs3aOq4Ud1xgA1L56pmX8DZQecP6jmcF4yCDNUSnKc9kPB1d+pL2/tD
ZqSwp94PA0qT+7XMQ0L/RyKblTlf4vtQhdIvJKxiynCWcEtV7B+gvztQ7EdC/NN4
07lcU/+xS6k9qTAqdItT0j+iTOYf6ts1X8cfoYJhfTGyOZeAJDlIToFFO/MWaXO7
mYEjyQu0NkyHfNbHD/4wdryuVVgxwOk1fnTuKtNX5bn6CaC9RYGwDBiIG/dpvA3U
g/pElqyOuqeOQY7FhYxUrU1u9Zs82bimAagh4BJNikUqCaslBn/AAnJK8WHN7Ylu
CzGu6pqILh029XZTMekuf1zGPKTbLtEtw+2LmsalWyXVjc1/pRBgVDAuXNBKYVtJ
Dk7ohqVOGHbByEloBN/LiGxxnQCblX4rnZhwOykdBWPbEGavTlXah9rVjVMMj35p
1fmaA3j576NqEI03hMrOhhFPvO0hzoOQbUn5ZQk361T8dHZ0D9PkKT/dv8VfW7aB
3QjCSdXCY/LZgJTqgm4vWOUKapgWX7/kGECP4m/BVMLP4sRmx76K2H66GF4dy5vk
TijpJESm34B0xgsF/8l7tT4w79Z5nlHvn+F/9hOhCp20r4b2N4blV1QaRcrIVmzM
rliIAEJ0/eQUSazQY6/kEntn90EFN6BN+fnJrxsfzXIw4zT9wK6wc6+gohD3S22k
ViJrRtvaj04Tvdt19kFT7eEU4jJEbldxmD1yz0u4xSPrJ5+dsFrueD0QDqzB2hld
NiRbjdozHMl9B7wIAPra12rzemF8WeJnHrxnFb2uEcf34fr91t9Wk6RKbVYSEo/9
DQtrBEv3yGvSzctUn8YwI1AVmEwUkKzSOE9vfpqoU8Um3qodJ/vZAL/ud56YkC70
6XQ4nR483CBm6HV0jC5cBhcL+Te0Hlxx0NtFlaX1N512INprDRyNF+Mt655yEg+n
MKPm+EwiEyUYh/tVQhJzMeLmoJR1z2e42O1XKvLQ7acGPp2ZBbmZdiDJ6CBbuD5a
mnhTJ5JqTGixCeJcOfrCrivHTiQd5Bkx568mU7gr3kUKcYcoTdXbLd67YUX/ZprP
ilmt0LcCj9Bx8rWfSKw9X4niOIDyl3bBzNkswdxU8cpSFetYFwipnDXZ0ZWyz2DN
HB/7TS4cAYPMbfMZJNWk/wdwyIC+qB8VZKksv9YwhdsSEARltpmBexMpPiyEEOXs
P44pyJbNDydAob1Sjyue8TjkZ2rMptTcxiZ52LXdl6zg0yMXiCPFp/IGSmfTEWte
YGz/9B/zhytkp+Na/5+G/PNNkMRF+0kfCMEi/77QpK9WqOka8LLiUu+VySadbeCw
AxnD2UdFDudbYs27BmuX+cj+xaifh0pOO6c4OZPHSjvno6aWsG7Xf7wuO0ppOUXY
mtk2e4BK7BFOOtD4AiyhoI2e2r9Crqi4iAEjPquYHcAwAsTBmKPTLC9mQYoTLqAh
nwDsMSpacbEYR+JDMRO6COSVE55s22h62YWso/mMZNpcWiY/1bYLCh3MuqGZx8uz
6t3pRwgfsv3FbZuQRkebRXTljYamw/sKKfT15Mr1CAOII8Hx2m84ZkPZUV5VSJqv
Vil46HwIo5B7m3v/7qXJvsMCYnE0sYP4tWelzMXfFRRqdi2P4dzVX1oKGsaL4vHg
E/GoRt5HH+loPynQ/ZN0/Zla7GRFiGDIy3sLh+WiESlrSq1UYhh2IKqF/AcugH9f
C4MZHPHq9AMR7BHV2tH4VdfSVIrjLGyWan/2wo9rIALIJPo//9PPnvJ8+moTRyFC
XzChCEMCdWmIMz0ZgvCunVTZdJmnEXGLoYUjq352djtx7DOLd5O+yv5N6hYE6Brt
0kxJpaz6svKT5TXFdjYUD3pP+Roa4l6pj7cvldn6g+4wyKDHknVQdLOrXciB2h8p
dOJFsX/HI8Q/cuAo2DZrvlNgcUNllSdkh1ZAUMFPgC8V9+9DYbKDU3d2QvZX3OcA
d3w3qYrO6Yh9ADK0R43GKJGz+a2t4iEP2u5zmWExN15BuibCy8YoYnCGtxwLGbNi
y3Yz8ZxIY6zNasaNBcBDl+L2jbttPblMVMAPkxrkGWb2vPj3BfY0/H5bmGkKfKbi
pG8VLPcF+yNQiZY1UsejcspnZAUIkL2n6aRabxBMerhVniPh9HaEt/d+Z/+roq1G
lKV2odE30W1DRUOZxIwJYbt2ONeohjTjbKp+eeQvOraAME8rYsmI8oGqbMSI/Z5R
DA2i3JCehDNAElqW2jcYetoxtcX5XpYWcwZopR+L+aF+BV8fj8dfygrJfP/9CmM+
PocPSxGqZ4AcV7h11F+vNtL+PAqV4Ck1xBlUm94DoCDkR39hVtE9WQv31d82dwRf
2oVad6T1uUKe/JPT22if4ijbE/dVsz94heDqZzariwCBGCCE5mZNtAdlA+r4vu3E
kLqag+Z82nZ/5KZVGOard+U3ZkgZMTOwuxZWUo3HmZad6FtB/O7jGBE+EAEaXu4N
1mkqxYJIiKd12LMv9Uu7/gw5pqiH8mfBTXQe2zZyHwkZFNeMydZSr2zNbQphwVum
QHY5u9ygVuvfi/x57O4dvO7VPN5St3E2AShee/fIcgJUZSh5PwqKktRt3ZymW0jx
sLjECtsGTR5Bw3tLZbk5hKUPwL89VpuWNW0v0S2cUS8be7jtietuxNC8lfygVXeg
FX7TNskUZS050UBhRwFk+PhIXWEHop+K0mSrN1UUOUQ68SuyEmbOvtTNbD0zqOSf
1P+BVzACNwh8XGx0MdS4uXco69679S8D139YX8JZ0U7JA4pH8/vU+c0c0aDaZyEf
oKGfEou1UUtduUq68mr78UxzJnwQY9Kys2n/kDL4X/I/QL8ss3ouMVBgcaVjV1gM
QYOMDv4c1jZZqJ4BDFqiJr1GhCLflyf5liqz3uF6n4pj3Vxg97HOUUHCtgbYZblt
mWN34qMYTsVVYs74gQOkHGXhj1e8SljGk28SuZOI2Oc4yBPBU44V53XU3gn6nQ/w
Z791Tc9ezTHl04Zb3KXI6OUnLXJ269YJXq7jCxdniOoGTcQo+CDDQ7yXlJTddTd2
Af3UbSvp34yj+1XL32CQoP564ftjPiFmnPhV4+dSwNYxiAR4OMHP7I+mwB6wjQbw
JfJ3yUe/889NRuPpgw0rgANKiq4OPPbS9MOYd/dwntWEZtHzr698gpz5kfvGr0wD
GZv3OBCwUn5kibEzX6ZS7mFjDh32nzfziNam5+pkUE1+RfMxGqVtjSVGS+pVCo38
PVi7JA8EdRvw8MlsBm8oOBUlgV3g6JBJMomQGl0Sms6bipSptbUobE/TMGF+sOZI
hvlR6eamiso1SxBnmTJbsOrPZf5SIKPfcW94VevD6zXnGTxzWkb6wZSicSM9i667
T2nqJbo3HyGG8dEvvW7KMcWmBJvVFPFSfqWDm7L9Vgj6DMUAUtJ9ETI59omMSGT7
ZoOtTlspNm3Udk2oLroCIbrIYQ5g5vcIb859oabu38l//DTxQHBh9xJFgkKms+h4
PWdnHhw/aGPKWU4Fwh9TsccL1ymL3VOVokFx0JAOjEvsmhAKwnDZa9tjKDsvr2jr
cZx9mPMdz9Hf6w6YR1fc2y2xWrZl40w2I9tHnFfQlyMbyxFQB9vvaoyr9+zzi99j
pu93El86Fc+6NEAsBCAqpb14eG9YLi1d6ecGxTfYeew1k4ZyJkhwASsS2u0kkhQs
IRXup5UmAjukoyaSbpjARMQwUzKrVM7I1ywK+tg+NnObdvLxQmP/noTPgsEdks5D
kcOQTLN+SK2JQPBroRly0YtWga1sXuyNzAsxSQAz5j1GHKewB7IOLJKtyelLoauM
cXEiNb+2Oq3sJ8IzNpCRfv1SIychm/hkyLIhQfWdML0I8wGqVpuAft5ZAqWA7CU0
zK8RHlX6YoI85dN5mptlUy+KdWVPow0fomFEa8PopqKNyGaoNnnJ6xnHvF0GwKnQ
lS1CvyrO6w2l/zHqQa9DG40e1LjFfKRBCzOpNu3TUatdkGR7m0B284TD6yOqXM8J
9F7U0tzor7u6Fa7IZqMH79fFMB4ldsMoBwbLjTL7fU6uXMlu0iwRngbddlEPG8P+
ZvEs6xavO5THnR8rvqPKO7tIZF9tM6CHuvJ7Y1H4Psmk9igv8jOjsRLSKsqeoSl7
D+CN9W2jI9GknXk9oaeL1r4yTF5ULPtb4k3a4ovZe9I7qCLVFo/rE6eSg8EEhXyE
X7f/+pBEzdXM99Wad0D8zSl0VKlRxGpBp9cPXX/OA473H1xSqzOXM7UueQcDRI1T
KyolLqt2ozxo6mmloisXDcN8jdFquVKSzSPihwuzFxoclb4GalyT8hWPvqSotpQb
cUatSt61suqFNC8mXbJgJAePJNIRNyzNIVkbOPL76cMfK1IlAaSw3dhY9YXV84f9
TjT2upQjH26TSZ7sUQXbteLrNM+/3wYDAd1HIP6cEV1N/PQtFnAAyqVAsEbTR+TQ
sSdrHE4JF5wo8l6XXqDSqpm1Ts21lZVkLdZUOpmOtU07KEcwo5oWhq+ETyfxo+ZX
2IUvJY4tUFyEU12/lcrljt8XwvfzULRRws6bTot1VYam8EeZVNADlxLgJlGCFFGb
b+jR7HKW57XAsmzuXVuGikFd8YUwgQm6w2/7dxsbaRUw+wVr079BfkB4mzpPVe3+
0HFQCAZOVM+42ljTskj7F0z4Ok0BrsEBdZ2P7vqusm+5Er1CCEY1KX+pl+dnD2ZR
ZpDlGbvSDcD3hV0F7t6mGa6NyhCn8lHfojPic2l+j9SX02pGmSCZMscV6/0XGw+E
Vf9MXhM7t5xtDJGIIe2c1wN9Y5CtFvXAtl1l2hOk1bJiHLBgZlEpHKUaKk+G4tEx
fGppCdfGF2PC9AekQaSNPpt9GHLs/Rfms0H/cO9Dc7xts45lZEvdDYJ76Up1sVlf
gLMRKnLRZujMBs5gHowT7pZ+nNXFNszBuphgRGUhYTjqGVrUe9LopVxECxKJ5kpp
19FaEoNSy6mNZQIUdQ2iGGJZ/onuepp1C8hLLHml6lJwbFu7YXFFWvaKg5GuD4Ma
mNbwl15nrMX+bGkIjL77UFgTnb8+d1wFSLmaI/hh9Ue0F5qD8nj7kZgQjSUm1Ojf
HrMScrCf99ImYiQPdjHCwkopVt2ydQ3pQQiE5xdhOgXuo25KILx1g7WGXKFq37Nn
wDHrtNSf5+niGbWNSKn1EWaX7/5FOqP/gFX8rsPv1TNqxr63PKK1Vefjt6xe3jkO
Hz9Ny0IACt6DR8VSLhuHWxykydkaeQCrvGI43Mfc1Gkhbn+YY0yc3OW701W2QqCp
dlYFxF+ZWQgaSpthgzqr1bsvGvmKhjtqTQrA6ovOqJWapvMiV3DSW9CDWwIkNrBo
2URYgXzAjYfMOQ/70PNIGnguXIcojfT6vW7QEdsdVrjMqXWV0lOVq5JjzbZroK1l
zac02pCj090iAwKm+jaoeEo1W5buogBy4vTf4kgt8nzQIup6whGQFfo7x8+vPRz8
+oVa6Auu2x1pEqRHhmPlWxqB/hqK+AIBM618/1E7rRFTghjo/fIZWF+1RMv26nmi
im4XTdcinAkCHhxf7PodELaFs6cYILvwzioFyK3OmCjenrsmJW84jMqW3Lb9E/ZP
arvw/BpYcp+dcd0tcvsgHUe0CcdoIAzAqxGgw2z3/wU2IqlQfwKhJ7Ob4EkOO3/W
oBNPxg20Xq6/2+9pQ4B6ajTN+FXK8Nyoj6UCwdFTtjm4UZyu1IY2mxbdxgsguJ52
ns74KhM9+5xnYxVrlSI9lLdLaXQyL2Q9wrFLi0+cONOZwEBNm9SKx+FiEKBiLVA3
cvO6tC1u6Tv/xt8r2KWVHzZeF4O1YvBZIGfvOYIRygyvzMKDSkNrNNYgRJa5e4p9
JdGK3mXaB37cXAlLOe6tYH14FHZElGouMB8b1A1X44X3iR/gNcvqW8JQvut82lxZ
7LwAymQuM4ExOYPvtIYMMi/pnQP1znCJFsIWDb2IGdb8QT8ICH1MYDIV07AUKDV7
z/Ma+hh0UXpDU+2ITTGEM8DepnSnQFfY0Fof5Qs/0x4qQ4wphILtfyF3Sz/MBVj5
CY3vzKuelMY6cI2mpWF/3GARbVFAHgGm6D7g8AaODdvEFJAEJnDBjucUgMajUdoy
PVdBg/CGz66s5YzGxGBrruqKzQ0hdnWq/1MkSC1c9DD+Mt47EUi5piDvkqMUYERe
7qiQuqDJ0Dp/sxqXU5/Pis92eQLdmvSTRscvRqZcrJnCcxbIcx1HIAgNKqPSoa7Z
4iVcVcdV9faNTzPRPayqJDCl2h6XkXytGPRdJzPb2sSJuo9n/lkBWsYOmQmtO1cy
z/RaNuHDAi3mcNgsJpEKpNCfzz2WcHZfjtfNFtX82qctBo84HlJnAtc/v4X+9V6C
KwlksgHexTVLw19DxOl+HIkF8pTIVNESzWUwwYV/8mT0qnO/TEJ5PgXCfbu86i3d
xhWbnjnC5JjLhUPzUcec+MTUMDSDNWjsnrQ9pk1EoDCsyQQInrDgdkvXjKcewFtu
yac/SzHdMBut22UNKOzraeSZ8uLEYDfC+0pOccruo8G/cKwN21q3FgFvMAxpzHiH
p1O01z7RQOBv2B4uIppXdzKRt/6d9Qwg1CnUnJ6x8qPdgHCP2zYQtcsp48IGAHvc
MbdeJUIlDUpf/DAFhHISaFotzQDmV8OaoU3b9KjW7WA6xCzhMG8XTnbNk1OTkOXx
79ewUCVWLGiKAwLbzk+k+xssgjJDeSFvreRzZFOPHS4DPS9atUKmMy2AzRM5cUb9
WCZ2Qeb6itHkOvgn0ItRYf15R0jhhSE1LO+PyR5V3PdyTCtl/N2Ah9FytJJBY1y9
KvVYiUf1ZuuWHi2bhHEQRoBXpHnGQZoSNvsbavX0IelI7hq5MSzBnTSbdeShTm1o
u5YhI3gMEbEZ8EIAN0voEWhBGaQn1AlJ+xn73xlDkt97iNWQQ8EP9LZdyeEM0lUY
FXP+aJ29xe3yzq74chkZeAcZy9R7ZD0SuU0gBmjfjU161f9XuxbYCjEEHAf1p1iR
9RIUOHrX1CVFx0Dt5k9E5erChPMfJB5cte4aK8IYLJVaAdQcxANXogl2GsaxHO6n
hDh4zVCNZRnwL+s/AK0lRUiJu7VN0cSco8S49XDDrcCQkbqxKEqC1G6JN87dLGDf
glF0/Y7xdRFpzad/nVBXRLHFh8qgV3U/p/t2wlxBmdq6t0OG5upHnfZwhqqKDjXW
1ZDwzMjC+08dRuDWzpnA7G49EfNyMcrrlzlvDlZ4gfbJFJ25+bmdWYRedWbF9ltI
M9mUFHNJzy1wYcedUeqzO5RWqrfzlRLG3BbCfi+qlkLWqmYHxK12C77gC23qj0PU
DQ7DyJecjtn0ZqcAcuVXPX2Ej6jVGtpu1i+97VebR5GZGQxfyty30jI5/ED5R28r
03hLu3ZkSSm+54Jw8UqIRa2c46N2IGrN4fdLz1m4evLl9mj40Ux5FaCP424QJFLl
qZUNYnWILT01NCF8hkrHAMRE2QznD+PbAg1r2OyPZch50wBBNyFlK7NdoIK/ybe+
uwWfCJw90FnpBhnqY69eMwBEuXYrvBLekDrA+ShNu2HwWtszMxPEjvN+xa6Z771Z
HyAK4GEYRBArv/3crg2ISpGlFtHbiZZQo17OJhGehB8E8fqYOZ72vMbOAtm5hsS3
mpj+KfaEcfIQgfVzgJ3zGHgG6Q8//UB/FgZMZfLocmqbAHLn4Qb3AbuwguTv31LB
Z9h8YKQDttrgGO4rKHeDsa4LkMpp1kvVyKJpX89hDMo1++ANKh3Aq2dtydCRaiqz
EmvlroyOiucC+ZAgql9Xn0YS+L4xzsjgGHKhCVqn93uHcdqXCyVyookHbiRN9TmP
kaVhrLFcGWmcfxcchtluvTr4jxR9/3DAD4hMFB9hJXDIajGh6076ZiObRL7igCEr
RT498zHFpx3Vc5UR6pQ4tO+hbda/fYSMcNv7XPKcA09JftAlsBFTo7CgmPMQRfa0
v2x2eDDZ2+Nah8fc3xQn719Aiar02ub8jLPNAcu14Z/AeleOMYT6diFXz1yVHTYl
9Xsd4JCdZc+KRAiWIFKANOXfINf1v6BRT7/Gui1emBWFRGLFeCXmK2BYV1tvLB9D
5vHJVEUJ9pec2CN2Kl32YLskbm/b/g/lbtCv+bWDQO05J0TClvMYwarSREE1fxeY
d6xogcik8TYEVgyBxgYJLTN1jpkpINPBf5jL70149wId1fkn9aW3HkjAHpi2arAX
BTU01G9g0tbTR8tbQ2jr/fBTihcUcOfgCm5dlbyn3vP3lT1Q8+mRFPfS/Hxd9z/C
4dfiDBb0r22PBRi62jhszTXH4lBeJ3tnOMushysAQ+n6PwIplNpfjTm8uzQoBKZX
t9L0vtUrlLNA3c+eeSkUZXJ7EYDRlk4RLZv91vuuwH+tnu4j3Bls3BQAZaBGv45N
E5zsN1d0yMn+BCa4JG0dGWmZhHxXnpA/QizFXcle0E7m4V9WsRC2IhJ8znC3d6XZ
HtvFMZTlOjczYRTuTb7JV47HerkxSUs97x4mf2fe8JUChAF0YJraxqJQ0sChW6qg
anlXqvu/MoCFMICjta9cwEL2uKSdR/hLtKQvKie8poFdRDaJfdwU6hjVxD193FVg
lCkP9093sCiACu3CMWTo3K8PNv2bd1soL//LgcJnU8QovcHdLDaXBX3+uOmLwSs9
N0KgJJUx8Rz71NGI9/lg0D3vysMNG36kZK+axXWAeKtDquvk6QOiYc7zZlh3JJzt
+ahk01PVCZ2ahXlKIWR0YTJ8DBrr9igLi58Tw5+JyUyj2bpbhqeFkussVwnIZWSU
91hvamRjpbGjUofYgKqMw4lX+fmWH+o8kaSOrfvlt/99KrBaytshJttE9vF1/wsS
4iFWayt5MrzQaGkaBiBDZ/1gRQXomj2guwirz/x5TTe9K+m0C/5n1lRIV1M/BoXQ
Eow3nzGK0MobwCMGwqT9v4cEeuxuaX5yFOw++jPVKdVmy462vpfc1jbjYLj9/CZx
GROLv7xG9A1dNNkWP2JxBVZOLZlI+YMtuoFivwgVlLTVKqa6nCec3yBrrlvnxT4G
RqlqQcFti5sMjjP1ORNN1/mY0kffwTsSwypdUKg4tzi1crT8MEvfrFk78pcoxlpK
Mn9zFarLxB00yCyPcmtvdds/EqzrIUs8JnPtgE4SDPGpNaqgwNx1Bl1qpiowHwKk
WBVmTHmPD3hyYNwr8RZ33siYW5gQ1hCGXvvXzBLXh9CGxLT47hqleq3H0o5a3TJF
ZXMAWZf34BVwBnzxjgEAI3y/2MWb1l9c5Iv0mCFemjfLv2LF4xTrMHnxbY+zepyX
4zYBDgUBEoATPq31yCNU0rCrFfmx8azXJ6uqc8PjfLIE8riRfNfMlgO4bGFufRBY
2DpGMAWh9Fg+bHMe9k11T8s7yXhSsd6VuiW/ub9ql/OgfaPvpLsXNFWdOobdeEde
+AZ7exFtROyktV/MVqb9DDQt4OhFYVfNJvBvRyzJm1ziEsDc8IOy9FseFEI8HenH
iTLhOXTXawc+5GdWkoni2F2ZaR4k06JipjPzd7XU5m0bvjyCitrvqvS2HUpyTx6D
nugHjqDOYPgEadrjNjJuqDG3rqqEwyTeHZovM1cuZfqEFSDpfkso660y45pcELYA
tkDyrqLK0swwdndRlCK44ksdbY1BD12wXR8aJdz/WPEq7zEsCLGIKnl+aYF1HnBE
cIqm1MhXPCvrr+eHs1SNQXOfu5/NjkLnvywt/WV65vxJuz1K1wZwBFVeAyNbUSD3
LvrIXr4Xl36EE7DVui/MYxqpBvwrWedwcldPEF0BSC48NoNJm175N7a9LB8rC1cI
JiaM/XrF8IBVxZfmaE5H3hXTUicIjKuv1oI7DR4uaPQpeJfH/lVCpwEX5XJc6bg5
PubaLjOLq0cYPWMRNFy+mxlNe2t+XtTtvvFWW1+ahuOYihdC0GgHTIpsJaiknhhD
A+m/dRFiWbwevn+9i/CEJ66NupcenNWxr9cDbmojx19KYjbxW/v2U07qPKXe+CLP
aqUse9cZ/sr02rmoRqasnw0wmDhZlrUHCVkkdTaQl+ruwnKg8K7TCa8VDXLy4GL9
eUjirwnINVzZTiKzecOXYcGAQg/eOy3qjH/3r5DhVs0WYfHLpo0jRuZsFkNAYnum
JIXT7EoAhjxCrBMhgW4gfDbNbRwQ7JbTmFPEDjAIM0ZkPLQtZjA3IgcS+RjZHDTt
GGy26xnuUGxdbNfwTX4riQHYpHd5owVKUX28VVJzyWFWJJtPye3HrjpAmEqXcXM1
yN9p1POHZQF8ogP8IqxwhxNFoKmSo4Zgu9UuSfllARbzbNxZktwoJheZ7+TVFaSE
Pvo7jdTuaFx5g4I+abdv4s6TxFTnL40m7ZQMlMvoLKGLYHeoazCl8uK5geQbfoAL
xVZrobSQ1s3IXB2pUn1z4/KERJePSzVVIIR34XCX+ihMprOhJImT7fcww/PXIWps
vSUBNGJhACe2gtMqVgtkm1bzZwDNVzRRJpi0NYFamXhF5cjgOUUi84UsiI8ELLjv
djgpc21Lvf1YFjERazRFxr3obnovULinJf6kgC7W2O2r2pJuRFQp1CWB3uYPlMV0
p9Ae8LWyHPymh6AihVMGjWWN1dl4Y+Gpe+yF8kK2QqKLUaGowy5CYG1N4j1iQcuh
pOUzMZQ8rQiV9JH/Z/Y0FQUWd/NMkI6VYvvxvwATsHmUvdulx5e5/5eKzT8zbu5Y
oBxcIdkR6xASyk3J5gjGO8eAoX92a3IsPI/q554/eEDVifviyHUyT4MkqOIARXIt
vgIgwWv3pHM36Dr3l1KclDVa+CNlh3Jfsfka3PJP/tKdvpmF36xdROh/EHOTzCRG
pmwLNEku3SOra6hHZ7/wnDpFUEM5Kp/6mcse0SvrbzcAG7lG9q1wAhOznAuS+nqb
JzUqQyYwzpkloFyYV0F+29ZboF8fYgJVvLPXsi9l37gG9EljqEhWEzeuwYC4tBjj
P1kbJ3qgUv5kag39g83NipHglCvu4hTtfDlF9RvLTcrZiHAHMgTGAtE3k19X/iqg
7ajZKf3vLmZ2VFN71tXt5I8Qx5t//AHrjcB2J7vUOfhsj3skr4+NrrIO5CoEJZQW
+NjVMsBTUEyZxSw2PVYyTjNqi2V6nbbRyrmzoeiRRu4EZgP40vT5pGrmiUYwXLdM
YaqKsDDRz4ES0x/oE1lyPBab3HiWKGyIXlJRBOkNbPz3yUbfN1rcqAXkjj/lQ2SX
2R+RKWyTZ/h1CbL51Pa0uNptBSiR+1IE9RL2G2AiruDx04yWBe/swMsKYCnN4a1p
YTGN/frcq7qEJempA2BCXMDhfBBDLmhxb+5HCh/E07mOxWj3PsQJX1R9aJY2bigr
O3gwKhQ21euvM6M9AZ5oSA12ZxkEbh8Ft051GeIwQKlepS4Z+dZ63B8O4wzBY8AR
QXBr1OFbNuBqy18DdI/5pOihRLS+qXsUO1kcpPgGKwJ6YgTgZ+VSog2uD9CFjMA0
D3nFwEylcIFcHq4XKX8DQiNG6ZvkdewT8Z6pUj4gsRfGzS47Jex4DGEkigCRbOTC
yXtI6l8RlNcvit3z/MG+9zgYAYuhEiqTDQ1eOvyS5u4k6uvlR3l841bEhYE5aDCu
hUm3NWysm16phus7+x4oiaZ091FOSBojKY8MPadwaJm0+/rMNrnzTazp4JtUUMTC
1CRocU4ZT5cRJRQcqz7FkyFVs+H2X+xpOgZfg+h4nLsrWIdT5QxZLEgcC5xGtaEw
lgt9rF+b+WwliIDvK76ar+gX/2xRcwjeFSuANF4q+ZXsfbJf9R8gX7QbkhPH72ej
ZO69xmiqUMLnn+WWuvY16h4gcb6QtwzbmS2nEEdQHK6a3xXEkwxsi3i1jxrVYJZv
bOSwNSod1phWuA3ddUbAETJnFz7+3TyWXy4o8RST4aAkhRfbTo97xGntijKRJrwA
dFLagRBYl7OqiIvcsBs2L2kE9Pkwzi3XPVchcy0e570q2ntz4aFvyJUPyc+0Lss/
f1SUEEO2Nd7Rjns/dxHosiG1z4m4lcTiJ9VJfSuqk5TvkytV7kbyahFXCcv47GoM
/9Fb1Md92wLjluGIVJ++cmCsAuppT+xJTPlF1vWXsUggcdPqgeFpXtMwoSdhCJdk
CARM3WjbK/Nn3k7TujKJvhqiSlKMK+cliAWFuVMyz1NzzDge4Hs9xikx5s33KenL
TYr6UY5LI7+PZtuhS/v7ak4lmu2S8J8ThtnjajXJQS3QDiRot3s50bBsn7AUQi+4
/7UkpKD+ncBJYUygoqK0ug43kRZ2wqLIpqe7Lv8OvbrRlS7mKnA4DAsemEhEn6GN
g+f08emzsz1t6X/vyqBUOwf2pd+gdw+snqiL0U/jEQxizU4ASpm33j2jXtw+xe5D
M7NbWcYIuSK3kQTepW6Tfk3hwTcjUc9paLi47yqtbEtPfCZSiEAk8QLsijIKjWTg
jEyv9feHoKbA2X+nVTxcwXLYtfdmy5jDGxgxhQQn0Me4Us0CYqECmDdamnx1lCp/
Fg7wF34xE6zDm6OQgqFeUHgv+5WjuA8utyIIVX+8Whad4HAPeXAZtNwRFe4rbYI7
0Dnf6PWslH4PtO+QbU4c0Hp6Rzpo6/nr8VehPGcUjboNZlwtQAj9AQeAY6BdmMjA
NGQFl9lxscYkjoZgBF1dL6BKuPAQktxFAA1WlsBM2eNc8MKofsE+ckD++BBaQF7Q
Sh4/0MXfjKtyBzVikS1nBfg3zbz9O7RcYvSLRjgjV1hswkmmhF4P0UcaLlPThKxy
y3noK/wp4cxVowbWRN9M1ECIxbXQUXurJk4QR1XcchuLRdNOimBocaYDHOu/lsB5
zL+NePqEm0SqFjpDQoY4fFsGi1iUjQZN4jlahR99RjVQ12d9OHZS2eD5T02rRHk7
2EBgngK9sZl2oTvMy8MRrLCDuCMU0rP6IEdMAF1Jz1fokmCaUvE9KSRnUeWOy4gJ
17rCJQ2kYjm12OWexmg4/FeH5RsrAIyr2D/oji0BlbnOAUwTktzmWT0mDcK4VX+l
gjIQVRY0626EIzxyU7vtYRleU8aMy4BNADVxhWd3K5cEipYBGKj1Qse0goRS0BXL
dTBdp6bfVRgc+vPQmw280w4sbWHx3bXhJAfcXDHCNYszi5LZxQMyGKp0oZN1y2Vy
cbDHTcfVLkzKcOFbgA6D2A+KE5vMRDi2Av5lnRdCqD2ymgiHE0t6KffgE7axNec7
bmsCA8OiN8wBLnysXz2E7M4piE1TqEzpoP9s9s2459sUpTAb8YHmr5rsAAWudZfo
VKZQM2Y7OmIMYD+53EGB2qJO7fyw3JxyYfKdFyZdFTYPYsW8km1LDZSG6SKpIlKK
iBsLRb3+XcjISmBiS3uRZXfd85wXJdxS5q6IqAntePDtiy2J4mzCLwGOlKSG+JK8
tlgP/oo+CMvxnPeRBoa5L2GCQXs9+RDK2MlF3WdWkJ03aerkZoMuvh628LA5tWkx
9xXdZ/j9yOIRQf/6CAfJ2HpWI5Sc7khx0bvhJxAN/mxC4bT92BLtL8db640z1M8O
d84Td9p9xQ0rOUZpyDJpTXYma3prmjipTkCtpRaeE8OxJxzQs5PLQSM4PeXj5aCz
3/3LMgzzFT+oR+vAa0uemy6hzf1pkThI3vR1HMMaxjTKomhmuNp1/KNGtpg9jaA6
DZNEWnVcghfj3c7BfeAS0ZUWVAXur+Z8K+xpqOLH+HEnxR3H0tFEhy0MdYy1A6zL
orHh12vBodsMoemJygd3eMjgcOCisZn36yTb+Y+PeS1YQSS0T6+TnnlDDYSaZ26+
dxkfxbcrv0PQxsGA3UX2nKxZF+bOR98cNa3KCcJmsndXd6fEhjre06BjRZKD+e9v
uPLtZq/SKZ4nrni501Wc9Wy/o9DHwrAcQZidYHNeh+2Tk6Qgul9CQxiozl4Zz0pn
xUX45DsfkqXnSZZ9BXXZ2M9YaxRJm+zqRblqT61TQsrVbsdryU60FB6Rhmxzg507
g4RH1aZ7pKJsJBn7syuNnPMbvZ9CxTgGX016WlO6HtGPc2Gw8TM28jP+Ej4E+TQJ
w7xBZVy3FzyGGEjQMrhHPdvsDbfGKz/t5xjJ1ARloetWAKcEn81EwG9bVEHzhOK0
1LMza2Y1NVFVQIfh2UZoQ7pqtl+177MSXQwCprT+MAUKoL90KbNe1i7RiCZx7/my
3Igg+yEpgDhIZAY7V0gxmgvbNt4A46mUJfe19j9wQmCAC9mJ971fg8OWr2XViRip
95LHdkMlQb+P+vXYHDCWCuCc5EeciXyxe0XoVga8Y6B9Y0JRkYYw4SdE1gzpBD3X
cErgNwUH4SPhg1BEZm157B2Wch1L0+ranTMQFozGiLRhOwKla0r1ildMLuLSUNUg
nKMrarDhYkl8LCvyxnu/hs5/wppNAN12xDTyRxxMBAvJbWCvIqfIhWKG8abUWSCo
ATyC/S9lXkqxN0Nptd6AP2ODBj/SLZUeGga/9mQlMbeFkaWxL/jBD+1S/w9kuuEz
ipvowLoaEGmwLUsUI0D3YJcGpJRVrIPgAw4n8iYg/kn2T0JHmDOlB+ajLHtvLreF
Ftt2HGeNujJdUsN4qFs15NfPwsETFlxVbgmcpYzaSxTxkTiU0OXsJr3fYWempkKh
PMFj/Kbx8nRpnFt8H4njjOV1/EkH7O2gwXFMzF+bhDwa+ecW4d0gWUFHV9Kpn4av
9NQgH9IhhW2hzFF/N5N1Jlu8L8+Fpoef/kGiaP3WaesE80zmJhaFxGjJHpKhXcUG
oL18LSxdNYOthxRIXc8pbfq7fVmwgdhfnNk3wlHwCiU=
`pragma protect end_protected
