// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D8bOKM6D8dLEeYTdIj7OWxtz6Ud7WCkzlIKXJLg156why3dF6iN8v7QGnatR70gA
gd2/GEgD5upuU3iyhXoVosxLR0KD9nldaDwnNIGVZq/riWLzrkA032Un+4G6wn/g
4kcAF4vcbMhoF7bOGfnuZ/kRN7dRXqO0ZXs61dcMRoc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 324752)
6XALmH0MNkcYFXbmtizgqKkmgm/212uF6k39uh4Utd/Xu0o30oYRJxIfJRJQ0YNG
Y9s+ndiss/t0gEPNt4MdMjhB8DdFwo0TR18TY58d2vT+ttUPS9utdpKxGAlL7QLF
NEjqkTGvV50SJmxpkouyMwBh2NUKQDDd1YkZrCuVp0Wk0nC8+OOPSkxBcPifzTHz
RqQgDLzG/IZhmwjKKJkfrQmLO+qFb6cIqpmhCJTDJWJoIRGgEAsYpcG/oAarI4OJ
yuoRZX1/PjgARFDKrWW5KF7NENcbe0Ng9BtjkevJxwS1MqEEjs2QvbI8OUeAejHp
qQfb1+WyTNcT4D+oqygsjimemLsJ7N2OSm81tJTL/ECLnIwUlyjVBWTR8wbBlVn3
Rsi+VJs66fMPTzcwusuCiruDTPg3m4b2EYY1KVGFiM+o06Xcq87FjTsEZhHfou3O
EYlaAS40ls53FHXrB58lW0QQ8ijuV24Ce78vY/I0r6z5Ps7qkecFq3ER6VS4mkBL
auu4XoLL59XomnPhxX2O26r6iQGpCyTopqya/xNqFpnlKAqQqh5YVHg8+vd2VnbC
Ebc78xmQkgp0uiyW7sqrixp7kmiHjAFb4zaYgOs5UERM+YXkpIP7sdElW5asmbf2
F5DqYBH/2aQ09eP9g1QS0np6QHbNZGjfuoQ9bqDUzZBxL1Cr3ZdLQAUyZ8TC5RPQ
OKKT4L4lo7zlfcIw55teVHQiT3bL9fSaXK7QucjBsfQdt9TGFct7zWsEh/W1JYf0
jMWLsqhMhK5RZjzKFZPjVKumz4YwxYgvDk/wk1+8jvUv5ZPGPGSy1l/SmVkw1x/M
HzX3eYqGw9zWFoutXwJ+wHHtJQLReGeWmsCR9p13k1c2oBS/io3mHB5klZ7t2S42
uEOFoKKoCfo0HaFsjTqGaqGbJYdCRHBUQDY6moyoaCdaWoX4KuGVZoUOF6bbwUmL
kt8GXk6DPLtjA53zRwgFzVMsQtXb09uIEt4UiRwTRDs3g+mTJiWeBS5pnijXNmZv
ZCNp9YpgehNevcenbxYnc/u79z61BZAXWkxz1GG+hK19OmqLfl8mIKAzR1cAyYie
4nmvZeZUN1teaq7p+T7VqXYpmGDHLBU8G9eXjlw0/z+ITkjQ47BsNQJvOaKsprd/
dhNqZLoXnuw0W50BrlEskDDNI/6m2PmE9gcFM6X6oPlatgv06+AVW9l+zCqPtsNW
xIsafJ274DExjiILkXQkaW9aFfhNcsLEtUItTIgK0hPeJRvnH2ogTwrLeoQO4Iv8
WYotQ4A+vrHZfW3e1NchETcpcP3MSoeHB7X1p9fORn5SiDL2NABgznsbYxyOA/V0
vhG8FqyzlFvDDF6B2HWF505CSmxxNuNzEMgD7njtrujeptiX9wkUgnL4ZTqOK3Oe
1nwlEFDKU9Q7og2o5NgdCRjHfFVTYzopAj14Z2HUuT58revZRUpqqZhiiYEWYPle
+rTIao5hTtRuqdg2hzsdUypCEP4q0MkdzcH/X57zMMXZ3aA5aWOkADXmqNKx6LVq
pbToT8nYhLcVhZA09OX9NWurQS2O0V5XFElLfiXr3MgtPXjxXIckW5Q4bvaO/Vl7
pkJaBJxdEJk8F34aEzOUTfj85AwZYIZ2v2irMXDi1il/KkEXdO00ypdCU5WFSi99
0gL70NfMGDj4LQJNSxo/D0+5CboIJjYKYgpnswqbXs/s5Gd1CPk6e62MAKI/LCx5
HOpx0V5padaxneVS2Frkg08uZrRDgi2PFqwLSoG7LVEQQAfYy6mU2U7QNW3IyOT8
qTNU5gHQyLxCmv8EZForPcNQUo2rs/Kp5vqwfxlPVCZJv2IsXH2KLg2oYorTVgc/
6p5g4HGNY8PyOhIJuTYb/3IPiXcWAM9DuOjgDnOIrEkV9+IOTImoT3hlv5RK5M+4
7HJYxxAr+VRYUJh6Uz67Zd4fp9zUg/JB9Zh9xWcfpZyuR05hqB+jlpNuemDys7y+
U2TQ8KesnSn/1/2hFHm0IwotC2AVPDRSKXT4EczxzIjELw85fyHsBebbOU8pFzMw
mD91ufED4rmOvqoS1KxyLNOx9S+jXi2rgPKd0flgyM2p8IUF2rQwGeDIAC/WSXUO
xNB6HdSmB7ZQsxDEwwRfWq1QuazlRB6b5N9lXRVq2hGFBmcxUSGoytz6+Kk3VzDc
0JMBiwly95T9s3jKruHNoAgS+tvt25YEK9k7ZuDc4WZTHmBJlSs3VVEaUBz+TOY0
4JE3AMNrWcyXDfQs9jL/RxglSTwE7yTdhXtpvjpn9kmM6Z1wTQEBrvevsAN/09oN
k/y6LTXJcUTx5SlETNZ/sKXyGHfry9650B0dCHdOPF+99FnsI8WsFLvqEk2p/VU6
zA9euannRUar39AP6hLqbL2IEktRsUMK/mqBrGwR89DrQY0xfBMM6j2WXuw8IKCH
Lpns7PB8rNVtSLaFDoqhR88G3wTqEjB2HLYdDUTsFBV9YsnHs8UG/xj73fe2d2vL
CI70H/yptaOb5th2PMGdJrTIgultmcybNqtrlEO1mDd6lOkIcnwGPIhkJ44I1fPC
1b0GgRVOtA30CGq58tYdCPmNQwnl64ercQD9/4tQKFZFnKN7osLQTb8Mzw1NLsXJ
JvZD0KIcBRbu6OIK0HonTg6RBsel5+3cnKnt5apxJJaI7vku9TL8GvP87sdag7DT
5dWkC5PJ1F7VR1G2U4Ocj7ayUeDlgYN63gOzP9crZfwBjP7fceZgjWlldD+d3Ws6
bFXLikq3uR4ZIqI3TKtbqyeFsy+k1zCTahWPdkgbPdWN68akGgswRhl8uubysNW8
5rx7W0Ci4tsR+DCB992PedBSZgvWFOlrwKGTtPIfo/mlISdOeXDkM9M7ueCVt2Re
rsk3+HrUpBofMnzPUn3iSt1F43+TPa3bQZBYlIb1ZEHtgJgcs8e+ec5is1f3wggf
/0MzfWlpiM5m0eNlqnfj7DFypQu/qWVf0tfUgamtFPjOhj0UoKHfrOEJGus25Yf2
aMy7qzC55kzqj+vKp7oIkvWxE/yvM7HKM5nGtY5PH7W4n33/lL33L/uxdUIFuCuL
oF6wbv80egiBTMeOCcuuzPybweGyvvZfvI2biJsFM03MFTmBUdmYIXnPE6b42MBJ
QKQs38Toy9AlAmHBfKP1UaNEMkGPZlTf9s15VMPIrfxyQ1eMA9ns0wSXoHynfVcV
GDLOj9qM/HFec82/xf3coSLet51BHJeSJMVA6BDWdHIKwyWWb8zN0TVgObRNWGi+
/WSdsa8A2IknUAbgRz/d6HB2Y/hV4HTMMqNpTq0EiQSqxVqulcodtpBha24m0jiV
T9rQTJBwiTFR40XO6QlUX1cM5c8vSFmNQEQkVCUT9FKwUm8HV14Gi75NFr8F6xi1
jDHNS/KQOmAxhhjbRxSOZVNcANKUmhJh2CCihyCkpYlqroH/Vkg6quJI3btvnKYv
5Va87GBPrtCjqwV/a0tEnkFdTl+1tgAHw0a0sSYE8S7QyP1LtD42sWxaTRm1ocKs
d6te///abY6ID4BZJcLYQjUx+cZfIJVL2H1hb/rbZ0r4Am3IrvwlyrbfJYfoSezN
0j6ifWboxMrMky+jKBUukwq1ht1zAXU+2yxSuYdqxsyRqv7Q0dA5m76DCDoFiW0+
DpKWYBSNqbtZbb7JMYyKG/KV8iO0VzhE9GubVvlzRKREv4GA/wFzBeoLqhytaKN/
soewyHvtoF9Nt7ETknvqCNkfnxRy/qpmsQjpE6Wbu8UnnScIJoo33ePro2qJSvh+
Yst5XJn9Yn1JfeqsbsfPJZUv7LDW0PDs4RdqQp7BTa0JrPo1cOMS5pTv/+7vosCr
ryzoiPFWmcnC92TMBxoSCV8hgudCwgoBCzuPKEe8sPXMJy2gy64OJcTTSfaA6eYF
cNBp1PiYl2211zjKVl3bV4IlFNz3b8LxbRkHE6ciYlOkPjDh+zS+f1rfujXD5hco
lKcX36ZxtgO56Cg2+FkyGgVzwRkGLSXGIdYNr1Pi1hJWuTllT7xl+BvRegK8WWQc
RzTAkqCQS7iRrWoUI40alAWndQIAQHIY7Z61WT62i5mb7TTDr2CupTyfqpbLVD8N
9ASYTF3YKQC0P/kG0XMlFJzx/+2t7I+hBND+e3x62T/knzsUxihZ2W4ctCppDBUb
y3Z+/QODLa3gF0zOMua6nlhx+Z26GNJoUYAeSsiKPlj2127GO/CzT+ISIlXpifnK
kqAKzRQ5p/9O+dY7LmouqufZ35QWcmUpdp6hcXSSXflGw+Dc+YVyoISLHX94VqEM
qqmUQ2X8RAgQcbWjhMsjyDKWBa2H1+CMEtRRzbqbBpy0YfwIDILd8dGVmYFRKV0o
j2hruF0ER2DvnGBrEh8GqPC+V5a0QoSdH/4F+stFNrEamYrE+lZf6MHbyUVfZ/i/
EvWT7J6rvnkCgWthlwh3vROs1uzePj0+yUPM25vljWFtwcE1ihtBj0VM+O0lDyYW
iMk6r+aBMFLkRMC4UCqm5+LWZ/CAjOeqaB365IDAUIxX4BXd5oCnuP9dwP1oAVvy
Pd+AQL5IRlm6h1a61+h5ZLA40UaM4vHJRLhtJYAGPfw6kJuePhItw2vxrWFKtatv
/batVnRR5XjYvZqZZUStyNm960B8o0Pc4A7wJTUVsZ1I0ycT+pb9dmEALDw1g1Jf
CankpxhpfcyFNtil3OAGPT1xtdW7RmZBZIODA/jnD6PmxXpUFWgmOp1W2nLmDML1
TQtmttRkjxiijUzJfYgcpRLlYUPH9zceyJvmzRU0KX2Ue6x4l909QJ7qnhBUJ6iq
sZDQg4XjjfICqam/QUb9MThmjflnybX5ni23JrQy8cmINstClvmdQ10UzFYjKwKa
b1kI7dAC5m9F3utegJnUAsjS5CD9RnuKfvx+4T7XZ/iSKJft4LDAdoLIw26u/I08
yz5JxdYjsSabazwIAChxTI9rRBhnkz6xxZWq7hKyLOw8gG8AGkFhwyKaurMtq8iN
7ktKY20Aq2nDR7NJVZ/HP3IhC86mkTZcdnxdAtdeC6NIYbZ7pV05y1tl6jJ1wVcm
/0yUYgIHHx/dEiLVCJ08T9E8UM+3l/Lb/bcWowgOw0jCCGnnWNwD6ShwZBpp1v7E
03a/synq+MltWGnK7yevfu9moX/ETwBzJBjY8a8YjR5tSsJmcYgHRRgrf4RfL4Ie
qFKY1g/bUZ7lYmsITmrLKQ51uBjgwEMO1ee6PfGs9RFGA1oYPWLNFkkVPjKBYgoI
ZduWnRD6Zo7ghxCVXg8yXEuOHJ+PBJx5ejbCwNUUA9qKiwQoRWOBjOd8aKTWlNvy
oJg4CCUzG6t/cZlLhbC7upOEMDWolNqSHim3WknKo1jxHPQtrCAw87+THa2d/Zy1
i0NN7pD3jCULoyV5x2Pvi+A0afpYSxh7ULjvaCgYe2Csi7+e1VNxIMtObgIijR09
8J0rm4uDnWNBy33ZSsFm0yNlymmcQxirgScRVl69WF+QXc3XeIpjvZP2wzeFQD4h
gxqsa+x7Q5UDji0+DVFp1rQdRR9fklApMIQZMvAx1oF/DAWwc8/nmKKeeRGFWwtA
80jaQOWpIDDr4QnCp/Y7XCV7Cs6Y4AQ6v1TF+1XKFQWXamtgPfHKcscHzJEZkTIF
v+pSwwqryuoL1KzG/JOheidxB9ZZYDuBgQu5KmAixDM7w7mWxZWIXzL5Mi4JE6zn
M21DQIRCr1iAQKYWik6q4Xq0kj1dtCHrn+6g+oUi5MFOL7k1M6HBmtSfYuSop1Dx
o1V6mcMf2xuYkywhZouysgt+lKNtdoWra9PlYiTBlRwKNYbr9xN3+vbq8MJJ8mzS
diuUkx4TLVUb76HVJcut93i8MdEY9A8108yLEBqGcq9FYlqFJd70eCtduZ0Wxcyi
O1xTkvIwz1uDj56NxdhV8UpOaoRRz3nogo8Zt9txWhK4Z02fXWRrIkXrQ4mDjIoE
pzCYeE/DEoD/ytKXJhPapsIYAi29QAl5FXXG/OlpFhKTBnsR/mZe1UIoyHPwLrtv
lH6zAT1tUdelIw7QYTIinsw+gQhOjLyTgqN1OuwCDlu3OaILWrp/bIu/xvmMKQrV
KV9KfNayoqSIkoNcSsVtWR9+Q4QDtI8KQgcvQmXknjzhpP6pTzzFstg3hHHPZOGn
xbNFIkk5eIef0juHjwMT/mIQ3ZnG0YFkF6DDt9ZIQ03EDqMYT1MaxqUF9VJRFKDB
cAXfbAJdkA6sXB+oXgsDCMuhxmz0vN9foRAv+ms7hOpu76Y2Gc6h8AmGLG1ldY89
zPH9w8Cn+m47sPcHZfkOj5Zou8uJCsdGUFy9pGxjQf06L0bCDxLTtee5Qiav1vyF
a1z4EVPwvpR6Bv5nR/QSa3dN9J7t17hOmxZYsO/1T0bcPdO91ec7h95P58jlBsLa
dbqkpLKE/JuhekdJKhuaZmUwxkfKGwWQk/1Tazp5zrD9mgmmwo28x94x9Ubrd83e
oNpvebGo68tXwZSJkUn+ri+i1oMU49nTkXjwYPkKwrYqGYS+N6M44hu0xsqdnSv1
LGXpRgjCVmUhIznrJs0n8opWswbtYkRXjdEkYl4UJ6CJ6vBrmCkz9z6aDfVN26kl
r2FdirPa+oHQNWDoz7IoedysrRwUrcyal3v3zUi7eGpSHHLb2q2Ki1AbcOUHI/AF
IFnzLTtJMJtJVqfkw9Shpsyw8bHygG2Wyn03DW3XFHBVmnk5MhFb4wU7UQfpNpvz
CX9g5LaE5i6FLm/9wAieQzcAKw59tCOfCWIEQCvksyJf5uM213z8gfOafRcMMIrL
UP8bJ1DY0SOVmKfQ5PbuXYE57wbuVX0xsABhij/LgzHVaAE18PGTer2Rkkj1itjs
fhd7HlUuFQ6cqPm9TJAL21WgCH45BS3BzCJRmVEJAJl30baIpbO9GDER6Y3e7zRw
7a47QuzquHN3UUDdsrqo1XtimCGDY+lMZ76VstU4o47wOPSab+MmU3JhbAt0Wd7w
B3IEU5C50fzH5ipxxricv2tC6G49gduT0noxDu/+42MoinjpbArxR2pkVat0meVG
rkua5A2clv2emT5DqfOqoVZgyr3YoSgff26veKmtZgh4SKwUTB2RLpdG3FKvwhi3
ROx/VxohtI/ynIxqLFD9+UQsIvsLgrOeYcQ/UshWuaKpi90bOiJvTD88StlDPejw
rk1LnVsNyTYrxkLgUIuzamdmKR8zWUZ9Eu4Rj7jdE2o3JvyobFYYyTWknlDX07Nw
Hnc+Y8pA5R6MS2ja/lFV4Q+ILdzkr5LilrevfJoqZ7GsBMT9xSQe8oFD+FKxXwXr
DZ/3TgvIqaP2y5zLQYoxOloiEVFxf6qU05CYaHePItRlVrl1GPDGzM5gVjGNWFB2
+2a8PsO2bqnm/g8nBqf2TTrQPVk32LGe6U0Tu5SqURmdb+RwrfEywPB6DCia0EMq
UBgV30KNv4OKgyOI4A+e7lS0LPzcE45L4TNkwxsLm/Av3629nk6OneHTqhVnkzFA
dpSKz6HaCtdUeMOVND+/Ok4P/JVVcEQrY5g5jJdjC8t9O9HO29FC1qIh7VWg/42W
tx1NTr+K3qCCRvVdevZS5dYVI1fH0IXKiK6TCcYXsg/b98P+CmGkluiX4Yn36+8p
VGo2m9E4VUb+VsiA34D3c0ssSAkQKA/vSzhRKYnCnZz/kdz/SOkD1RS5QHGZa1+W
cn9XC4Okd6CJz9aT03KQYhOxyDmdqr6Dyh04ZfK82eK/sxYbpveqqZ+rPWtgLm0W
EAMqTygfJ9wtEOGbkJkA/EPnuS0U+Z81G49p6xN7rxxi37fYgN1IGK1P6aCJdy8r
SZm8Q74gko6FsWGKs6wpiZ5Jl4cHKt8VPuvTG/WKJuVcHIA6f2hYJ0RiD2aSQsRq
zF9P6KHnkQXVD2IXcmVmYOgIMteBok9U5haNKNaGMBjk29JoV9rKzTgW2y5cgRpG
F2B+V20BSlclLyjVl05YLsJmAhlymdus1SpyuZIKEdBDk/qEzGOB/QqIrQXAOsqo
AjQS1i8AmdPFDu8F7HyPztYS7I78ExYV0eQou9PtJkyRdzJ/GEaGdV4ORB9mWBDW
/42IBc2L6d8YAyzypMmOHPxSRs1yWtDhkpwfQHSoRW+cQom4g6N5bUQDCZdMqDZ4
ifkuY4jfO0QqFUplKcBCFiFQzZngamDM/eeXp/qs4TodRUs/SMoTlo97Y7xP7H20
MLi3SIz8kZortZGRnlNHx8+PEVwwZL6JlZwjR2AhrDrjRg8KSIpxN9kVoXvIuBlF
i7TuH++4YCx5fd0DIfOcCUQGv0bgo6pwFaUi1NcwJhUBMHBZEyMKutTCTEineeMm
5xaol8FJ9yi3KHJSJjMEkZUUB4wdfTEP/ovyX7Ha5eRAVxYdZ2zzbymGxkHy5gRi
Sv3r2EP4HxUAz/LaE59KEAZMVOy+oae+bFKAqmtrXrBVBQgaxDL3Q3UsVEg8yK4j
mxaU2TFukm+qbAk4gxyuBS9Gc9gx+BC0a6JdGtDsKHIdbgjb/vmnunMNVGjc4weC
5NMaOXNe/1AtgvocVQKkSiceapEpqgPEQHSexZODhNAq2g9KAOJAg/77QGIg4kKU
UKtbdJfr6MLwJXo+YsMkFm0gYlQuxLDLAVQ3xuxX1z8tHqRyr0LqUnToHN9Nfxp+
fM+TkhQO24hprP6dV4fXcHNrJBgEgNHUcdyLYyaulNFHz1ksVcTa6VriYfVLmtyw
zQXjEi+XFT3YZAiYo8r3uatLM6/Z18OdQ79gqcaFm9o0BTRTV6WfjTI2mc9JOrQr
knugSbUSNzTPktKY9v+eHeQkVwUQNunI3wVggJDikzlV5f9hb7WVSFLuG8Ong+um
rT399DWNW+3AXmyfrNzVV74cEjnrqflTb1JBT8x+/XPb+sRL6VfH/jedWqY4uY7B
fjXcOotOsc4mcExq7hrYYy9IEb/sdtF8lJey9ipz/QWWgKV+3nKV4kz9Sbusii+I
US0EaK4wx5iQMwjgrP2PqUXuGYVZ5LfD3v+0H/Mb055nWf7ZKzw3boHN1oC9M+hl
hD887o8/MWWqAuCV7t8m6XIjnRA01Bmpo4sgHlL3D4x//mRB7vFEY0tEYE3ypfBx
RvhiwVR2vajteaZqot9iTAk5YaHs6gwLs1vRLOj4x8vq7oBN79/Mx/eY3OiMETyS
ImAn7iJx/QBoRedFfZpNlnLyZPRArIU0W6ibFTtb4Ibulv7F2T6H51Nct70fxvGZ
TP1ZGNoQY074PTKW3cCGY4s+O4RO6jFQRzs6xuZ5Mb1K5FVXqARY7Nf1JY3fXv3n
DEKUrSpCn7sMGI/ZPJufMktWB5ELH2ygo7/RhYxjHXiHhVfAsGe1WPP98Z1l0sA2
xlSkDFZ1+teJa/qyFkkPQkYpqanVolrmkWcuR/+EGd3ftmcVuX7HGg/VYboxVybc
4LfpnKKFpD8d3Z7l8s40FGOdBxb5/gAqC2P8F0Y9w+VjEXU1fS/I4oUri1C8Cq0K
c3sVB8wwkhrhiXl08quxpKIoZx2VyiK03MafIFFlw1NTR/wTaBtpX8892+T8Y8fL
B+cwSUm1Mg/QGCmd0ICV/oVdcvEAnN7KeUgXydNPAxcVxsHuD2xf7tGQ3mVFjet6
dCKYW3M8iBL2kV18fZMACt4brULmJhmXOPM/hgLb3oVWGNBje8M8crVlKveo+szZ
lxGxK+H4eUvtPDyp1zPCnRYVLzP9Ta8hrHzrNkAHtnw6mHaFuXfqJSsGbdD579EO
xtKMtCYidEPC1R2xMh6HmxeMd16xELf9pOfRipogvO20blqwPwXzNn+mviUhQu2R
eF+kn56NErU0KZ4xjSeiwfp9vd11uU8mQjwm0EcJ238xBpnZ4YpvQBZHCmPkIa8N
EWIuM3vJMjHOOBjnd0/moeHL3Lz48P6HW6e/RWg9hfA3ZhBUN0V3KdPIwfKo5NJH
JZSaVvwQIQEOh7u+ZR5cu7Bf1U/p4jlcZpCCRYWAWxDSxTx4B3xeukXTcYbQleb6
L+J2nGiG/WERrTSV1HymDUE868+27A+VnNqAjknCJGHyxtPaTF8sXGuNxoosJw7R
wdezEIF4h9lBurdhKEtNyd6YZxO7Kzs48dmnY5gngloGVnOUoeCsVSOzlVziWc34
rp4AuzEbs91TwjwOMWgH9qOPrxgAYn37ZeY/wy2E2gpr90IMmOfhQC3SRhY70nw1
QFO14q3646/oXH9josAo0ym/Ed3aDApqiSOJAeZvFYUqT19fN7Z/fFueh0+G7/Ed
u35j7bkGystGPF8oBdJI1JrVN8OoN0EI/UgsH7gnstylaQAeVLhlpy/6zlkTL6Gg
eyt9HoJIhncaUhCBovO3fp7oTzi58Eb5We3ZBaNOUN3XG0ENKiag6/aZz/txUewm
2xOLKCOCbFdIsnbi/h7nBAZ2x5LseghpRS9ZH4QYd7ge/Tm2B1sH/vvk1CYa0i6c
qtBFgnScrE7Cjq76japQsMgw1Ov2vFAiGGIduUFEw6VCqyzPN1xRVKstQt8M4AXs
3v/jDSICw2H7/7YhrjxC0YjgDUmdD8Dz+eb6wqdNO0VauSlYzr4//2RHLqd5VS13
exxjWqAeh20qOKHVbJ5IHZFFm5qpk8syPo64KhzD4ApBVMlCy4MClNyGu1rzOa8r
cs7qwkwMI4kI0icElrGp8vzgt02eVcF/Am09U4ZtVOMZ7DehE5ufNcTkmXcXwJd3
uRFgF6YjzPniYALYpmZaDWtrlgp9tLDldKWbXxWRSvo2z3aYKfJG1Ha5Ogq7D4RH
HmaD05m8XYSAHORFTJoZbMAqkxo0niGi03EhIKq4KnbZxqYsxmIWvJ4GaMrwYdXF
JMgKG2aiSVbFvj5TjIglndwbcIP/cQ4FjHGKIgcoeDuLBfW8gpp+Z3AnRAjgD+fR
PIK31QasuSfDKQwBacyK7aaHHD+Gaw6ZABInAR26Ja1nFTn5BqJHNJW71ZZ6Lu79
hHQtlzCyylZwZ6+BKaS3aM6mDjEuYCwOJnopVCiao6zOAr5B54eJRbLxroE4zXDu
MIc01/naO8RsaQaOg9IdKdptXMAijArunkfcCXoTtz+9GHy1AkB7IbFzCaOASr1Q
nXQNMBiL3Xoa3n/hQDq1jCnziNfTVm2DkGWwVf76JsqHYJyaFub/0XScjFB+k1/4
cz2ISrQX/+7QsId7MdWlVjX2tlyl2ODEdUR4oMLlwEqzXSV7+kkWDpdHh6h7Usq8
bs0CKoxrR3jJLMzUCkUtYOCo5700ZKghcYgmd8JHTgpYbqDYgnIZniUPQRxemeCl
/rkBX+qSfF/eIL/96OBlepR9qqNedQQQwqPl10t9VPz2TsU2+t5xKwh5fg79tOE7
yFQFaeHb8zkmwuk7zhV2iSuDwyZOR3xylMOgnU1kxMkKzJ64nyfawgQ9uYiJSLw/
aCtW+PmEj5z4evxg3SCw9QwBA10swN9+xzT9dRC4u+CXVqDqJQ0PYpU7M8OfkbwH
Y3NLNfozl+WzWYeASMp0MDqS3Tn/NEfv902uKt0TaBUU6TVKC35a1fHHKvP0pf4U
G/Cm3g2QIUrcNrYBhEZyUc6eaYy3o/brA59KwioEJLbDkO1vCyEge5hz8oe/b/HT
bbr1AlITaj6WwyKsMDlXLOS3b8upTMtB2HEj+n1GXydsL3cRUhfiYW2ok/IJG4og
O+gQz94+UEchMFHNUBl0xk2lxm+/JHivDkOylW/A1ux0lHNO6BMSOMU2Fl0SvH1A
5dwi2f2lLuLTzRRIKa5rEHZJNnSvfePWrUIWinRSJ0Rl/SGeX4xb/DIIWkl0e9vt
qfO/daaU3iBFnAKsJsTc0XJYmx5LdvXPVCwUybriG7LhwehmFNJzD2SBqLkcs7/b
sjvXVuoRQklT8qSgC53ZyDKTw4JtVy2afU+qXLn8t61ffFM0OrXpGV+qH1R0G5jI
57Qg9rqwEMPW98ORW4+XCHRZQZWPyXrIv4booJgl8mH+bo0cxNrU27dvX5rvN0by
xXzte+rj/GBX+UI9Ck6Ifk+ZNOVlO9alg/2KayAeJoMy5+XwJWF6ActrqENj1mPR
E6vl2MMPaK+TKBMTCn0P2z2wLkjebsd1QrFdfKGVCDl/vjbd9cRPVjF/Ppbm4ob5
V2pfqkaNc0PzEMPoFNLEhKScWiDrkgcUfue1EHeyKfdSpTsugzB5rzwmAHaf1ZJt
2ViB2tdcNftDGeCrPgDIxQZ3Fl8XyW4bCTLul1CNcuxBL9ovNam8IYuvthdngUIt
ap+cp0aTadBQVXxLM5eG5dbMhJFFZzdTRtX4cBRweCNPPLwkgKW2YP0Kghv8nXUk
Rha7e7WfTGXJC3nNRHqsGyzKfsT1LUDSs+tQWKESg/+yLUEDG5E2v/EFiVRzgFPL
VaTRpjTiz4cA9XbP27Q7AKwJQHWnSqxS6kHDhnGYolU4F+kf2xsFW07Hz9rHZduW
+y0rxaKhVe/GuSPU9xEUzoLDJXyBoOp2RpQqhuBZh6g+uaCJVLP+ir6hr9dNAKC6
hWDzj7soWLR77VAwpfPRntEZwHRucZs0ejemLir/o30BHQvulvXreXluRysOCDKJ
2DSi2Z2kTzJY4XQqpC3Mek+56ewvl2ug65LmEm+opz7aA6459NOr3ETgguEJFmDt
+fGlT+IrT5k8+wQ3mtVxl1gaIn6X9dePfIe5CcHSIlBlaYcl7nqWeMctUoBDb4hP
HoDkmt18g03x0a6JSdoMR7eaUIdz88W74Zt5B+yuLrdJD8P2dn6Q1Zqigup5lD9T
hU7BTurZkzN9Edx37ccqDST1jHERMR4l92h2VFebie/5r1rGDg6L/mlDVFThxx7h
LkjQZlAab9KPMMhQt/hWz2WHVDUOHYfir50Gsnsl6fBOV5TrZdWaMxvphnlSvY0Y
yh3IlV7Jv/kdxXASCeywhSVDP8zNIMtNNWY0EaeFi1l2uRf3ut+7uwZXVxmdibwk
cPcklzZHgjXFv5WijxkkdLCm5tspQGK+6GvxGilACK0dfB6pVPlSU1cpdkwvRPG0
ZhIRq17dqwpWBC5foAWcRJ1/MOENElKyX9JsZz2ATlf6MfIwJ3s/pqG5ANTcA/8h
B6BGEdSz8cxa77WArj8N0EQfP9FaX1BG+6pXEeRjmm1/KSNtVCEOynmmszHvqUrz
EAkcwHuye7ht6mb101k1HDsyan/KhVOZcingqR+AEv9lHsu+LaCm3kqRjeGN7FV8
DlVd6WTCRQ9sQEcj0TmROvsJtF56BekLbp/XODV5VDJvnQC/ZUOpfRytO3MkE5nv
Y9h4JwSZCBiG9vTrKvLEDR7BuroVHBb0MK9OgoaGaQNCJNc9OfeRFbTI9tYHJ8ed
klFWGBTx8Hbol9TfJcEMS7qcaldoMSIbmafwuCTBCGBAZ/3CkbSjdA8PfLSVqK2s
rxox0hoxiYgc++VUgFow4VRDikH5Lq/LbgLa71pyJE+sJXWt8FeU9zLTj63Saqk/
Gryz/6aUXEPtG5ldooE4w7k+W67lZHO8RLulwXkrcdDxRk6wkiZIfWMvGhe094Vi
s2K6mfUmaJ13IChSnSLwMFWaQo76giANteaddlFB1uVW7/Fqyt2N0wLvvhmK31n7
wTo8+iETbxYb82+iCBJgE3/oamSFyHHrOboP3ydeBHlK50efYh//gMzo7mKS0tx5
Q7QCG9w+K7xHQlWPqhytnl1BXWwOnv8G7vhfzHAKXEQmzA8o9/L9dIDiPznuotWQ
sKn/0HeZLuxhc+ByLr31ylwPlJEQ2vXzj/odyQ/ZXcuJ8waCKbr9kfqQMspIxqDi
mXkA+E974BLc4jYSsdTb/OElRyY3zUhnVqcc5MHr6B83cGzlsfNs3GnaHaJnQaRO
kNaJ+2+AHibIb+FjJyGAKAqrzxXW6npKNVl16Iiwo6JQFZsb9rAwQTZY7R5HT+Oq
fGr+ZqEAFpIgjeKfK8FqnPbsy/ZCQAMqJItYn7C8jBzEZjyEyPcVtFKgBbps8ZAg
dsv2p7x7jq7f4T8U09FbM5E7rHW+W8h1Hw86/wy7lUmveHAoFjAG3r341WSKfqO5
ixFaWvy75N5/uZ/FrvCJ20zX2/HlcCeArBkbkQ3flX0TxTJzXNi3PgCfQDsHaYNa
q+TwcWxFk2VUY27ftYaALBQTHZgidh0BA7hmFuhJkzB0d3clfiYtllcgjhZQR9eK
iJ+qegIGrIrFeQ5D8PFV59n98XV5AJwsPpg4oPiASrMbnZnMICH4LPl4amYsGn7r
lOwXPZLDcJO+zd7mO5VxnnVjOVF0OO4VC5/yU0cgh/YzWMaJ2OY5GU9wJDR48BAf
/fpbLGGecIx8BlmyFamYMbbNOWt/stmWxFZoITHclgStX8eByRwMB9ir/9ULIWg+
YF3KJUictpTjYJ4g77zoHEtfPK5ItRbQ3x/Gwz92sGF0a4Ihh9yjMpsDVFEoJ0H5
ZzTWF7k0lOpNtW1S5zw0YANL1PUBMhdZWuepRrFq2JsDiWlyc+nTnQTrLxP02Sw0
2a60R0U0+z+TAsUGNX4YWdFG9HFi6bOPSq89b67NPFxRV0buWatm6mPGWWHIQ5+a
vFbR6Pimw6rd8P0Vk8yVWJKycULwX5j6bNYNPI1eR2ncjFPaTvEPRSX4I0rsbaV1
W/FXXTMbhacmAkiv5efeC3HgFcVN3mOCnBQbOT+byiuEwvnveqBWUTKZBK4I/gup
qJ/hWKQPrcIcOpbUmjoji+hnSTO04KaXwor7qyg6A18zRrVw00rpwxyitQUsblw5
3+JZlKofgEAMzg6he7p6TEsfOgJPMtAs9yck2fDLPjC2f0Cr/CJbVhegmLny9XaE
xZmjC+Qa7o/CRRcjyxAZpbG9OUNx6R+rEHKO9B8C2zdYO2tBKjPYNfHUZhZmQ6YR
SEJSCf0+Rprqc0LxQDFJUm1RUILc/wCmoHa+VxaGgzRtGnUvRimLo6k6bZD8qWQT
/g2aravuSoDeRVJtnDkOtlMxfYTQO9J4CnkgydLZgeuubQdcmkFKSh5yZbsK9+5C
DfaVdU+eRHNX/gMr8cbZhCeeDcGAUd0qWaoiwypxIJUJ2HtHdlWXm1N2HCYXf/my
ZGkG5nf6gxRkSXJvGLLQyFJ51gj7LMvQiXB7JBTBXDuvHyG8MSzHWeZ+RmJwhv1f
cEUyWxasIr38drZXccdY1Me7J7w9z7TSSE+wfsvLYCY4jjZHOw5uLZIFKRXJTOr8
MFkwXC3JYFngVCqgbUiCxKlFvXXnMxIMNWTzu/Bnsw2nfXyfdGmU75ie+wGce45P
wk6aXLQ7X1LOyUmdQraowJg5SdXyYEmLaZElTOcVzsWWobi2y32J1fo9RgBPAZiL
XyYE00mJzZlOJeoqrK2mnrv4Rv9WDydme75qUSj3atpqSfbcExotD5ATfVy4Uchi
lqugJ4COFSgmDeDoG2Pf8udYXUDQjOZPQEPYukB1f5KgmE6s8q+LON09xdOALF9T
tc5hlkPvWOmTLl8ygdNfZ02Gb3Xb5D4ifeUV8CMlphpan29msg6j1Rn9Dof41z3y
h3saUViJ/JCN4DAM3eXL/EQzvfZGFujzzIuqTkux9Arlt+cjrFQcBtJVL55iCtrU
GKaBXXrjYgkmJjOE8PASnTIbw46lj6ntK5fIuaZrCGwy1SWkC0b6BgpFP74PA8KS
HxR4RynzVq/FYSrb+OJy6T6ozIqgI6gcxqKxkqmE11s+/mMqRRd54FcfBZUoA32O
i7B561sauNo6nNbYXsVcnkIAHBwHlCQqS+0wDsWLnfA8iRs2/4z7OWBNeCN3t/JH
JNHL0LgNdKxWcYU2YtnOLDI0Yzkj+itR7twF+8SZ/paOwxAoa4O1Mq2BCpoBFAhi
PxtgWNLTvHShDcFANVPzJ0D7n40RyZS7tfdxeMS8XJyFcVDokNp5dWI/IUJWtepn
lWLBg8MuU7HTMLNbe8ZkAAqyTT04S9Fw/DVWei31BGtmbiEqnxoeLMAYUYg+btmJ
3SG3WnY/ToY7lVWYFERX2/pZ9VD/OTNs9+MsJbXV9PxZ4QZtyie4nUztQp+q5kmm
6fH3SIOn8nrwapVx7aryJi4QjWFa9UD3FzDztyoMLCC73Pfo/ZnGiPswbmmQlfBg
mYgc/F63uyFpAAmcs6lbFR5I1fyaA4jUhG3B6GVKfbmcSmb+l2eEySwnJmx2Oeu3
3QnGRizH8SOaMab7IqHJI/CEve/lBess80edWzSwWjAOguRNXOE0q+CdwIID8Dv1
kY10XQdHQ7SS5NJXRA9TAVSXQnrEsx/VNLVslz4WnRAj+z0pEIgaWeb1vKi/5Zjj
nDrjTpL4Q0rvgm60CivAVoslg8Qert6/Us8Iuc5fvk5jcltGUsXDw4z1M68K5QJh
3jNCG77q7fdTbsHqiCqt4lMG9PudtqiG9etfWx7IaQfPccbzIum6dEAbDqRv1RL6
jLxnXr2ya7nLcX6PDImMBfmPlPjRj5msnEnesM5iROSZuvzj0jT8ONWt2dJ9Vw/u
vWq/8JEgUgyuZHMlesRuLGnKtp//waYE6mtxFosui9O9Q0krtkMZFgMW7qkYo+zC
mAdzk7E4YT+can7J5h8xma9uK9EKjYg04PpzF9xK1KCwGHohY4noEJ5EVgTDngEW
IRAqouzgnuD2ppX+w+nyTf07RGdP0o7UHNNJOMNRA1QLRqZBmuBEWmj9OK1Hw4M3
zCs6hP+jD00//BSke0ObpniSwJQnHJP3QPkginW25CLzZ5mQw+DjW4CF24tfmMxO
wXakYOp9gYWaNKWU79iYwOzdFDuagOZ+noYqvCtskEkBZfQtL3qRApwHJrHYDjB7
d9Eu3mG5QhZB6/8RM9w8qXY0TBwbIjBNCymOaNc3saqweaYhnfFACK4CIIULcFKu
COMCafNLUjuibroFMjt9rRrt16LhGGSHT6QmjzzBrr7icKRRfw+ZbS4pBhsPLBTg
G7CS0BTfll7lFjo4eMBhdysNVfuyznsy8PmYqPcM1mBSuFRI59WSbFckVUhP6Hcw
E5QaDjxmmQSd6yH3LnStzbtgWNfuQ9Rhtuo+0xoGKb0v+8i7b0rAMAQ5CCREjYit
NiKl9b7+YsRBpPjtgqUSmQ+9TAUYFedy2lUp82CsEUu9ppRDqoa1PkDKEfbioHmA
JJcUPAOXmspeeOEipt+GPGo289rMgfa27x6vStsUVZeyqku1jrjc3NYtTkd7tXfi
LU0L0MnIODOA9BY9VdrNZ8Gq5B70lJxyAudCxy9NzABrLY/ccGGy0PvNyGBwAf1C
c/A7lWTpG5HNI7RPC4+DWr+6aErIDMTHjAUMKRcY1FCg+cggvpVg57Wk9lr20aMa
U/w2Xr1Bizuc5kjJgt4fl6dRogV5XTCXfS4xO3I7i8QLo4jW+/kuFZ1jZEex0vUp
LAklRu/eB3wpeM3jWSLZojc7a6M8CQkgoQxEdeUvFnS3n9PrOpMBvXtvKTaoTqMf
HJFmXZmcGETVViFA65WFwGjp6aczL4AY7EjQkNAYohQC2yfoD3pEv2dhKZJDGLPZ
GpCgHjK6Ju4xunb/LKIU3rbtKBYFlhCTuLNLnCBohCEzVxb0bag2jkuOrxdqSYC/
UJmnAXC0i4Jc6T+XdoAUCsAsR0dmYLgBBZWMXOPz5i4Gfu3ZFqiZGImGBZR47aJp
jcG6hPMTHmz9iOE5IlCb82EKzTwyVEThhfhm8SjSluU33Jr7bKNvVrO1p60sAiA9
dAT96Fw0Drox+O/1xuNH1W9Ob8k8DW6dbt+hAjwMro50k2wnM+2RNBPIH6eJLTUH
e0z2egKiPW94V7uN9/tBPlVLPYktM0uKQNGmP4xBC/nR5KpBzQel+h1cp39hKDMY
reKIn1WTsdQ5ztmerPD7ngueNYGZ6/IP/jrIh09/VKt9UF6MQfRdWEsG3IettQ1u
Th3lHX2z24Jqb91OlIW/dJeBT2a4twa6+AKLsc80VepWZc+WgTDObeMXrgUjynyx
wq6MN+h5q8bxddAbQdq9FYfkGbaHWeQfbETPLBUJjfjq3vI23pjdzJa6iRjHhrH1
zoOCBTMgl2GGx7yl14HLEqoh4ZZCJLPegFkTWlWTYc1ZxbVmtDmJRmHGwvaRwLFX
Yuj0FknsbawmAabyh3fgYAD8sCB97wfFc/bubsaXAMKa3eTHbjQnfj1BVUrH8Qp2
1DNvCvwhWUiSOatUjnL8hXRGVwVtT20SyZJZ8N90Sfif4weZBmFoYCRwl2DH4fjQ
OHyFX4kldAcURraj1M9z3oUt1wy1ldTEHElG1mU5n0UjzAqe2q4ztl/+X2QfhDTQ
GxoEn5Yg2o/PZFJo+mUIcpSl09y7Smsdd+wg8JaREqfB/uKHCqVYbURdx6xsHUlL
2LXEWGmI2hV/sJp0n9HidKZMlzU/Ad8qzAQiz54cYNbNP3NcwK++VKPrEpbaoATC
EZ8pvsgToOFbWv8d/tRxeAUCxH+Hyd7nK5VvhgAP2I2/KAPu48Z/nnbpezJ6iEBK
QhsdKCUy2POc6EUadtWo9cWEfT2dxXvZAhnzlPL0ETO+VxGpueMKdDmvCC81LHdn
9UXOmUTyokX21rm695W91+P7Mh2cnDS/LuuUn3d1t6osCVs2ATNNEgVECAyJcXrE
gufFNYtD1jAcjZrJTEN2PJJ0ESPC534GtQbcPdO9t5x0C0DabqiKRu9LwphoXC6L
ufFsGDclgxu0VyS5yMrP0iolyK5RCoQ8InPZ3xuWClDOzhPoqFaPIxP/Fz53mbHF
mXwIwHORurT7s4PB9LTayGvH9eJGsHM00BuaQuQidtOb0+kVV3bqiiNrF7ND7Dr4
ZuwJN2OKfsI5CZkg/XkVQfYAAKfuNOEA6KcbIB6HC5T9whCvIu7xdPprXOHsdu5z
0b68c6HQHICBCyvChVQebctt466DV8faRl0WqZbKri+0+bLihNrHiUxTEtdoFk1S
P4f3GlBMS9WEixLljJf1bSqy+oMgJDS2px6ZOmXvLhD9HBhM2SrSCQ5w6b9mM+jM
c3lq3VkZAYP7m6bOPdVfA9BQtwLahCjO8i9k8d/YTHI2DKRzBCT4GVQMwB1DtSN/
umw7luJY8ljMqdzqEmb/qTwe2L+mEQRqjUwGzqNAkOXB58MfNO0NMIR+WB0WOxJy
9P6qopu+j7NM/nA/x0Wn839zM+WHJABTda86+voElBQqPgRDzA76lcnR5IF7hfua
xcF5P7fjGTcD3t6IXngKJ2BY9P8cvUU62R9cIREuA7B86CO14ZdE7o1fF5/ExgtI
qy4dAmc+ozEAuwB0DjQ8U20pf0cIZlFgJ3u5s0EipFrwyYgGnELjr2xP5ARDj6aG
JIC/H2o8LVemNMV0gSCpWC9gTOPLyJQOBIDjjsVkh3mxggpPtC8tttRSj3dE8pLe
GWPqdBx6RBMcTBpPUKyKBmE7urlqVx/pnc3TIrtH1qPT65oMCY2sWVN4We/srB+B
ic9XLapZ7NRC5L3sCxfU85HxoC/l7ijNaZfVVnVDj//+zm1b0zmGEm1/+cr6QNW4
teGUsYNVM8D2CYDaEgzqGbmLi5kKEoZyaM5Jkk3p1UrLPa/LbjQ5neJDAIU8OiHd
8BsjYoNKlfO8UMEZG9OQX/CU0J/oRn+urX+prSILx8wMVHPCDuYUN5CUgcFhniX7
EVrFBAhc76Htc2+8WlDmxSxncW6ct1C59m/atdbrAIahfJJ2TzXvsXiWorcCv4z0
uyzAGNgFH2hqig07t/pWIgR4i4G+Mm+L6ORv8vI9/0NdZAn7fOyQgCWJHv2qmj+i
J8JWkX0VNMWyRTmrfyoWu3MhD52HEoKYWT1J3GePtI/8xvgURgnMk+eG6sSSltik
A3CnEAVAO8SdtRZX5pRuxjfQ+29XMVl/lbcEeCeV5bVmwewzNMstfQX/8PbR5kU6
6C2U3UADvRrTQWA6PtDMSWlSWi3ZYqhR15GFxRTBZ7tkGedY7zwf0SPBOm1SSExA
ot9GxOWsjUKzWLzAwRWywVh2iEXUbfco/sLAELYtvIo5NxNjZdOoTt4yctAxatvo
3nFVVD/+KqDPgpfGOeouR1kfP3ZUyiQz+D7ucjPtxKSGJIheLMRTsBNyLYOmBEKG
9QIHFvserOhSXIZBxN0RL/TM56Z7LqMFLDBKs6m1WzMSIOmNqRzdoaHOnJnFd1ec
zemzFLz8ckN/jpcTKHNgz+KKItiSMQtIyxnvHrXNifXKhPxjRQ6J06bREHrI41Qj
iD3Icuf64lQpuqXBDn+RP3hSqzsIRAx3/ugKchVJCPMyXGqLAxyRSvnfbQDOhKnI
w77dHF0JjCfWeLSFYdsXBsvdSc0WjFGwqGyQpPe9fuH9n25zswaHEGLW5dEMq2zE
4dvr6QsNSuSOZ4vhIc8lU3lL0+rVb7L+NunKvUel2O8qY2IOM2m0f9nSPowa3T2M
AxcWpj0Slbs3uxPc48jrS9PWZT1r2L2WO2rFoN4FV1WDqGF2TEKwFzxgYW6BAnVB
mcYcBGlViaVEKaKLDpJAYtA98gEcnLGK4YnqEs3Xfh7uomd6qGmAWWdPJRa51h5A
35w/B3t+MEQp6XVpvgTmox2hvKyX1fTcZTB37nLTxZ6aBJzYmU3Wu7GviNOzYqqw
bFFc43ndC0EWsDjkdqKrpD8W8oEhR43w66ZNanZulq8T3N/F6cyMfKzTsyGkBhrV
LI+zX7KgW7MOgqkzLpyksNklbI8ZRYMWfZU/+ghLQOac7ee5dRmalL6F4dFuDx/5
mKVXRyBK9RTrrsk6QObmfMTEEUPVRwSM8F+IRzQLPCRK/SlLIYpSjlSkFYqqUpHt
V03RQVIkqV/kIxEAl/Kw6xDnFPrpse+0xN2lP+1qgP6J+6sCH+J+Utfud2B3c/c1
RbqeUurEWjEMxW06sTtKc2L8NPRqzNibJl1TR6ootB/hXwnZ7M/ERd1Jkb9Fd0mR
Tgus2jgiTnk+9Wx3gdy1JxygNcp+UzVFUxbO5/MDUK2WDTfNGw8RTK90KfWBEZVx
qL9Gzq3Se2/WcycTTce7wZr3ZXvjqFoMdbIjLPWjizstybfJPdXi2sDXbCXyHr/b
pW42jzRmMuD8SpmWhgUo7ZkvWfpQztINEgh6szLUAvsiWBmkmaw17Yq8JS1kt1HB
L+KoxLO9d9ewWsJlbVXF8G5KW6cu0wTkE+6lm0fpJsSEJvcRD3MNNiFDAPHbaGbZ
udyJZskgVtPvKK3XaXHzBl4vDyA/NducCTY8H3j/+nc/phQdpXZDFodTLGc3acbq
FrF579DogZjg2LiRNyj2JDmNaUU3KUMR4Hn+Jcf24AO20q/VhlygWvUWpWweUrdm
Sx9JhkvXQyEXPDSaXIsbjMcLaQMZgdZmy2+mU1iZOBRAmC9c3w3fqnFX/lyYuaap
nfdoNrXF6AGJQ4esmLWxywzimsmjOH0kA1B+4BKowPsFawZy8pkFxPzarhBTIEOn
DVb2iFktQpO3rjAa+ToCSugcWsl+96rzk8itmaHz182bz7Q8TDFHkbqndRJ/Ayo7
u7I1a82aXOZKQy9MQNO+8VjavWtXQXPW/qZqr7MIR0CDLhPdWchJfLLSLLOWouXJ
xt7n5Fr8cmYzvzPjxKVfo2OuGJPvXiKlWhnInd5x79WnIQ5Wb+mG6qZC7bm+EZZY
Uu5s4ewLzH2jzaLH2eRkqW6/a9iV8H/9rwMoX+RiVhse/mF7OOCZ+Ewp2pl1nuBe
Ru88rHTTGmhOPyxm1A9IRvcBqyFQJ/M5VX+VR5qcVFDADCO94c0ocs9wrYEGEdBQ
wi5HWVXbCHLp3q4vtqv0E3BIloaMW1USQQcy53BY1RdLLRthOSmuma74ZVwrOazR
sYZ+8jvB1mhAurCdV5Sw6ULUBdouuhoObfWWz1sXvEBCIggQR1U2JZkhPpALAH1k
o5jjfuGR4/40pid/QfOqX82isAPuC/pKn4dxr7S7z2lBEGekKXe1LezYuJ4IbxQv
gv+GikkFi6fBSifeiIvJQXhM4G64r+109voL0mRtA6bO5LhCxvh4ELyLDy2pFhNl
auFKPfm7I72UFFWerB+OjOxfr1mouLLEIdLxg5VxOo0jiSQM4ePY4ceaeveaCLcy
BYf2FDmK1UgN+Njt36oVLHirMnQZc7S00MpnagDcodo0O6Hes4PZHT5wxOlrF4pX
/pLomMTvn8IqSuxP6g31N+0Eu66DkqYqGE+p/QG+YNSSWla749nKYQDyZbvJgqTV
maA2UHRN6FwUzuv0ENur1LZQXaussvigLhUrytw1Zbi+7jkfrPvuLp7hCpgxw6ey
tJygIDbVkDSsKNUhoOJPETrO1lLxKOO+9PrQWR4qOBUPPXsi7hDScTI6jjqERlJB
dpb7/PFw80SGcvZp2OIpsuW38sR5qDD7sZ3054phcuXzf8GcoDGa3jp/DTZWomB7
UVjBMk1vcleRSMFiwyTP0CBUIYX2vyx6CNTpmO/eNJgt1T+Boi1VuwiZvEI0Khah
NlUCFGBZIOJBvGiQOVbaOi/2hVJNRznTipZ1utv053r47a7sDxSeHeYh4JH2n8M3
6BHt0Y2bmk1ntCOVSbw09443y6GaDCb5mfzgcUlCjyR+p7hhdF6CDnTy1W2UNe+0
Hw3vVW6it+VcBlmrLGsTfeuPScnKRwkCHmgMUYLfXZWvC5gbbj+kDOo1Nfnr9+7h
TwvQZgig6FUFS2SLGwb2E3zCucKXWlkck2IiMNPS3GZsgQw8wDDzQ4uLTZ5l/Llv
SG23haREs69U9zZDLNPVOBGKz6DR+C6NRivMvO8VdWTofHeBS60HatBEvlbP5UBf
Q1M5If0U2Ym/HocP4Y510J5vC4Av5seUbQKIoY1N1Cuq0vbccXNrI1OGsvsMQSHG
5OPNhP2NubOdBYXkAB+/QoLeEq2dTTpN9Vo7R9vv3wF9zNof//c1wdGy4G5z2QRB
gPlNXa1KgiCf8hgfWkMAXEYOXa39ShRrh4MEea/g3aiKu7pLgXtMdpiDHkkfS33L
D7iZS+YPPUeVuD1oOyWdwZIPEpuAtQ5yc9AeyCi4iQF+H/XXDsLXRvrIyvosQOkB
5sao4FUhNqT8ZcyV1HmrfZbKJy5ktNN4/l2PZA/LNFASn3TWdpchIg4NK5/0hKZt
PveM9OP0aQcxjyqRI6N3RU7idVH2r0r5FZyJGTO4oBn5IMeABED9sd8FnCrfBId8
TmJouxXDx25JXLtl7n+IqtVX+f7vV5378Yvor/oyj2Kdc/Cvhykvp0hhcQiLTbPj
QZhmdrEVswCiXM8ARj74u5XpP3nOB3YouOYJNJDKB/EDiH9frnWdg2FE1NYB1omI
uq54MDYkvsrzZuFrx35MzovApI3I1TYVSws+a2dkT9SjBFp2qfl5kzWKK+JhOgl9
Kn287LP8/4htz16f8SIX1tL7ekMvxzqFFaCzw5d3vcNlw+7xvlAtMok8FVjRyjME
OguvlrGbHGWEz5ALmqbHPtuUnNOVhZ6N/tnSAEsmLwS7MFctu9Cji2HlJOMZUc2n
WpCSdMqaOqM+dafgJ3qlWYgvcHn+kRKZsEeZMnJXVvrwuGS0e0qGMrrrd1ggc3qo
qbUT2YXG1Bb5f19LvjhG9rx7ff6y7D8N7TbUGqRpC2pj03ZKY2EKsiGym98RwJjb
AS9Gu27xA/gmT0RmhJSIV4EbxJBhJKTp4gXSGwpaDGNCNIOc1uGP7zPpRRnMsZ5x
kktW6WivvOOIDt0HBQFUl25RWgjuzZ9VLKsJ+mPouU+q/ZhNIPsWE4Y0IcDD5s45
+nU6c3yX0doXIhoNUHBxaRwg92tq5NCKl3GNB97tg9nK00fBObUwTshQkI2oEGP1
y9qPB/UwBfMv+mV24z5rWYEODCNNwaTTSBJGt2yd8J7O+gZL5nnnK/YvztVFOVdS
3XauHE+zDW76tsGq5AGePmnHFN8IOx1Ln5E139bQZ4U6+wRAfGHKtK357bcsykJc
dcHXCp2wIw2MUvhVXzAxCu+I0+zkAb6yU/w6aa6MgUkcPcyvHRxoMAYzq++obLeR
4yuV9ALduFVszIQ/aQIQh8ag67m7ya8/mxyEY/44Lwq7ioXbXRvi5D0WJ5iJoMka
IWF8MLxMnZfMp9BSk+RQP1CAJy2MHAUqk7g9zhKdn4DF9EIDwl9H08+SGNw43TAA
/dCcYU0Ms3Z8jskg3gmN8awnQhiUed7z1GO5yjtJFXlVnWNX9t8+PyJ4lOLYXXDw
/D76qbAgwFWAXF8p2zq5gPHmEzZekyZpyMchiAFi180/Spuv1HRGS0Pzdj7RUwLK
J8hAXcrGnG1i6p8ipwCMwBjA9l6qRHJHkNmRfwV2CR/x7cZePM87Mg8LuvNE8SQa
lGO/qOtzaXtdVkUbqpOXg/HdqkP1AYc+KKd9KsVr1HzueN23DzRQZWez1KMA/xXm
unhUqZK3c+sUSFS51Kr5olHf6sjgoWdsd3QGR8G9iqRvOLPl5i0ZkmXKphMryva1
MRsfymOeh9KoRppUtwh/VoCQp8nqMvLC6ZIcWPav5eezG1sPObBuiuxcQz0dcbIo
4LWbL1nMYN3L5LFHpSL++EEpv0ECaj+kw+1BoJwFuNGZeilAqQuFowmHvq5q3MvV
zZadou8PY8YiGCLWBZWu6XKJW/od34D+hbIYa1Vj1nsAHQP0kWdgjYoC1AkLOxHc
TZe919FmZetUtevyJdC/mvNTbP+Dxzz2CxpaALjMmXWJRsyNfRCgX7ynJ4Jerwqa
XBMB007RD41ENBGRPMl7i3DqK3XarVNWTeI/wkO4gJWFjbb+UUJfgzYm1Z1UfG87
iSY24rRFUWV5mgqVuFptRbVMJDlhi2QLqVXrKM4rWGcQDSITk5VXanDCmowpu2bb
ZIBZa0FLcC0ReMKlslofKmSuxgvlthB2ZQI2rpk8bg+eHHiRJ6dOl7l9f0Vg9pWI
hGTOA0aQWA3pad9Ef8LHjce8vV/2fX9WzSvlhjGNF5Qal0fYm6/7cGFalxfK8+38
TiKSpotFJ+we9BLzlnv3Ydo34vINThJjGvITgGo5nip8sccZcj2m9/Ho8XJ+7ONK
wto546B2GlKGir6SiM4FPiW8gegbYRtAwwXJiJWG4lAUeEtJQVal7OwWGFMN7tYM
10lECj07M8KcyFyTyCO215WW21C37dxBPrpVSVt634GUkpeAPZYA/dUi2fz3NDqv
hdUV8vJUPl8mP5KBz/Cz8xrW13kXYaecmIWIOQTcdVs1s4qNkR20PdnNiUhorDXL
SqX5NwJkbO9gbNyc4eZyi0ezJ7Tg8OoPKSKkzVzCbrt22tHb9vJzsZb1tyw6N3fD
briK9Q6DF3EepusA15CnPd0WHKKOjvL3+b1Dd2TTd8W/MyCbjZ1D2K40j0qDMUg+
cnenSLEauEJHpCMlvAdGT47C9vYe8Y/0SIuKGwuchspW+fat0K6S0vL3PSbHajbt
j0nyyUGG4YpQDdcx/0IaL1flpSUngmY56Ck3k/lS58POmHx/PE7fQVPYowwkaN3S
zauD4rQ1IuK70eIXa5yHLzjpKqpEJ63e0BgegVdmRpQJ1QYD0FCVcUAzXiANyMbN
LEuPRLqQiNQAJszCxEerZRwYPZ0i7kwwDx8yNaJCm9ZBu28zV6hrm9su3np/4dHf
4oFkQVLouj+FPVz1Q0r8lW5xRmEtjW3CdJkmv9Taml347P9c+7ckg9Yl6e9rqQis
zbMpHnPi8PzJ5r1bHghssS0RAqFsPwEG6T+A+Xn+IXSgx9h7ihhpKgHaA73zUBgZ
7ZHMaAbiHlgXJ0lphpgM8MYIy529TqxrVRhT4g8uwDSBnYsgBnw5sR4mVwhrI/2p
uyM/E+Uh4l2SFkqF5w+rlZOuoliWSdth6KUNsTyc4einyDx/dMLwREqh1tAYCi1o
bL1DbUl4F+5oFB31aO7jDwC5v5yDSlm1ioH3a2+KzViQYbxABZooeWsVOlSl0fKc
I6c3jQPJPLKJ9u6Of6GOctPFMi3XgAA0KYLnEhAEiYYxnuwwobUCIKTKVbtczVh4
FkyRmaXu7u8r3tD+n+aSbDV9OByC7rloAJdVcGPe5NzspUdnhdu1LRjchoCF5rgy
tuonSUIXvvLWL0klaK95tHJ2NmWtbXqru/ajL2VqXBuLj1nC+Zd7m06+r7l2Doxb
ItpZ6oUfkUn/ouHs2EmLpPB6DhK5cEVgneyYiDFXcNVt2+DnxPzFmYt6KqmkNS/t
otrBhCbLb060y2iPZSgxEsIjLV9NJKs2JWM+F4GO/9j7SpAS1zZ0Gqm/T5UAf39B
hj1B5VrFqEK5slQ6FARuAqJlUg5PMUNtWhSeHBqZtzCGvznPRznzOR3X2pjcg2DI
heCW19dSaOh9fSl3XNZk9BDIav5s8XoeMJfaF3HerKksyLmqd5ffe/gliqom/2C3
Ws9tn4YJh2pTOSEItkWP4LfTizHOn4gz/S/O6Js0vVAQ7xwyH3kFmDy8HEIArH6I
F0ZGHjF5m21cnRbqi4VItze5cJjchZQt93k2NEX+Gud7/ULHdIULUbR5l/Z8c/Lq
ZmYbrOeSBya4kHw9ys3kb8Ay1KuE+kZr6yctgoFlIdlgKC2PYkSD0C41m0RxHOX1
YPtWT/f1mgPhb/EWbONssTKOS1xpVkB+i7MqyYgDaElwoAvWpjWGcoBRHdApoBzY
4YsuBkQU0qT1CbgYgMF/eDJtbhPWHBPIvo7WOHNna5YUmbZw35OU482PcNrAaP/c
PR05BoMr8w9Mos1vV+o91Yb6eNBE8LCJvJ/LaOoJNzH2/PdBSaLdsQkoZdC0+HMH
uGtjfsJuzToeTA6luSK72cw2SgzKk9FkVRpby/FpG5B8E69M3KcBqdAU+A3rVzzi
dCRHynvLYgx9oSVLlVQoU1i/E6zxIlx1lW7E4F8HMfeFsVQ8qshubNDTX/eBFtqd
JuYHNn6xcrRYrt0Z4T1/7rmwQgd+15Sr22hPwWdSpDP0m90lvg1/UMDmhUsdzS64
1HU5w93Z+QiAH4zmJ4XOhSy3AOt2j9BH2ieLVsSfwG7GT34nXGDGhgxYFjggJRC9
f6AKuhoyW/uQrk1LaQvVDl2gbXZv7KZUl7qgIPpuhvKOcVN4aO8+uv3aEVBlPHQC
3lwwQYiDNT/fDLxRvcQVj2CMSbo3BVne2y+SO26TfjDqv46YUIDqfPpV9tjV7ise
kXDxAG0gq1cszcXGuVGhbBdJm9EOHFnYcLQvicah7ScfJ79plAMma7dWYusCDN3R
1rMq7MtFHo8a3OnpkdNhRZF44Duof21OPq/b7l0OCz0LLmC2HeQgsP4Ef03QEyMh
oH30z5V2juPUGloArkHtip9Bipv2CES+X+8aBRdRf8MIMK1O34M9ElwPlPqMKJuO
EtZUTlv5Sre9WaCQa/VNZIwbfu+WwtkxT/oBcotI1cwe4yz8OMMjjMDT6HpH8O6Q
xrfOzQeJVyXcT/QEL76DGDYS8rbxp7n2V1PK4P0pg8C4eVJ6iIsHWPaqeKQTCzOd
vLALnU8roNuML4PcPxPL8/HRnpniajuJQTPnB2pgsTISA/k1CyUTGKnbQ3zri2mH
FriRwLWIlP7Xma8HhC4BONB4LCuZh2GW79lSctu34zDao+P2BiDPFiJao9AYE7q+
J/Jv7JaO50CWHXG9tAmvZcF3l4Nmnsys0Sz0maVnJHm550TRa7G01kcQN7+0jN7T
Aa01Y+ULjIFH7kbpmrgLO3xYnRzp6VAS1gevgfcbfstMAMPGRAjx3pClAfRhGhvn
C9I9rOFD0/FzUDe/i6ryHdNpY+EceyLs8VDI9Ppybk9a6Tuv419sfJlg+JHeJkAW
upPeemrbFXURHyBZ1Wpkg7bXhk21v3Ye6J1kReJRVjDoooKJHIRlXs7ZQqGuHHQR
zvbF6pAhJVfZsKGJgsFAbEctUmJa3rvgQG44UFmMrDCUBGsYxjRNr6osSaCq9CW6
4bOt0cBg+DBkMuFx9dFoOMpu+TKtetB43KHJuXA7folQ655yPOwirrpzAxzOclET
+YlEhib3f84kzIli6I9laTMm90BhnkNKlxO1SsHKy059O+z/7fwXWYtmooYEjmXM
qaRD+EaORvkzwpHbXTTIOXzDY3r8WFzxjaIqPnlnBiXiEzJ7y0+Uk5Thq5zWXEXc
NyGTZYhXRVC4RZAHcU7KprPNRNS2Uslaj+hZhlVftdp/b5sjfRS6FWYTGJvkh+M/
vQetyTqkEohDd88fW90wJ81tmff9w8RedD4uHPadlJaGDeSzAFck+ijTX6G8KHlJ
2fWTzGt6+um/sJS5VQVCC1T+LbRS1xwB+QWh3guraA5WXvLWEVKvhsAT+Rf5suZk
ivMtSemRc3V8g6Y0tRldrg6VvHvDbSsEvacDbuk6+XXh4vZxcP3kpBiGuQUr/Twk
yBNEseKaBYrWsbQScHG3PAaz0whFysqwnOfVYseOgjj8tECsSHlBOHAd0iMybVOs
PPMd3YF1riQz1J7thRPqOmNlZyLdRQDmf07yO5Y6hfMbzfWxLnHv/QDgff1ke+e2
Ypl0qhHZwq8dNL/Gq6cYklE/WEJzz6iLb+OlyWfkhCdHdAcyCWWLCnI+iKYzE1no
FMkvCtUhBDmL5m/vE2hcNF9vaBTfIiuVpcgcfbi5pweJzeiODccU2XWRMusdEu8g
2RkH7Bh1WhUsIUSLFyNUealup9xcNuIfsehy7dQB+BksEZtPSPHmz6I4aDuDgQLb
p5vUF5yNgBqoEfJIHSAAvkAgCNK+43rmlGG2QV18yptxypxPHccf23DF24MZbg6z
nHKcD+JWW6s7j1OoxSv1FEpka+pmfRsPN/SZlISbWO5ZKynyaktmY91HhoM4ILXg
T8wYyjVevClHSX2+rATkX+m4NPLFxGdvOB+XSJE4h54q1VufIczoi54L07WUKMh5
RwWapZVtgaPRJm+wTZ9nzJbfSOWk6Z2uI0pRDY/bt13yHjX8KZ20Sdpq/z8ABLql
20sbsV+oPDA8h5ZUuzpY2q7OMB0jbAfLN2Tc4r+vREwfKvKLrpK6bm6SOhrBI6u2
dghGr4S7Eb1uTUae/MusA58B/rOcavIiOT3DKHCPBzYiMW0olTEGDb3tyvJg7aue
yP08lTlLD3Bbxlq3CQ7Sshrg1sBE7WOeXJ076PdpMeKlJ8T6ekzvjkE+xMEyuoTr
M15vq84xqmE8x5GpKp35BXEmzQPNZYrASj0CLQxhaFeqLwSAsyWetsK6vbSVsnFV
UAmvKjcLitaSBVYonS0MqgQaiKdEuLJOF5k0ZtbdSyQMKrN4LfAvTxfZ4ER9S56Q
JwrlBFuWsQU1TaRoa41Bsv8JIuS6m0opIo0nx66soC2IC95d+zGrsy3wpUiInojA
LUqrJl4lzQ3H/vMo9dGsVsMvMUuksh2DSEdnF3HQR9/wB2XXCJhZ1lyApTOTuoOx
w653zpk4jP2cdVcXgDFwb7gV6SUZtmaaWfSWE5N39hvdX2QSfKnky5k07Y/Fj89G
WAdQq12DvkKoHprEEs18RlwGJXcZxEmmM2s1DH4gcwCnCCAN3de40hKijZKebDW1
dQTdFP3aqqsRBAWGgMhzF/xzKjfHWU00+p4aPzVWvVYMlnDhmqyWZNLIj96o1Pgo
Z/05s97mMYBhRGrXKwy9ljU7sAUOB72sL1xTC2Nusx7LdrfdJgHyho1SAPQ51/wD
eQXzvnKuL3JScGkW+FSZvzSLaZ6E9LxJh/1+tP4Rx7EM6kfGTE0oox/7WgUkGV0m
++fpvvAJZ6ELSc85xDQxkAiGGlXu1mjcBPocpsqwaknx60kIc2P8t76iFWAI5CUV
yZZoJJSjbGGP0B8vuzurd4n6Lm8Z/IphplaqiiHhxqeDjH4RYSdp9659apIM7zNj
rrMjEODFlZaQAhLBMN5NoQBrb3EszUMhaJ4m/DOCSz3EBwLdMcrL5C1iBLo+FdWd
C9Iagk3Kk8KrFXhR2mUrRKKm+cVV6apJgFtaJmUy9TBcR4HwUk5jv47POMiuDFD4
pfkhX/ypV/8gNISYxtDznqbzsqwq6QZhy5rKD9BWlUaQRazUuUTXSeA5eHQj8H57
6UP5figLANVNWj98DEVzbmqUNESR13U62JyAhNvDfYrXTh/+Ni0gGWXiXohsWBoG
LKEjzkc4GUYd7Qej/53Tbc0gw7HUsR/qGHbcx624RnACGprt6ZUnY9sM4/GK4YEg
6tJExsLxvsQT3nGL2RZcTASf00mH/F6glCdbcTmxdFPqvsloG8a0ASolsXX2gRFj
zQLT/C8aArRSWVZvN9ybXZcfIOftlum4J7MSS/v1ME+/ZZZfpqkMBta/lMxlbblr
ae+Bl4ibIZ3usUghBm9K+uCiCszoq5ECp5zDwBWwDtxQjRIVq+4kZXcIdXZ9WTek
Q/GGeyLenKBdgB2IJVSVHAlHINkAIURvUu4LDfM5cHW/dgEh5ALAthdBpRmU3vDa
LFRWkVT14V9jPRC2tU6zuGxlG6dFxbv5wvYf0w8inygX5TVw5w2ICC+QUsBh50Sz
1yA+OuibkmR9lpCk8WtlaMvI1EvlRjE23bWQRtK5eSl0jyEqLUu4rmpESnUqtNSZ
BJdTEOZ6p4LMqCTMKy7f76TnxEJ3H+yIJu0rBGseK3TG33u8O2YUkaL0MXHfmAod
HpJTrxKEfqkMHJz8a52meSUiLump5QiKRcb3aYq7sz2IlA7h8cnzGLibDdk9IOF2
59jrIJZ+maNzOBKY8q7tcQoAKUyvTGZDMLVsTKJxZgRDuywHB7UngYR27HjctVZx
KFm6mGMyok19u/UXtY3ZxnLx413f5+UmxTjTk8wRShJpbMyPESdVsDsx+c/5E8yP
drbH8JxccWzPIBWmctwY/556JrpNubAaVdQpdWvQubLIcjJZ9Q/fk6dVn+QMjD2X
G6+cD+h32sw1X9k+za8bYAbNdwK7kaPpFzaYI0TNA8M79THrlm0CX69ADTk/jsSX
/kBGQT+zOlPR/25OZwzG68hW+XHg24U5Mj86RsokCn7vdzK+u9Wa0bzp6rqrplgu
ysQgYh1poSBoMZDiDKOuM65fVZzzKg7VL345CkC1eQrxK569LX8LFIC6XzKZcsHv
vZMj6Dl8KaaE7YfSKFmubuEkB0vn3Jr3XyCVKv9gOA1b+cUwO1vmsea3GKxdXXet
avoOBYr2WCWYUJ42TPjHn0up4D8uGX5xqB2wqVhkk1qOUq+2rVu5TM6ZiB1LKaqV
aC4ytCTxAhk/sn47O/7A+VWygm+1aON6qh1emB41BCiS6IPUdMgEE6c1xJGwsKPP
/9WrdHlpTsCltq1ulQkd9cc8jE/yELxKQ9e5EGeybLtznMaXTrwKOg1A/05gQYgs
DF8lORSjGR+8iWordgmreW8GzF9t4JZEI2d7VcBUjAf0v7/AZ1pHZ3jbu/xhYRz8
turZWru6S5pJyRAEp8ls/L9GWSwn+D92StDY/cCmwA36JiftDAq5eXR5WQ18mWII
53fQtmzpsrI1WwSTdsWuSDA3s9Ma1mgAUHNln5B8VQDsW5tk5wgmbX9MM9uV7Eur
iBmt0ioWgUkGn5M6M0G/IuVMZR2JnXVtCfFXJuS/qDD94xqV86J+7355BYJFwVCA
1XyZ7AugIfOwuVSe7ZkoKnae4okQo8NeBjpOR7cKcqhTfnnSce/necbq3LSvFypH
G8AVCQt7bDF0WxnGEU8XqlcFe9PFUIIdLpDcar3edUKUbd5Wem5387e3GcYdVy9w
wGCWfRt5j/yAnXKhChVrqRIndj4WKhkPp6GsJPGH1GPncuciFvybpC5cShYIsN3j
uymDmGSqP1LxwtPxRkOWDQsgkPOFRe6uTk1rlm+w2WbQukIGzZA9T6eEKMFK68hF
/srRbvH4RpTDmiDFe1DjoH4LuaaPYUrMROkjvWjLqiriXU1w8ezgEZ07H8946l7Z
CAIrGuDXTiJyHAeoe4Vb5ZgbKbsj2JTS7sQXYyup7ILFOYmyNbg6gDKLUDi7+BjV
ApFw5M8c2wI+gNOtep+oxAC9mtuEtbqa2gvMRuwQpsL+fe+MqOgvyTPIYL553voY
iBsfEjETcCNiwA2VoIEuKUauBfHHU3bG/EWToAXI/U/+I7xUbVWLGmBEBfugwbwk
+w4w3Bij1OhXxKgBidEo1598oSd63YBosY9PvhCD2kOvN6+QYaOQxGsXcXHFSLDm
dKvw+eXHWJOIi1yxYCYZWfhzyop46L7GARna4/Kbp0cwUjXHpXFIDiCyHd9vC8Yb
68pgXQfSa3gHIGM51ITn951GgkQSATHwAJoma1BxTuSpRW4eEJYDKo5QEylGGhns
u9azT8Nwaj9YZ5iZJdG3qTMj2IAWmGQJmEYXMyXMoGjVNPBX3uGI8oiuREb6zM9P
QUcnht1PJN6LnxKfTWgKli1CYwscWnUK4AE6qdnC1K8cUe/l7JGWpoghKED4U005
UFTTtfB4VEVvXlLfc2uiQbsgSH9BXcx4khAmg7rJm0w9LZyVB8U12aFr1r0pGkZf
1kfgaX14cULPwtWLGs2UgKSs0agVCGGiSvU2Bqia0cjXh/1w6cC6KuPYEy7QAbDT
o0fpNAn6vbq1V5IT0sp1V6uuz1ilyfX9liXbYnaAFYEa3BKGmJ47AFByG3XT+Cox
vCw4EhEqQ6BeK6jEWjCE6chuU3SDy1Ov8WlM4bOSjWRMY6AisvP8wxu+oLjka0gD
nso6fdnS3va7prYNVcxc5ckTUSzhhPZ5WeXaiKt4h7NPfkdEvOgseK3aNGutku2m
V/G0kHErfG98CtWUznKNKbRqGNcqHHIcnvgAfDk+xSYls10Q6B6FpFP8VGSDVyYm
uZtOWs6StivIs+Cu6k8OLT7M7lAFr/34IbnNd988t1/lEWJzjPAYKPhYCU9oegKX
mH9S/1pwqTomgQZJ1CAmn8qqJeNIZ1M53nVMQN/MIpD0rjc1ZFcWnh2E1Va3FPmx
Q2Qk/TLqCBj3oOAR2zUSog3PYxhg1rGb7lErGoo+EElhFYMboC+fcEYnA3ItfDFD
FSl8icyEjGYYei7/e1lTKyd4oJkZR1t3Eoi7y+KpD5sv7sVQlyEh4gCkXuAcGyj5
jZumCO7rimHGy1Rt4LZI1WQQaBnGLSOnoMv8h+WSRkkJfrIXEx/lij5MeF4DumOO
0N80mpaQpKcKHfw5URWLsyl2TER3kfrjG3ebK4h4MlScctBY6D18rg+reLsWWiHT
ROSLhpVuSKEyrpzKBheV/mnw48qVjYNDGCU4OmD9ZTVo1nJnCXtuWkrtbDPC67pB
4usPzsQgwrD+MO0YiVx4hYBfYK4UC2wpsFjo6iWN7mw/2yDrNVDa2Y9WkRBJRXuX
RCzcyErJWx4cSIt9/CJgaSgTpk7MBwPTGnoaiC3WyOL5NkfByU8UQRhmBzb/F1is
6Ez6nb147gF6EBylo5J10vt+KX0EknJc7EzuvfdCdvzb80x+qzUHZhUMsSo8wk8N
UaWG0VBaiiUq6v3n5EOx1lwSXK/LGS8OypvaHtuvAZKjlojdrSBEpxQJ7DW80xpj
igrObgKLneCc1+zLm4MgivQYlnEbzsJCSYDrLnvwsWZBrqNQsLnlVWE6JCAsRiSK
sQVutsCR36jwavZUByltKLWgG82e9HRSA18KnwPjmlu2scUUx3N/QrGMOSC170FI
VgDkdt6y4LeCJ2MuzjstmE6k8XcfCAg8JpZqfJ5XGlMCMS9IgzByA+OSr/i/is0Q
7c69+Ho1FZtIkS17zqnUDgKgGcN0JxTaZh7v2fZvu0/eT3Y3UuaULR3y+kbgNER+
D3igPkjs+dhgAB6zTeEOxC3pFxzVxwpObRBnly0FrizpoqI7VWoGpY0y0Zc0Rvsa
UMd3gjDIwD1G0Qz1WR7EjAbTdAEwmYjoHs+cUy6WdnQ8w8YS1E2E4BPg5jFLkAaV
uZA8KEW9tQWo62fD64LayVT+NOV87wYoCZJYDjlz0i58mXXsMOvKEsIbeAa0R5HN
TlTYazT8dq+tYEeSZmmp28dBSmqUQLWx+r4F68eVAwazYgwbarXWCaJTTazjV9MX
gApaohBpVKGiewwxvNhkVczJQTTW4kypvWTaj2Mgu1v8L24xCmC5TRoi9j6RZ5Ri
BzeE/8ooaARP8OUhhMIouHqxzNlIq50TxUnqd7CKQ/Ozp4DHkaVDKoyyxqSUcG5A
qhYwukKR+SHf4SGrydeBLrQABb22wlPAjjmNJdn9pDDd7Mygt/fTn511BFtudhoh
EnP0KHIuUTAHCNsNTxXnpnoNneCCk7HtkzxGZW3ye8YnQktvFC4GDby7/lWeD8lZ
vejSWU3b65WVCimpDopKd95lYXMDUk1CVT+YIZ4cOYUKNxLRVmM1NjZEWNiw3FWn
4RGOsAxV/DNkguF+HgYiUkXkcOJgweWrJuEhorTY6jcG9PxWkuuc/EMmg7sbTdbz
38hWCX86ETGYpDQRSj15r1bv8whU9FDB+ookVg5LELb1voRlWJjRUG2LlAHaVTzm
o/5cfe2S7nqqsPYPDowDTeg4GLJ9hlxECzAioAA97FxHyBJHege3jVMBW5hDenkN
PLzarjbYYNDVz3Xu+ovfWK5d5VzbiXVGbKfrggt3TZhRu8B6COKWsMggOR6cMahd
IoWQUoalTw6DMI9TepxLfFWK8n3Ea6PKsP7RvrhnB7nKcfiy4ekAQyYI0DitPpTu
BxBXaKR9Alez/bGDTPLi16npxTFq+Wp2L/SfwnUmmJ0Z/pWY1NecY7z0wx3A+C5J
yQAxIkWGGEaZwL1njFMHi3DvdoBrlOy2+uFj7ymx68VwEzHj6ZNG48igi6cUoAPi
xrxRVUFnLtRE5lUL6kBogy3VMu9WijBR7u+P1kOocirDfaHLwQNSR1xNFCC9mQFw
StDIlcrre8VzSHkWohqZizIE8TR9esUKwfSfaNACkJ/5eCEc7t28KFGIGqps5K7d
jsSdt/irFZgX9WMwbX3quuJYD/AYgU0MNcbiaMZl7qMc4yRwrXpTQpUyTXTyVTVh
UwmA2qJ69e7mNuTh1akKDFk7o05qjcKpu04uNNz17keQ08dH6ZWrjb+XdjMAQeQB
CeFWfYC8V+VVxyMqpHO4qAVWMFZUfCINuIgnMHcqO5j38Fe2JHbGlKyiOkQAwGvO
2dLhOIYKSJpAbGIVpgd/LQaczSE8rmc+eRbnpziUG60MXjLdXoAhb9zi7BsfOSL3
ollr9S2OYezpyVuwzJI1apFKqO6CbvJNMySGCfj0A44b9MOQdhaX9LQV7mfymMV2
uSUDvvgT9/JojzywyHVOUZxU/jO4bf3LhkL2Mv3CtqeN/ryiicQ5YQF/ECAz31xt
eULv6neYBHF5m5mEnygOVjK+3IHBMwCdrya8LFr3FDm9MUOfyf39LiRXSM4B0+GY
GLEPW0DcDhDJ/bhXLaL5ScbAd9ytJ47ejthibslOZx1IhC4sMhEQknWaa/eLGZM8
IuB9us/j9tuCdl+ZOyzZPImkb017B7UFXinTRRdhUcooSyZjH88f0K06JS/k07xO
18Qyqc+gv4eJAMUJB/Svt3FdGGMM50TxOTKA+QgaXgUVMtejHzKhacsuZ7Bsb9xA
O4ahaPV088hT1q6lgmg+a5+g80o8fwGQwpNywxj4jVe/go6zGfL5KRZYM5/9xxAu
iurK76X7XhgKTd+YqQqEY+O2cLENG1KSS8IvqyoGJpdPRkBoi546j9xUk4eJreCc
MfxZzsADPmFmf44qPaOUAwq0wynMXp1+68QjlgOzn5YJ3nGmsE8g5659/qJQHvlw
Ya+3cdu98I0qCSulDLhcX74OZSoIwIgpAB7ljcBB7xyuzLD3Qn1/Kt1+HQC4wyqw
zgd/e6yxhvSuqFMpfnL2BHnroHeAncQ31BwxVEHStKwZZ4AntlfmtrjY9toFvllI
TOChZ8AProNzm7vyXw3o9gF/V7hvKYMWZ85TjSzlKMXN2OGsFp8lt0DS3XfHiK5B
z+GBAErw8seV+yagzf4n3w8MYN4CZ6si0RlYCKz7X00viMYBkydUyXhTLSao7U6O
i5cCWCRHWK8LdmLPnnG6zTaYCMUMyA2124VPQQW88eGDnWlttfrCHo+dQqUjyYMn
MpiaPFhT1mZfztNRYqef+pEEb5D+k5901V+6/KjaaJtvp4zL1NJXlmse4ahxQ46Z
vQRb0hK/+EPPbkoE6gdu1OmBrJgXG0BeOsqDunXJXA6QvHVrh4/iFAt5a1yYYVtr
Qc2c15ka4F//tuZ8SUjrvklbQfkaz9qprdX8P08xsAW9SH8vRxehSylA/FJI76yy
udsiQRCNBt27j+emViJAPyBn79iw77NACcIlacH1Y0H3M0JnNgE1za7sWzLtSMz9
T0JmTEYUrQIyvA5BALnVCFht7fPd/UbpqGPKyaS9Nx+Y4f1vCql5l5F04v5C0p6S
miNG7t1MuIiYd9Juu4r85qiICMZuGPeKY775q98JdEuWF5l1d3rFslC8dwpgB3TM
blkZyceLmGnKj+0Wd24WdkpPv/dAV4QBLIzco3SdP1ERFCocMm7fbhBbsFHCEKWd
H4A+7JuNsHGh2ibYBjJ1bDWnmuWQ1e0RYN6Nt4e4ABZO0UBsGrMIp4TU4ol5pOiH
VM4ATD3S6+XnZDw/rto/7q15D8KwAF8BoidbZS6pGECEryWStMoikT1hySAa/3b7
+2QxTEMUb1BPyhQLe7rNlfa9H+vsVz13rBCERftqv+7w2ug5lbBjdNnGTMK+EFNR
7dDq7nCffpI0yc46FDirBfzs+BdLnDhGtuP4v8SfbUCYH0ALYTDqE3CqrHQJEZWv
KXu5LqJcAC0O2qtm/gtRaa3QtNlLLdYrHQARc6ENW3EsFcrqHiCAPuWc31HMorCZ
rm0itojntIWpXcinRrqGwhxt0z8ylJsn559IWoY2Cz8bGlRQ6ywkaWKCJGG6mUxH
VlQlOwt4PpqgHafNfEuMPj4DlhWkzki0n7/MduJBGG3YkhZnV1zLCrpMZWZ6S3gf
X3pd8q2SUX9wjieVlBrds1vtXdZPpHtiICuwCpko3SDBavo90i/4qoXHVq9we+GL
AlgBuRrVBcLp6SIC/KewXAcKYoT+V64nK1iZjdy1ODXmVANs2BohLAZ/nee/hDmQ
dKTo0pHHxkNrOlGTB0n0ZliTxg8WcRYMVxUXqYgNk//SgQuipUoy0q7/ztnTm3ey
/ED7hvga00qBvmGu6tlJXa1cSa3+Mxt3c1i5gKp/X0zDkikf/kSUmiFbDRMlC2U+
Y2v0JZzQUz0bCRJh7PwvdIysxmavfzp9+jw5Bgtq9CMFNRPawQFiGXDuIWTp689Z
LGvF9cEOSHqwHYtWnBVaZ4ME12ZiYKm9yM0wf4JD6eVpsTc8Y110UHgmM7+D5iV5
hiKmVeir0fcLvl3A9GUVx803Q3HhJ/g4KyRNTJz1D476i4XfPs+ByBikWYR1L1vr
Wt2b9m4PJjB8JbuQPkbafBFPS8/ELidXig3A96X7xAlATuFxirNRLvmxvwOX+wQf
3fmi7rGGBEn9VuQ79iX3iXEjfxLrBVVfO+iy2gGL//YmqW4ppOKBA6g3UmJ1oRt+
Tf6DzyG2KAXa3XiSRqNpYNifS7qsLSdFgBtYd1HG5I8ipXn2gNGOr8+eJKgis8SA
uBHiTItRqzab6pLKwzpYxJrYfN+U5YsPk6NfW3rn6HDu3xepiYHTdmufrqhXuGTP
CbhE7Xs79vKrptpj2TbOvXDqERR+/T0c3U6E/ZCdmxAs4equ8gukF34eqGoEwxoT
YyITocTa6qyC/LsJ91aky3osHYLF6yo1Hk3XLllAz+bX5VZK6TPyC2MKK/lG4LcH
HidAj+un/IbIKj8g1Z0SwlP3m/AwYZ4R2+QEco237eMVMtUzZnnoR+CeU3Rgwh5q
/0K9BvXifOxD1Dkp6JP6wffA08OmExM+reQUa7bVdZEYRT016cmALxZ8xG7Ps/gH
OQXTmEoYEaEj4ElgW3g3T9SclkSVUrzpBVuhg5B9CJynBm7Y1k39ALkVjsmskyyf
6RbQVxl2IGbXvWLGv43xVesog6PRgYiG2zzziIP0DcC/XB6MLPaB0PldewqzqEft
Q4iATs2hYtkAyMFgtZSngLiqYRoq/hyo1eU94yDdHsC/Ta22vXUkbgCV9I+zY6o6
VbAungmuqLzZ5pR5BXIpb8W3YRBB4B0fNA4AsOKCG5fKOPoFd74kcjiq17NWPbGT
9cVn1OanK560DK/c55l12V+vC0GB3OHA020/8W044PnML/sl2pojUg6eDzN9lzlW
XO/wIXVLf9uYnG3ch3+/v6mfOj8ASu7z0ZKBxf6iX6oIgHbEvKmj9wNLFA5VoBqt
AXJ5rI3fXrOSL3jqCPgOCegwSKHfkh1HHJYFIxt/RR0lko02ZpB5xMrEo0fY7O8f
ADZh49LXFf6rioz/Y123KxGFJA1LDef5wXYL8PpY4iQMdZAfYvmRpHx+03uswkNH
4zjuuCSd8Q/bvovQGAvMLZR1kwfcOBGmxR6/Mv+XP7U0FApr8I9j8/DqzRRxpPSK
6dCxOrehNT66czfQoXJCf/InCPM17UyazdPjEUMlS8m0Eaa3obKAOD6OBwJ0+7KI
6X2TlhtZkLtiztW5E2YzDzSxxgPLvrHyeemTHXbTz5nF5BNQmedj5igZyygsr3pV
H2NeriYm1Ts8D8StRo4dPo5/mEcY/mgZ7gZHAE1ax8lRR0Sz0u8Zy72I2ar8qr5v
LZjGeND17ILkeVBYoWeBfmErGOfV9+N+cWQz0EJu7/M0wyoSpj+q8OxGeQE68Mqz
jLdYFbqcOwuAjNnFzuYfkoCVZke/3kLlTu52R/JQLYe9XYPxz0M9DZNW3GA44D0b
2d68eKSwORdpJFRBgAIwGTkOHByBKfvrnGaioEiNH7byfezQ+ItqBVF+OMUkDBfJ
2THTV6CdNYEITVZkxareSBwMSw+TZpU35fctuXETUle1wKjJV/kw+IwdXCHXiTD/
wuS+tAINZ1DvZdLLN7b+McwZdPtEF43ogrw4fC2igfmQq9+HNKn/ZjSYqPxlSUj3
qcaL/j4ElX7+CXUDGiThGdLwiHEHGu6NTh49lypeJYZlf7HEcQcuVzN/mrVvyxx4
ho3v50b2ISu9mHUjKJTePVJ5Uj8dRUynxQwVczLYWUo4MA5wt8uwCqSG4CutwuJA
LDX6Hvv2fudoeqnhL+SdwLWHDvzgT0JsbVa4+DIZMYw3UvCTFAx6ZHPEfJrvw1e5
id93nF7maiWG85yR5cVQlG5ucp7h0MuDw6006kwPCXMQdB1drHbOqGjrhcQ4FWeg
vEuPW0rHc5viEghBnUo93tnOBF7gGO1LymjyN5Rp6weWVW6uGRdCVcLeFFXSQ5OV
r/9QeYUtlgPoE+inyK9i8N8EEueP789UATU10VthB9XWl9WHAleJmJFQ9Xrrb0LA
8Yq5W/jqsoZr/1Afk7zhmKpD/ec0UVh16QF38twzW+XWSi6xchCjjCarTodFoHJ+
3ovlvt619umr4/oZO5EA18AOZll0fY27ohggmJFfarfDCGG2TxXhPBwx8iGA9Dku
+L9T4SwyImz9ChmLGIiOGtoQSRUWTqAWH7WHLY0CztyeqzNlWO1hYV2x1wkankdb
5oDB5NFcU1xb/moJ3RXXIy4C4zBKMLhyQcy+bD02ItVTxXuDTyOEvEr3es4gvqk2
FJIT7eemvbkFcGgafsHOjvTbJ/ECX5mPbGUgReu4mhtjxTGwbZBuvuR/Xj/xlpUC
XJB/OKD0JNSH/gUIkRHD2df99xS1tp47r7dX2bu4EtRD6leYAhihiE9x2dsZnXHE
XOnWnaSJsJDSqEG5f5jtnnHlFMTILaa5rz/3Vk/muv8CSZuIQmln8hK6pX8BXijZ
wQqmvU3/4goCNmHEtDH7D0cxf14QIm5I4xXDNRdEwVdZWHWHQfhTm6fW71dJ1lmK
Tf/IPm4xw3AwyEPP00Rg/x7YjUlKIb4PB4B7gfcR+hOe0eujjkzCoQRuKPHqXXwa
c1E8AdMPBgIofCTUITUfpFNyq98xMR0VtQc8Sf/MeIDg3M5bwVNG02pLgrCBKHw+
vuAc96ONYDFWQdYCYVqOhQTiaBGcKUNyIY3jm5SlMgbhenXFOh54nIWnP/ZIcuk9
rGMjHOGOPGx5TOwaIM7lCNm9BfQqcAXG1fMp9Uu9+HoZ9ptYhKoAGFHbEmoGH4uI
sU9QhNf8Tm1NlGtJX+xK/BSCvUMgO1wgQKkRZskw//0TE+0wtXsVxdzt4wYhkPhq
UOICfC6DJU1twBVYStcKDOyoPnd5nim/YF6n8H+dXmm3ffhkC+mK9l3nJumQXneG
un0AKq+12ptMC0cbToiBNt0LaZKmAQN7a+pnp4lIOEK1pwKDFVm4wO8yZequkzT6
l+Tn11YUa2XVqaI2Pw0aUMl0FQ/DhwMux7qC+mj6PLLNx9N3C/VzDA+rHZv/cXC1
EThNzevd42cGx3HR1N9m5ri7giRjUPU+UKMYR4HTTtmKehK5Dt1+3p2giblYxsPX
5NhH25BmKWWJl0EsUmmORUQWRZDgypgnBASVh0ePz6CoEq5nGzfbaVsV7lactIUF
Ce3YFuW20AtBHHGx5NdC2Ka7b0jFsqa7P/fqdwJRKPXXEXAs4KSKGm6GN/FBlUQ9
1YkVcNaZBXgrF9BDmzDjCCXJ6Q2qJdme7MzSDkGanvQ1HenrjjxmwyvpQGuDOxe1
1jJGjSCmvR7bObXkQs720p1JsDn9UJvllzaphbGUhAYdCuAu6XKcU08JsdEzWBbZ
XXsdy6kSTLzMbOd2HjmpKiQQpCSahXoFrDiEO8mCPRQfCPx7AybRky00ZhxJtUZA
Sbh6UPcJRBL2TIOF65JO1m/sHYTH8QtwUfyNnf/XS/3UFcl6pSjvmvvOch6ybJ+A
V7QmeyWxppPuAGSjjg5lmJx0GJgmSW3Cme87PkYsRFAvSpaPnWKdj6+EhmSU/qW0
CI/EWU2gY8g7XfEPMvSKH7dKdULWYVnTHGGcMIQKVgiU/+MK9P7e901KtpcTFdN0
XxfyX7ct/zQsnuB3DIHLuB5jUrp3kyOy8sSrO40QCrPmOgAfs39SJz8VFvk3dw5j
H2EgW3NAOX6u9LMQHc4dqFni/l3metDnXD3iAV/Zs4TsdYyq3Krl4mPLuGXkr+uU
gLtJifkS+EOvo1MwWRX7UvwRGHs7va6rhXoMNCNYs7UP9HsJJDnXMuf+tR3Etzmh
1bH8kO68I8B4pimxnHuQSUEp2FbXDnl4PCKSiyp1H5pjg7Pj+1Wo1gXsgMjs/Yhe
2tkkqi22u4RkuguVK6l0a+yl/wHOLWcX9VUfFPcuZ/WPe3EgztGtcJuTHfY9ax/2
4pJnxfUH2OXdeY8ijjO3oZ2NdUUVzXcg1HwPuJx4RLsWGZOD+ZgU+oImGE2TBILO
oBxT4jEUoeUk+mgFAVCGJnxSW1wL+hDthsskYpTshMwEwKow9zFSsE9xxsR+rzOY
/kpkc1u/Q6M65G7I6GAQbdRX30fUeX2F0ypVXwtMiBPXZeuD9E6CwKmbhIFbhMUM
SaBm69KpP0Ih/RYHcRLfNO14kDabG54Wiyx4MwAON023uLjTG0+wXkIxH9tYuDNt
mtGk8phwOd+UTx2rgeIYVPoYbkDPzTcH0fxfUs+YWkLq3Vlz+GOegoOJrGNMaELo
Q43FZ+1kF3izdwSmoYq6w/bPyfKBwAjpNShx5tSHotEHrKb+q6+EFCoPp5Ttx2Tv
dPw6XJCDdzYW5h+QZbebcwasMYgRK+WGwCtAeDRiQ0+4GJB6IiV/pSC1oWiLcaOv
2mGJLJPNYGBWa0U9yJzG/0QAolqQ6Rp/L1X7Q5RyKU5zj3tVpaCzUNt2tyTZ3+bL
imxT90Tk6EAzrtk3P2iulMDE8EtOeo5oBWKbHth9seBnBWs/YG7IZYJI+xzMKJwt
Zp0rveh9b6i5QRrPALIiry7vnNIsygHsg+bkgAFa3rlmwJNFSP1mtz0WYq5+zl9N
OsHzKw9id6jL9A2IOalu4ZkF1jZMPEqU8ulMQiYMyIgVPk8o9KlfQKMgvThm0Thm
CdRN+uH1J47eRIxRjdJ4Gna66w3BbAOKN6ieXwcaPiyPFZHgMeoulcC/r+zObue8
a6gMujinUPn4eDumXyzh+0+uL0gzZwv4PnTqDdFMAJMpyMVB30QxKldK2iws/D1e
Fup3FHIcjl+oPc1mUxwHJ8HEmetpx5eqHWWK2onWcma1NRmpWBfGJLIt7lfVR4EM
HZUCab0ys2MAwZqD5G97OUrUzWmJnEJAtACO8moV9LA/1mTgzexOB3elEDxsV34E
f9pigG8kIIAJHtC3giybySngFQA8FXIUlgOkUMYU8OcBSRzVtiHOuVugICvniWEg
vUkFhXaQaU5PnvHxthKA4PVn7ARTaeh5A5guMTERmHjGiXzCNAKELzMmW/T32N+N
lNBD+ZCBatS39HFY86DcrpuHtg97hP1qDnHxiMYx4T3zg0J7ic6SLmL2JVj/sg1k
cczp2sBQCizcMeirWeC2Ss46julqAakAguYtm1FhEzLPQsvv3KTgEFagvhGX2EV0
AJsZOxDsiVpV5J4iIXI1c0QkkcOwDaRmIZL2xeFRcRptIJU1CwUBzTA0QiVtSFUX
soQsJ63Q4HplzqMdrUe4sAeLSWF6jKppXIoVPQxK0bHS/eU1fELBUSqEmfKtDK+N
nz35VEvy1EUuChzBWLDeVp24Ef27GgIMVb1qdM9LRlvLfNI5KAai5w1RUPmjSNTn
0JlVSDSOISByMfvAmcoQ/P+FYpnt40yYAwZ/76CkGQFqrGeW4S8Sl6xit3yNJQXX
iXR/EcDbi+cvmmQWChsq8T+4pwEDxFgvAkV9A/rsWGUy8tF7bRif0h3dtcRlDB9E
k7pZnC2Lko20iUsWA88RyHYMM+Q1ZCE42NpJMJwxy29HCma8mTd2zyIWNwKRPOLH
meEUmgdhTaOgSSzC95iLgYs1aPqtndtCa9e9hdsiunDwr0J2r/zjbhve+Z3Xl8NK
4ed0b2yI327OCipCrL31uGctSjc3NAtqOvhU+BWVwNKaPzHaTZD95Ekf7eMu+B3Q
4vMTLYFr6CEdnjTga7xdaqAyd4PMJ+6M0tWTqOnqKkpOSrTa1MqqiCKnNay1PYsl
i94CbTyb2D3m9fcyBrHP8qabGMudGi/aOcKgiCHj1tTbO6oNwjfS6aTW2LpnYqSu
r58UnGa15SkCDEL/KF5hihbYhITk2GKhTVQfAv+3HARxmymVbMaWL2xtp0w/49q0
/gHUxAa1QAu/jcCmSA5xZmCXkkVQgdAeKKBEb1geRA1Jeu+wbTzHObYTvwww8RRd
xUor8MWSTbUZJUhFp4C/uSwU+L5tdFmiqATM7UnPtHEi+CgTbtiXhNPG5NsLh58i
2gAT+ecTgPsBmPH2HghU8djfk8tt5MZjPQPf5a9+O8XG6QrikwTRxZm9nYZxQUrc
gmQac6D8pUGGNGO9cAUn/YYowWXw/TGBIxcvgqN0DCuzZjl7rI30jqv5CNbSREDX
ydVzzCEh2EEgcj6vPMSqwvrvw9RmCCgkZMDnmapDpwSQGsetEbjIRk9tchiKGzCr
9f/jCDlaCA0HD5gGlyhuODCFbn8n5rqj90qV02xadE00jC2qrfdeoO+Pngx5TiUN
GxIrdkQgamEHTA7LMZoPYl52j/Xs0SEjAxdTau4gYBlJVJPwbX4SAC0wrXYdqpxD
siqJ8E4L5kq9KHK3vw6jlbYgGQTzcXvWQicPjNF3vo6wH0wAzioMHVglL2vNRofi
PszPU4ArCqDP7CPehtEdGjzqpAjMh4xvpVoycdMIUgOYaFUzi7yG1J6RmVq4Fr0q
4aq2gQD251ymgTf1btmKcvtSRwajkcNmUSS7WtQgLU0O1swgJiiKzirRlgERWevT
3BzBrW3O8HzsCCB2MfGcgnRnQGTiEskWkRr/55XsEidLMm+tyG9R/JptOps8C2v/
NX0iygMWwJZIzscPLKvw3UwHf7vBllGNSGec9WPRKaBnjWRwotqbWxXVTn4fP9By
S9uyFKR5t5sl1dQLOkK8NZZjrvb2+yxK8y+cqBRPxfecHi0aFgXxx0PTL4NjNleV
lH9rREr1PEM2W5gePz72zyysX+3SvrIJDkYnGG3pCC63GTq/uWUHg0LwYq0utvjC
BMF/vEG0UQ4kxfMgpPFhgVe0/5ME0y24gPuisrKeb5MFlNgbehW8dTgRTsc0SIvN
KlKTIrjp6MzvwroX9seZbiKA8xzE3DvapGSTS8hNZdKiIHDBMnkRz1FJ8qrYmzfz
rWY1BPB09urtYuMEn017k1FYp+MangISPIfo5EGoSP+x0yap+alWIU8ymP9crq7p
73edmwk3m/Izr5pPzehLPrScr5l0WgnMIMZnjP3Bpo2dYtkvu/PI/+c+dorb+wmn
f0J3ZiKPzuXWJGmLVdS00L51guRFmiYhTXyTpmKHTCMlzVH4oqgjl4A9BTIfGCKz
KJW/OsyuliQL1kPjZMJhZqpK4i0ca0AsIwvV1vED7Hx49wUl9osxKpYQV66QJJUB
s6gNGKlTsvYR29x8FoXNIHOfDgNjUDgzDLubFny+1u1vkfLxGZXVdjedVeWOXIgS
/Lg+F56e2eUjykwKUr4zYSY5BGWkU3A0RPvsliGovOsuKRCNSWLE3jAubWKvoG/L
1QEtBwmkURgAse/LNS29yvR3wwK7NbSAQXznx72F+wh8E2CHr2N2avMWFIGbFbzR
6LnBUTCw9sCSWUs1Njz5+90Q89y3P8F6bSmjOfnyy0VaKJJnjMzmLJ4n40nlj4XI
kuy0A0bqPPtlsZQEXhM954qjyVTWhROC6Tz1grnSQY0vv9gojys8UeUpcDIF4ZA7
0wLLEawl+GBe5o5HLbBrr367XM5+YqyItPOQhp/oOY74RtsVSQjc4/hes6qqA9RR
nf6pKkKhWJEygUW+WPsJemxED1RN1FfsPjA4YX/HLG4PZIIFsTvp0Q4juQlNj5su
zLmgMNGDyLtzrHMwFE8fFvxyZkDXa8TFOcKKLdaeR8VdadSpOWEjhz3VYf4gtcXq
eLVM5kMZptpNBj/l9/+IA1Res/jGOZ0lqDuBhrp3iZwSZo2Dt4ezN3FhV6TxmiRC
Bd0nFL3MaPDpwb80jIsCI1ND715abNh1doDgh6S4REaRaXZcDaoDR+2dLboRC+eZ
Tcn5jI06iBWE6hrSXrWUxMxAFvU6nx0eU1FytbvoYE9kAp0HGDeRdWxSNvek00uT
G2dS0dCIEp1QVJpZwl985GtPmy3Rb3eXcqJwEvrhqzx5D/Gl87zbI/glNIZQM3dl
3Z522lgvEZSU60thrBguT67oMpRfHNRGc/If6qR2yn3TZS5NTspacQDJV0CNNQes
2c/wcF1l9u+0uYeGxcbo4k/AE4tP7R5d3W8dJy8BB/maSwT1nQowTtOG7TlkaNDL
F7mt1ZcCl6BwRrc1jwVtbsFpQbJ/I+RqhDc9c9yygMETfpg4ocuB/uwYpoX+g6x2
Mw37ETS7gBNYwp7+K+N8xwAvyqyqDj+YCzKBDSx5B9w3z/IE6HkfVjKF/I9d9h/q
UF2GIk0XcJeHvKAQF/N756tg99+BrysQg0kmTxyHyOROl9qIM80lUUWxKNFC6n4Q
6pVYJWczVFS0p/LEf7txwfBv8o9NPBMMKh4eNyToGdGs/RSargTVoruwpGIJb+MQ
qxCkGbcq8QUEfa53xLjB7GPKLsypjUDIwbHsHEDd3AW9NtnjiDmng9slAviMM+7u
Dt7vOtp3l0+HS7XOu+Vvbw5D7S2mKszZg9zbJCNZw30sZnXhflPNJFLJar1kAyB0
ZiKwmZoX/9QDaWNzknxiXkLUhnwxv5l607SjZgrzGE5v8ZRv5qceAoQViwqPJ+lH
G2iWXalZGJM2R/Z3OUTAuyXIiR5MHRG7wTmwO+56/YrxzNC+dhISvQ1yu42G132C
KwyuEmMn3bEZeYTvktUwNa3oqXUSeMP0oDUpQbnswHh8pkW76dOnHRXPsaSxn7v1
9VoT64iXms74fC33Sd+akqBc3Vn0jAugz3NK5rT2GHU/I+Arooppt8wRcBfHfY7O
DgxbdGrPY01egQxnLz3mHe6ijOXt5+b3KfVMCjowLuLlmlY2tGpcMC/sTEQlfeO6
mLeG04Nqnll6o0jnqBzWL094PK/7y1Xyo1IblIDECLdWoz4N1Vigv1KRTFrGQptq
IDux1avh7wy3NOp2wmVn4ywUzgs5OeqJuYXZ4B86xfGK2B6dDNGmJt/qfC0cCbVa
nUG+iSStCAieFEYLEC8eWNdPSNZfXS/nMfZwUIDQRu991MS2VPprjv14oVlf4Uqz
CC0N6Lgd0z5ptBulrfCzr8vF9U9sBBmmwIVu9l56o10LAAOMJGGYUjZhvlilq1Y0
SBWaPO7GOiF9V5HoqghXUL8SdmkZWXDSFHSlSXrp4+ub2FJcpR1COLniY8ORZL2L
FKBwbvRIQWsjOPP7orzHFVnvQvsvBIoTUzq2JBCkc7FR7n+GiCfOYbUKgPZMKjCe
dhQBsbEQ1mKUMCPp5BBp75l2WgNHZ28mY4OWfPRj80pGB8en2T3RyAqrXFe6qz86
P+X64EPtCyBC7KjJNAtCDu7Y4qiFwNQYSDljcaIVpMHQWbsjCjDe4mcH0jkql+eY
OHYUOkzfjipFI6H+t4J3B4Nny+MubNftMFVqot34z9XsSdPOGA9GzzB7TTnVflT2
Q7SHrO8nPaPO32UGALnoDB2XHd+5ew2fu7viDZ+QB61+SD4qsVf7mn7o9jpgsiXF
5nwU7BzLLDAARdnOuJGm+b/Xyzu2FMGSdpCdbrY66lkzIgARwD89tW6pwWPeENWU
5pJ5eGvrFv/LOAHHj97U9b27coO2klr9s641J0ii92mOi2UDvygS5tMs8zUb/crp
1YYLwqV2SnBgNVPlQ/B7fZX/tV4EUHNUDALfbL6Vti5DNa56odc2FVOq23Zsp73D
4yJehKB6s+jIHIwbMcPo2sTcEOwgKLRdlRa8Wm0DU4qTPOt9reUK+aYxc7mqSURi
ad1iCu3M7h1ms1lOJox0DMhNWieMy2ojKPHVRXOJXT2Qmcu7BCCODRIIPU+FcKrR
SiH4H7+ga+pY9P93ZP26PKIJaCep38iUr9L4TNTQQOhqzenNf0sDVASiNAINajSU
PFiYCWg5arwDGYYDEi27mrYBHO7GHn+xZ3ir41Ert4P/tAR1XB872jQQTHU/cDS/
96MnObQ/gVopctTKL1jFf+EC3Lgv+WQOx17BA3dynRgDFfAMFP3Y4uD1V3W+iMUy
+8NykIvn8j/bXqYEGSqVw3uDTNl4C3pn5dDYHfd9i6/BOC7UM1dpTSUWDjSJf2XS
XP2Rvc65+Btve+C6qQlKIW0DQ5ntVJVv3YYSF4WLGtEJp40BrKZcXYCAB5K0ebHl
An3Tcg/98jANzV6xuI6OEXvIs/p8MymIDkNCo7PuBQhJE7ZLqCLLys2XiElN31zQ
3wBvbesotxexgI8F9UL4XAbsxfrhfPc585O+iD7t/kHWssOV9N5ospSrn+uAU++A
viI63eNNCY/IB207KdvnLrIMUChSbElCpaU7dqj2hyGMZF40Lj6x65n3pe3Xckub
FoLS3WI0dNOaTumzDaUcuKxn3Y8YdDWbsiyAJQiYLZMB+WUSXDb0pnXn7X6TCY0d
CCDfDgbnhkF9od5A49G5wQJTmW0xm5sgidTt6lEnpFonlOyXULcxBPWwY1vM1eF4
adnGfiOGPp47SW6mP9Dewykx6ielIdnMLtjRYaR55JkSDThe4ZHkdSAk9Hv1+RAi
nFvo/njquKUgqo5LUDaDxU3MQS7iDpqhSIN0mEk0OZANGGL69njxdcmOsLDsF+Oo
UqVGZGtwXM6aCJ8ke+294Rqkf1I4/gULynCVW6lEkm5Phh+1aOQL33HCg4DdMEcK
7sjsrnyi904bdM8GPo3obqkUt8wodAUdbUgF/ylKVX+wCTcaQQ+zWbZeTqZFg87+
4jR5DYhW5wTqYG+lOmtbGuUIOmDuTdLWTMzKL7vCtkYXKFgByJqtoxAuRh2R7/TJ
xgo9V+6+QH+2DoX9lOgXyeD5gYp4s7AXzT6tQwe7oU39ImwMpQYOcoelu4CVVW+x
Vhot8A3x/eLVKGI4dRztgHmE6Ka5Me5wYzuwsm9eofl84PCGslBwhE4Syu4HoNaN
R0MLC6tsOsuNRm9IGNHkbtQBkkD2CX4PpH1G5m+28zGtIp75TjHd5d/lSSc51Jjk
QBynKUgTC0NvmmdSTF7DWvgtdEwUaVP/umU8vUNzhzZPc1yy7Le/CORP1aigYbO/
hnojTAEdIgNFqtdRDCSr5Ph+wnaj7+JL7COq658L8BuJsIAh8uuy6OBHdoexEhiP
HU45UoDdIs+8VDmPwOHPN6lAZWwh3GswioXFQVaWJA0i0TMlpxfv32o3kxWvQVGX
h6LfDxlhHiEA8hDbTBAyJ6GSEvlOgYCkVf+VsqDS0OD9ARidN5+KiiVCpR2vPx66
drcMc2cQIz7oa2UkYYbduo/f0BOEMiQwUSxtvzjsYOj2KC/OXaSE/x5utGAh/QS0
NZViXCETnxyvkSEWLeDpWDAzVaDXjSMkcWl7r+kA0fgnp/wNtJT95Ai2V7I3Wjsk
Sj3GVjF9IbsPEDfXjbUKyYzXgqSnTAqRUy43HnnJCehd9cZPXg/E0OmO/Ka/ywcP
SdT8XD21X44CHxeMHsQ8M42/9podNxqZxDMZgBzxGvQaJT4mjjBtrJ6KopvNbz/b
IKcPqQTJnyMQJqZ3fM816WXLuKwvunwA8spkksDJ7vcinWu0Lm072ynWNkoKVP6X
VjczEG0lvQOws2zwttz+knA8ywpjEoUzUpEb/S2DeoDFAlva23XFxz366MtCpEKR
2bebYe7/LG67U8NyX7CZX4MPtxpwI4vpAN68M3jg8veyaXYb/ffeGYibNpy8X75B
UD/LDbQI470uAxU7hu1dD5NAlmQ+AngXXkZLCr1QJiDzrNCJlc1fAhOQxaA0fzgx
fUInA/xnzAylkZAahzeLHNYFfMDt3vjRCZ07SUOPIIPonxrAOqFxgYhdQ/CbZx22
0QJ4zPNWIxvyUcarkJc+8sI/PD8fFxnJANH7T/409pnLyLbEwo73rJ0as/iTS4zo
rGatlcUga+E8T2m1uexacRYCgtqt9yyHe7cnxma5OLmXfVkLV7EtBQjok3ZFqDSs
80gK4o0J4ArEDh/6JBmOSpxQCb3+E5LKg52m5sE8jBpQCdT3OUsRKkIhLDJ7AV8G
6vohLJX30k63MlUC5+aamT8spX+LZk1UCXbP9VSyHD2SVE3yARRQVXD4BXpUPMMw
DwWTMsXsmX7gchucc+qVoAaOihemCZH1TSSdQ+T7EwORfu4PMPdf3xk5uc1B12lp
b3+pNGmhv7l3gJZGLcyiNXPnOQL4hwWfT5i8tQrgZ8YhMLwg15vKcxrDreVaSjQ0
3+QD0O6EriTf1gh6MEd+Grs5OahZmpk9fCyXxObCBsRwHm9q4lcfuwiP/gZdu+5Q
lWy+1fgyjj2PCv0PFLM3FG0JLABTXR9Z3XKupkDCmQ92W4EYsuGBGP5VPnkxUdq7
fE8cO+ZlU/V7+lUYqSZ0NuEE4J8PDrNBwev6/zSNLjR8ZD5nY5CbbcAclaHjLHfJ
JCrOXdjLICni4EVn2MXTDT/P0a5Ihlk/GeWM6XVqhL7R+XewIdUZYZmaxKn4Qift
OrmrgWrWa/eLsiG5Ed+UB+uJWqCX7IPu0obYsYpezub+f84ExrmlxWo0TS13YJHM
T+tvCjOU+0t7a+7SrxUwwfV/Bv/rqUzNTAEYnCLc6Wb3Tjk+PYPLoA86PBa/TOos
T/8vQmY+laqA2ChckFq/COdQLtdzZFuqufUxKMLubPuwAcCWJeEQp0g+yjksUPDL
0EwECI9ChNKHQgpzwpPBIlqJWK3HpKbOdB50MCGHpbT+YS/qDw0EMXg/x26ZctPO
taXHlLqeO4V2Nb4UntX3je7VN3I7BkjEySWS+yquSU2sE9YlQK9AFULe898fMeMs
Yn/WOUaOuvW7EX6yAH4eqX6QQP5PUph+AHt7EMV7X3IEZG7dgGYCBW4P2DcYn2Kz
R/TP4UDpuX79FisygYwNSPSgmlO3Hpf/myQL6yFZ/8DvpNcqpq+BuuRjxjI4OYxQ
AzWs/ptzn+PagOBPGz6kJHRikimWYq/NNCQ2T1TzgtyAXuUmx6I/TOY9L8NOBOyR
W7KkF9gqMkCh4tGUPh81ANXySWL0Nd4RqxY1cxWO4f/xgd1iFF5DdPbdEpsKWqT6
uSQRDt+1lbCBXL4rwJ6TfjS/eIurEawIiLf9i6+NmzBiWku+Thbl/yGgUmmCIqmX
gI84Y124jJtIcnDrPMXGqZS/PN8PV+xVU5dBvn7K3SUwIWJFtUfmoSxVzRA+E5B+
oGZk4st4QxHaGZZ+rYkhPOFiwIDNf5Mn8VqOBIiCsDeVpdxtuCpAd0vdYcD0hyfU
ZO9ShWRzEE4vid/hJaP7uvrsaAOELt1Xub6bi7ZS5gPoCFuzjGv2MrEsekWe4qPJ
sk7NGiy3xr4Zdxd57yUPbnYP3iHZ9Hej2paLZUn/qCpHHihDSV2sYocQl0kMGJ0B
xiPXCn7sJOBKdf1mb09BZ7olnDEIMRVsmpE2gCEABG5oshVrpBvf0H7lpaWhwsNX
FbM8Yex7UE4XNtxnON9vCEH4F011aB/ogHFGxn8Gx1q7KxVYtJXYk3Wa0371xnKy
JZlgfUmR60qJ3v4GAh/C76Ho5VqoRG/v0jk1f2sr44yiJX9AEmGIjTz0/wSTJue9
S5qhwNyJQoDPVgIcJj2aip+UdJWhj0SwETUaJAoKsBdwdyMhpsy6RdnGcHx8mW6E
wYId/X0g+5ejjrsxTm896lLIJHRjeI8LxpFLvEeXqtAUyb6nE2oNhMwlQjcE/Qra
kspHNkzo37IBCUclaA9S6GFqlIpwmsz9jcKlA2dmXM7wvkdu++q+PXKc0AshaUpo
/Z8cScOZ6ITP2h9wIwBTwcIY+sDEtw00TpEe5iGdhMllJrphGe7Yh2V55tnqPAKI
X6/eUPdI2zbC8mbLviKmo2GafxT4Vw3o1YTA7ameBvwqlc3EjsQo0nfMNVWyhHqu
iCBjJSNSqd8BQ0pn5Bk+XHws1GNxwKej+d5+lAkx2cjC7nyLsD+HYsKylWWxp7Cz
e/H+pxAfg/qIAWWTnvOuTDET0Ezg0O8oc5orFRnRiFU2izlAr8C6zbxx1BxPfkO9
96iaecnXYcd3uaNVhdReO3G6W5I3wKaj5BZQTWY5TXMiMWdQg+pwCKBYINcFJHzT
EudxhkYYJxS3A5LEEro/QgKdK3PgMBMrAeQ8EsN4F5zl8RAG7aFtNstzSm/ya+p6
gwwZFS25Dsx3YHjqEUqPziVcm9Rd3WpMhCFUmOc9sm/QHlPRJnb8LdnLM3NoDBnL
z3DzwaejBq8+SXAx5LAyxuJ5jNHk/PIAVlSvBQXU7PyW3md4tt/x2FnqNrmLwB3C
KpvPxkMuUYeqOzcD+9i+wB6NvH8RAg+ABfO5dRqTNbODr+c/IwDu+LHZKMCtXi29
xsKpmQtmbpiS9wiU6AC1iEaocVkW3pMlixsFxkERqIAUqpDhDE/k2btKCX2Vpakl
goXiCTeU0bcuFwrAx+gchyefeQcG6ITsDSQUJb9EuQ4c4aSX/tFb7vnHMuqIDJrA
x+RPrFXWPbC0Xesz+q9CMQIb6+GyLayu1OhJWpbdgrcjVvdLX5wgQYZVBmBRszWJ
zbLqi5dYEZW8rvm7JmF1D9Gz4n9OvLzq2ptk5do4OvKemKeNzp5QCpVNMXn4tGEA
nCG1C8k6IPYD1l7eg6zEIRuDh7Y0R8gIvzRfSLN3NdUCEh2PvobsJU585Efv/zvY
Hi5+/V2mxdeENQSy1bUEBZFHbEuA0n7YqxHhVbzmbWxmFEbqCDwVWooaeqWlTvbi
O2+ZueFKHqJuNs3+2u9OHu93PcryF7JbhCx+6wtdB0QYLvrNKkEb1j1aCKAp85wp
SoC2uAQtpTcEuoLOTN1qupxalWOvLCz+zNQ/6q6I5EieRlwMFGOgD+5Hkx4AmZdc
vhtiYHXbL7/j9LlIB5FC/RoibtGS733IGnWd9VnTU0cJJ4aLPNNUZiPe0Bw7wkEM
Iy/Xj/7TiYnRBtQoSJcKOKbdcoRlMDCHjCk6iytheedBvP2PZb20w1D4ftQhEUF4
+TCV6oZUPlOgVA5QULpUCGKjWm3bmGNcw7BAeT8lzHHxGg7rrc/UY/F8q+j190Yx
IumEeY6ZuiFM3LtXyi7s8Le+XqhHoP/51je6u9EqwqlyJ1LPIr/SxAykd02PknfM
r2Tzy6YTi23dsUcSj0Oeu1FkVt2idPRh1MjGms4azzQ4Erm+EGdh1yKS1AIn4sqy
Ux0p428P2QyljzpG9A51XKQOO3KdXKwadfNiNSnn3QZ/DyROFA60MlyrNEhUSkDT
y9Ii2J7OhPOaS40PntBdsstlqxbNy6Re9ZvlpgT0zOK5gBA85wh2Fz6/ZzOCsg/A
f+w3F0HICUahvtXwYYFciKEYDeE+WVRhInoc6C6OX0uQWljJOWydJ6DdjY2ad1IQ
hKp+wOdvpwytqHsrYEu0yC72VzcnA7OZG2KDaF4D79b//oOFTV7IykIUBnFKpkf0
WCAG/HrnS8aWmmUnPtwj6pmc3j1N+TP79ZgziEfcg+onQaqxLa3TpVqnqPOR8/Rn
2NhvQ+6pNBC/e/9AyKyoLcNhWPYyITaCjeF2+x8qAwvO0YR0EPqOVDJa9hTQwnHF
odYUUDZJDj+Rgdy3PAeZkzl1NuBBJ2eDACTmA3h4yUvmgYyWVyKcJeNqJcAHGD2k
CxDnu4kM+NFOrP2xaCc3V8+o+7HrOMqDHIwtVX2pKDDwgz/mUuuLrR/8kgWgYPOG
lNES7p46jsMwgL0OrFoOxdM4BYTok3rqsGL3AwogDfVloXOqqPhlpobaxq/I4JhF
71lIy7/09R+WVRf+UGAML5neA3w0zE7MNMsSvo7VvnjFBTK/SZNVw/l1c8NWV3qX
pX9NG/dQekkWDQJdRQdaeN3ch7VHOdkc8yzCUmSUJjtTxjRaGUluPp/vMufMv//3
AGyhz6Lu1BVmZbyYdKjEvEjPDUzyWlTLo3O1bZ/kP1IfGV0bmfBx6hIaiXu1zhxg
l8HF4iBaFJOe7pN18xQb4SUIFE59aknH0E6ZqA/Z7sp4yM0BoR1/ybPZdcMfVPZf
hqYf16YWlN+9BM6fP8sJpibuNgE6rHB60LhiHEthMHmOa0jIn9IEwpyRqn3X3kZx
nEIfBKGSEZGmj4mClo6X8AhwcwsghtysnYI8iGZt/u8SktaDmR+inc4sYq0Sn0Hb
ztozWkSov6qMwf5DP4OBiOVP6C/pDu7eTzyc/Tux5v0cQljAjUSjHuX3jBn93lTe
oNoJsCK3QRMs+XJI1CKkH6xtIcRQ6qLGA3MlME2VWFvaeiu0FXB9QwXN4VVPI9/k
j3iTiEW00SUNNHSgCOXNKOFP192IVqfE7yOyf/HcWa9V47DWhBpEVzN0NOxMjAgu
76JdCLuJrWKHqRdOLh4C/phx3LW3b4Co8hgcJyy3haZPcQQeDPXmajFv7RJcbhQb
p3VFMxk5X1y8yzavK4juIzx+j8hxZ2vu42+sVHdsk2Cjml/VsBt5yB4behZZlXX3
VFKRJTkgb4kzm1l1j76IshtvMFqnm0i6rvxZ/PLiLQiTppnjrJVk87043FmnOB7I
FqCyFmwYfBkRWNYof2hKjdl0AZvvpv4usmBfX/7otLFBIYa1M7hdA9AFg1hLXZUe
HGAAJFWvrQu/spPXGOmuE2W0KPDCs3i0+at4TrbnpDU40egdvLoZBS2xVWCL2C/n
0qHBvhuZZlCmeN9eg1hDr4MBk/ZRoepG5EKr/Uy8OeJE71EOELYzYDeg4bMpQgF2
uJx9Ln+xmaA1dQdFs5lJFgQ26zaB2pkNj2Ad//dESpE0VwnBO613r2ScWO9acppf
H4WtqN5z5w2YeGCEXcAUsULWaTWDeLXDRoq2pR2rUFJpd6Xb0BE+FE0dUDlqhEnR
TzXk9OVR8W5A3Xb+BpwLRN/eIi6aq0iKN/FDdtY2MrtonHTZondzTEj3KGSAtDrE
udLYxNgUQWxx9OxieAEBIXEKP7LonGL28swHskHULNrh+4LgPbS0KDdzvbRebbWV
LcQTsqLgUY8Um7GTmiA9o/CeZ5VzcmifN8+TZaU8qMT8LI2OO7aQJ4XEJwKB40HV
pQddpEuGUv+nqIjoNunGY+FdaxxuYRs1msGinfcDWlNRMJekSaT9iZsjaqJGpVZo
Y2SK9PA7ltVVNil4dhTjQO405oRO7c3xwL4cq93rXBrXlg4ns8kNVkffvBqAUhr3
lnf9VcjsxZtt/AjvpduS320vgVHr1WJ9PLkkFfyPEmv+13PH+AZtFKuki+DLlDC4
C430hTmcF1164UAtL9tNLCs1eCCovpEFUj6Z7FJq2t12WKjQQyz6AhGYKXR0Qsx/
awSl+my3MClxJWx2yq2nibvNMTDCzpcI9DXTHrzdoXKJ/0H1MCXtgIst8H/mJVa6
hP2wkruhlDnx5CbFhLCCGRAv2IZ+TmesZZJRZKve6MQqmSN6HCs3I2SfjuXAArXm
agsS0lh0uJ77flVNAm0GMI5lHnHf+Os7gVrZg1wjLoBUOVVaKLGOJW+4qKRcDo3X
W0Spw4ltYFnBrKYpElYNeIve1kt+cxPxrFia+bqXSPEGTegxyTygSuUzDAKSqkDP
MmbI/LmRRfic3LUnAJ7+2PRmhuTMMoI/JH+t7Ui8RZQOEvsVuz/2gw1IKyp8/ZLl
qBvPPzlVMhSTTkJz2LkdUTGitgvbxR0SyNm4SBXJHH9CQp+IhhMch02k53Kcv8pN
GP/3KF21/d4oXAkwrAGCcbJijJm6x15FEIqbbSzj6uyun1fG0GLWM60WYUgQqN32
YMiOS0Be7XA1dKMNEqdkUpvrAYZmk9psJc/hGUyeoKA2q+G4md6lKkg00di+IK7w
WNkWMS9MGi2IPbWAb9ktCf6Z0YfZYYIxrbA1V+fUUcGnh8JSxrQmwkftVZNqE4/Y
qFDSCZvSOvNy39eKKF/n8DMKfuV1vSd/GOP23/PKVAU2syCxbWHbPMgt0XAg3f4A
84PFEMIklVPOvrk5OgE7YrEHgXpe4d6zfqmb5MOX/J+IGmfguZ1s5BjAImT/1qkE
dmxB6z3pUipDsSQnkn8WXiYpR+Gx2ndAtOrhpqkQeCPOiKxRsXOBvtOGeDH3pdZj
XayF8xcAQbEfFPbznpmkkjCf5ge3FGX2/RbVyNMX8rq1qJhjjDbBwzqaHEbDZx3v
1Weq9LQgqGQ0lR+1afZ3Q8UujUO+icf2Ew4lzRla/A0Ffx5C0X2l1cID7YlYlzWC
Gqcc0qof7scIYCn6jVDxvJG2KDSqgxlZn/EH1owr12zNfJLl7ydtK7WnmLrN+14L
BVHSq8eaOyppSqpOZO+3aWkJlqerh+NatVGET8clxlymrVqA52w7A/kC26sZgymx
wnwIDbB9PE3JPTrWlXun4Nf3f2C4qqz22Sumtjk4VAb8NvA3jmbt0ZpqKuXdDQ3D
dicLS4qYfc8HL7GSDgthTduePO52/hhq6/Wx5Q22ACviGm6ccAYxlJmcWWhmRQ42
kCwxY/3aBNYmE38gDVf4FOiZcOmYO5aBblsknhhTlEYzyoz4RBybo/WLh/xTvOz8
9C+HPVR7xglbz5HhCwmAXXVUJ1zZ3yaOxG1raHjTZZBvan4r0YnVKOvjTMtz1iB6
Cdn6hQmqAL3hMxDyYk8B+ulooMrax/6LeVqzkIV/t4Pl/mDbiajiahOeCOoeohNb
N8mlP9HLG4Hkj+q6muw1kohs4X3Ip/9YD3ZKc9M3kdQeAqWyOLADe4kAKL05yDn4
qn+J6tQEulYKbJfbvqzsarTeiaVVx9i3K8hHWI4CEFO7EGR3jweBoAi5ZIONrsIq
m2qY9TDWhVnHlC1d0GtT7Of5myl+/ozAR1HvTX18gs65axDJ+StvtfiW8rkBBi70
wngiWPQ4ccHayRLh5AwaC2TWTd4DmF3+Oy5S5RCKFhKY3u/ZoCBEOgAa1FKEeliB
MoHJnQWdyROM2p5arhjIfXe78AEuZd5DHXINyzS8k/2OyxEOl4q41YPjR6giHWUB
qWu4yjO41C3vxmoXVWDCEHVzaNUQ/6Lw3B584F1m+njLBri+Sv/PYC+W2NV0Dcp4
IBny8QNm7dO+lKabwb819imSZOasISfW1dsPh9lToXXWNfHQ0ZxNarHkdsE18hF8
sJJTx6zF7DA1DWwGX4Li21/lEV+G2CYgJeG8Kzf5OYpgUuirLX0U+QxUahY8Zi2B
edoPjxYf5GRj8+N6Ni2yEGvwTKFwJd7rHMwfCAKlcgDl95293UQGzECgGOvNaSsg
K80Io+f3UEsG9aJvJ28bTJZhnY8mfey9k9Gd50okkREr70cXqIfVRmkD/xZv29+Z
wtLDUAf2kSvaB8uvqby4yr3lUESmmUFrssJ1r3sZxsnAWxalTBA8N8XAZTws/8TG
DBvyCJCj4fn6H38RVzUxVz6GjybWprpthRcZZMQejeU07iMg46ML4MQXfxLPDJog
i1MZ5l6AbZv51TgimFVQRqac9eRmxB7J3sMgYYIOXGEfr7nNSZ3BxdLCL/7Vbqeq
ckPHlNiyLF9zFB7hJyMqupATd+ejMvinTotNdnGAg6d+WWT5R8Ua5t3NhWRczN2I
hZ85rQfRiBp8EPn1qUEFfwEPva8EF/LAbJG2iCzM2WDEXFBfDuIIBhE6qrppmZCA
xU+VjxWppqJsE6r4ZibDEKrJjZXwH7ZycdFnFlwK0/IlEL9Cag/3xnH8OMZ6j42M
h+22BPIhSMt/BiMvCP9sS1hdamXMDXXgbd4E6lETkGu7PcC1MMj4TLlEr5PPhPvI
5atTyReGBI6QKnxZIB1srY4K63yKNc2u5ATRLkKOX5C7dJABlcaJawrMGESKYbwg
1Nq6C1INKubUPXNS2koUU6MoAeqGchGP+BGlKSTO3SIvhbF4znxGOYQT/QNWN+jG
2y4FQ+/VWSQsnJJVYJLQFix0/5FGdbb2h9e7aodt00v5PCzMQMtBDo+4eIaSwCeS
OamgzKxVrVtSETQhmw1DyG4MnMo1c99wpHUQy6oUEnOjW3gKCgExjaob0ba0CQt5
7gDl7AHav8tqwgUk1rwUGCC7GaMiz4qxI1UAzVwULJQwpNN7bq7zCmjBPRbFZNwZ
W+VRdb/eyI8A0OqOri9ZMkat2iC2+sLBrfp/bNaRI5AIuox20k1pOYfpM/aRQo/l
efvPtsZCmPjSB8+ILmfoRzKrIR/agmTLTDvqqqcCbNm0LmFZozZbB0Bbyx0KH7QI
+1Jig1U7foUegsWl4odCNqUteHVGQrVyHZBdFB1bFkwtgI9/NOFp8SpzM3XlZA/N
mvc8w69MKBYddvI5phMnPUAlgR5+zg+FxUtBOurMmR9fBjhdqbD+W8C59Xxt6Y8Y
R9/P5pj/xoldt09KpJy0j6sDHmQ5XCx59SlZ/f9imNodphScN4IH5JTrbo6SJ7n7
RRLA6GMLSTTmsGaFRoC56wHCPZyNaUuGlOgbOI4xTtnzDbTdJGTQaspB75cEnMaR
eFEDGJt0QTVCcDHkOjUdJocHK2JCqWmZbE+asAgvLZu11r6xj2F+VCO6tk9pIYvD
Pf8KKFIkKu+uwFl9uIgeryjUTqiN1CU9zLczOhM6HlS3pL8LhvpoIa741nLgZjS9
75LLZ8c1Zf8F4han73VFIzScS/oc2LVpx3/PMY+0IsS0KxIzPl4TtH/k4ITj0PiX
bZz3m/xh1DqxFUB6y37Dwj+cBm1ktWEX6NnmRK7jh1EQwaRbuNVPI5lx51FlwnG4
6k5296Wck5zjJsg2a251zGSfos7oEsxN43DAUP1HnA8JzRsCwgzf4qLtyxdKZDQb
R2gz8yJfY257NrB6M+oAmq+yKVygBjhKsAqyHP9H8lppEZT+69i7uYTFgO1yUOJ9
XidMIHWHi0TYNMD7GD17UB0vIEmwZJg3coClIqQGyIOYINuvNm3cHn4W2Sm9mPlE
KhxsMolyX0R3wLtyYKnkbCOVRrXKfiMzwS49pKCy8gVoHNXs+u8YA5HzDrD0o/3+
lV+LgdC4vushFq4dILQTQ4zx6qOSBDnitzRs2gi0AyZEcELTRYFNYd5ax0Hwxutb
IltictvnxUPshYYyPN1Uu1UIywvgTlcx+Isu68oNCSzRORXG/EbKgDDxVTrA4O/M
gbNl4JMNCM930QJZy1lpMWiVrjaiiF4sGd1QQz6HFl+OCSc8Sx9gTJFZW+DtWFnw
imurCCErY9FXRIjJwLXh0qq6uApw5mkYIPurjBiAhoH7K5HTbbLB5dQ4E+W0ebmZ
W5hgudTIg5oFRuDufhS5WEoyyS2oPu8OSgudSyuPbaNfi0r1FbZv+NI+PiXXTnex
8WWZUh7dUxWAXcgX+kUFZVOEP7PIIdxV3zHAFdHVqX4MSpbdqQq+RzrSVgbYiSBk
TP126MtCPlNlYK7GND/8uz2IUWslGU4KiTvP/njUokphXJo/80w2hTwwCOrbeh+C
HZLctadXekiCJdFSBYvYuYFze+M8HO7S84cgNe5ynC+TgGWYjLZJy7781si+RdhA
nzTdtYz6JoZNiSpuTovxqcFtsuxxtyWIzjChuTJXuWPuTJh0aX4f2QCsgVrhoZfF
M3z98EaFcVZ6B2rX0M8JanhMC4hjKR3hrzuN85wigsBId7FcRIiMqwNYw9TIJfB2
KNL+2oIszW65+ahOR1EY56nMcejWSmo6VW8ZXChFJZKe1uVZviY58iP49gb2Ox9m
RtQUaWBmLdgDz0YKJuqxu3mI4gt6WpwmwZfKQG12+wbRXYsAUL8VL8yjrR5g2/XV
U+g4Ib3UoNQzqaVLdMht69q/cOKg9AAj/1Pyhh8aDK1TxDJN3CmB6wDov1IxJELD
xxjvFVZoIsfIkFlt1BKaQX3RXw/d4YkpKKA3nYc4AG17dZhB/1YeUbJ+VbMNd1b5
jH6uFBhYLhjAWPrjGIN93KZ1PLVg2lAz0Qa0ETVVUPuG0uyoEKfhEn+jRtBh+ZBG
eJrrTTaBxOW6oYZUPSxYc+CQ+9JdsLW7iC74oq6ulae1L6BBuaPr3bqFMh7aKVF8
l6HpLTZCYZYtLpMI8AdwKcc45by6qRDV/PukwG1H9IlBETCNbSm3z5t8sBt0HFe8
UNw6Hx2HZDsnm8PcZ6DQXQrpklAVzhD1sa0ZNSnxElyRIa1MrDgVMRS6xKNwSzjO
SDE8M022hl2ynounzvZ9lbf5NL/+dndCn7vi0deJEGyipNHVrzrVcjgcaEcVvYOH
CithkYdAZI5qQMfAfXA6wm0g6AkHeFRrn7EHXwYs0epycqgRYuUQYLFx8g0PUjGB
e+VajcjNXZCOW7Qr4+t03HbVZITrd2VuFedtUMAnVgR05AQ7u2PgHvjsTO4YDCTR
FNr3SZo/Zn2B8tvZqIx0wE4EyUsW70eH9t76hw6tNQZkpF5F1k79h72K7szVoexN
lTha/IhIyQVIvwobzxMoQCtDPZv92Hn7t+8FtTOLFptvlkmKF2UCsAK/5a128pmw
QgUvDIlu5Lm8EjcPKD6A3i3W7+ixGUv77wknx5iBmR4hFL7GyYQrAv85BR3Eltf2
hiedlfUQuL+VrjBllhCSsNmoy4ho6G9v1LwHYGmFa+9OqVuG4swIRl3LQpa/071J
lF50OKLesWjn1DSsnDb3hZHkUlvXnCwg1iqqpkgCsdYx9Sb7i8yCx0WfbefJ21Tu
Yorh5R4l87qhNJxXllkIapPOeIIsEvRLAKrJYa0Ip/77chWUwXwouugE2vHNp8uC
k3oW466hCZ3mJ0qkQfqhMR9jvgWUykzJaRNriczw0C6dKPKxsGldSxR7KDP6dFGO
jBJGIpZWsZs+DMpw46En1EJr+pZ5G5qGYtMqrbLZcBHUn0tXmOgK0h0CCrrQbPZT
Yty6VthKoAQwdipiP87tFLm/rjbNFTP4KuavL+P7Vt2XPxpj7VVbMw63JkwFLsRg
djzb/UgeDFyeDtVSqEoP1+O2YdTgRj2lSNqLSP7+x0qJeP+qIPQ2K37vpHEMNTE/
/s7EYjVCgmzhqG675X+sEsnmx4ZJOn2jYEWQeND6TVGW8kT9DDoadq4n/zhLILJM
z2wd2mQqzg8WVdeP0L40jDK7UsAtLYhzvbeibhweHI/KAOrgLiF0LzGpdByuV+GE
9vvuw7dVwzl2zX/fe0we+U2bNDFowb2/iTU3aOFeulHpSwogJLrXRkw+XJ5WakNL
7pxm8HehHCDjnvJUpwWRJO3ArlQhpK9rVLNK6XVFKFjuyfSC3Ij9dCXI2dDD32MR
wCaZpyLlLsTcQpErD4brK6vLgHVYvKy74in4/WmBx5bV6kJuKMPkBYQZ8EX58Ggy
hWYL2cIqRRDZPaPqqGf84Hc50VOiDuEqGGQmB0WE5aKUQAkwZO7egKWucr1qRYZx
3Rs3N4FSzCtbDJKRIWzoLOez2MpxPWLJnFS3F2h1Hl6MeWZ9VFkJVI2tBxaAe2JJ
BzVnOODB3mCMZ+duxZuThhpUHfhg9TOCaUHKpamf6OOxjLXed7kLunFaLEUCT46Q
KQ7qL9wXVO5HOUPrY1u19DlbUPJKduJZE4Y/SucfQ15xVtOBs/BEa2InuTQcrOwu
4YPgvqbhvE9kBRgnLzpcZxHCwOKWsXQU4G5CmKwG4zuoZ9jlLrKsQ6JqqIZoxWmN
Wke0Wra+PnreezRdyPOHgbnaD9D3EhLdVNanDzgIbJa6b/B8C7wvsj6dFNSEXKtM
3KptmVYxfnnBjmn4ooP21Dj4scQuQ843AZysU4YKsaDvMjzda+yA7PpJEv6MGrA1
1bb2Lj5ylUJOTalxActAszTn/TZgrSzkcUuv8/2gi7Yq53oWAszn2kDDogGQo7RF
QKNY/L9FMXbwC1cG8wKvfcoPwcP+aRsTYM7CCl6u+wlpSONNU25el8dPTVuUTJRX
QDK7wxZfHhwVVMgJ8eSV8UrHXYU1xgpnGNvVlg118/idKV1Pfb0jyKub1J778NvA
UXq1KaMSGKExIuYPz6lKFoth0BggaP9nkH2cD6OIwH+1XO0ugew0MZRvoZEjRNcx
bpkaZYIhFUnX5LELAx/6jTpAOPxWOIOkwak5G/5wXi8n38/VTMHnUjsH7abkqNPK
BJZFgQapJRlu7v1azWglFahvDLaiXCNMIz6xMcav55JDzMBku9Sb/1k537D5v11z
0N/P+rnHR1GO/Gj+lvy5qNJEh0qMA7Q/4BZbaKv2jmktG0vo7hITMhmDB2x+jKBF
qY6icTaOr9jqQdd5EVacO7UGrpxGSK7Zi3JaHD/qBofVG3dZLbM5sV0DOfpICTgh
5DFb9LVYlQPY6IfJNDO3O6Hw0U9e49OFnmktjCIKo9+91VpvPysFrLXo+LgIfoHE
+m30O65kRHTWz5CsdO9CAZ1xsfyVTxLGDtpa5CQwrKlZNEFgdoHnej/Lb5+YgHLJ
Uud9OV5S6V3GeOgZEItL441dKQbxZ0/o+TH+JGcypnlwOBbXsNda9vLIJ94Pi7Gw
peY2F+ueqCW79gV5FyGSur//Y+ld/1e0C+gBPslmd1d5WtKgEiJ0zHrHY3jT4gss
sGAPvp1F/bMlsPITjeSC/obPhLgX0SyMFssx3kMVDMScBBbZhAgayObHzJUpo0/D
tGQqCJq5E2QuoD48nSoRzIVGd3XeSpTVDz3KzU+hLXCnKSxWRFHZ2ck9R/oqIDo/
xfQmAxt9CT46oid7pEsBtpHsJtp0IA8kZNVph2iy3rGg/G2xZr82LwSTcBwGW300
SMI2fpB9rdXwsbk2Kl+M1efPnvk39h3ANhOH78kCENRsEoilA64yd3xRlkL6UKjQ
Do8Mbw0/Kj8kbb9T9bOa9KgVYy3zj0EqoTM9j0l5Jr1GHGH64ftrrFKHt0XsHtdv
G5T3rJ0nm+kjN4eVVvZ39VD1TU33jcyu9bHGhdokKzPGGja22wl8wlCY05PTR0Eu
qkL4fYCy+7791hNOH1EeEv6tMLNS/pnIAowWM4sQdHMqbj3aWNf4iYePqHkmZbco
res44bubhYy2JeWW93TkwQOg6M95aK7aPCaO0MG2iXPJu9ZhQG4Okgb0XF/xW4ts
fBT4qZZ1eDAnrVW5a2G9/V+G93dsPhF/wgI9XOCCoZ20jXgsMEemhFst9H2fL6NL
4KJBm1GQFLQ03yn+b57L3swKzUe189fUgeNylwasgbM1myNI/1qiohM53Fg9HM9t
36foOyKCHjIc//0QH4n/2WcATgz+DjP0J9XKbUGgiIYg2WFQeaZemVQIYS1OfbDq
LNmQHP04uWLm/6GI6N955PrJiQOSS4TeUFcN7hs0HMS93/Xtt6GfmJ/jkei3uk9P
hbQ2LU78q2lbE+6IXbQQSUBSLgvfM7rTfKQHPLWC0LGu6ehK+/GvwBkI1Ni501ly
ay9BdKvDnzPTCbZC/bMtDedjvvDGFY7e5k51tO8D4j2bjSPdxELEYCATBdQf8HdX
ZZN5rEVLA4jAC6sD++XWapg22+bg5HOohQ3+5TwQI5n5nX0izyoINqcWqzGpjcBu
IF3/bJL/AJ2QNVt5BXXrBgjZrv+TvEKClJsBlNobDLu7nv6KzEDNVFZCAvRDu3VQ
dWmbnUQZk/YrOIwFJp0h03jXiym1ek8DNau391vxOEcI83RubHfwiC0asYkKhepM
EBQPgKIN1qVG8cbka87DoJjRWscKQjcV0SBHIu15NZfoxN5Hy4PDKiZzcxQ4E182
KOMngXCXh4e0yNzyFLHM70XGGTOAfUPPFb7pvLDvr2WkSajfFHWRIPBvM68N3+dT
+83+9gpcig1pNll75XjGpOknHULlMeaDPNv+HtX3g7G05ksd+LSxSvgNlU/cxESG
hx/d1KNoROpRebSiQTRmnuFQpUuMU3avV2tyzsRAEAaUZcrZs3UIsfBl4OjUNqSC
bnQEHOmQubOEJ10T77tlA21NqXNs/cnEughjyQ+U1CMGm737Pg5q3yoM+GbS4A3l
v3D9KrLdOWLV3x1tdCaBQPzpHiqhhFFJZ/kVoyQP89QJ7q2WHvHdkbvOKhEn2uqP
A6HbqRIwfADg5l+XBxvXbNp4TQNlavaqSgqSuWbebVIu1YW05FHF9fXUEOarZ3PR
MfOAuunT/yW9OZDef7G0ha+waM1s5LxGbDCLR4PGVbUswo5OpICV2nEkEvkH8pIA
tASfw+0sGUwEwkFQMlRn0pChNqwd3WO/OZg1hFOMXjEKzjTD/PXMEASNDuLBKKy4
O4+Xi3AdXVUWaQJR0W+P0QsDRZrEb3sciy8VF2PCquk/qKgPSGNltoKd1UOeQhMD
ewJd7eQLR/DqnoCV0Yoc+/KdTfMTduhrOs+MaVzQKDF/dCYE6n9MWyK4D/i8eQdI
mPDsw+2kLStBH+RMjbgn0gwirtNQYEo919sLzA0t/gHw/jOf/pbdQeLwhgLvVUFP
1TXSPIPVnuFJi2RJ2MzkWg+pX9H7GF9MRnx3a+/Z8QZMUoDskZbGFpB39S3AgR4g
5mFc4NlIZwvsVDjHddWwmAU5a/80DwLcl8+kLbW4a87KKe4XPD0aDC47pdps/QRc
ThVs1Dz8Eg0sZate6N8+bA+hzgk0rwL1Gw01pBlxmQxNzZCDNkgXISky8FZGcCmB
u16CSgaPIVsXxMho+BcsvA6ptSgBuXWHq90a4H6Ja+O6/MqZJQnjQwWuZ+pXLKwK
MTHTeN9sLidEDREJ4nepnceV/DUVcga1Ifk/ywmAUZuZTjj97LEnas5fzQ7qVyhq
tpFb5ljW9dCF7MrkcEQLFh9FqGMQojUbDXvDD5DEj3cB4Eh0DXoMN77P+83d1O+S
dBH6Fr3Y96IbkxjJfXrtwqidimCz2zBPUQTQQv8Qv3bzCPaUdDLZv2AnrmAd1JcS
S+Oee24kq7ZFx9/bnslAWYtF4YOCFNz6gQGvvAh3HNVb89xHmfE+n8f3HE6Z6BwN
8QigGAigk59OVPLMEpmrxF/huX6KzYsDIJ40DtTy7SgS7bSDBlVOf2S676RCID5P
btgK/Gu0Y0GvwUKa4Q3h9xIBQDNJFZjZzZjTtFiJo9MOuTMMF8gYd9rqczo/ku9J
Gj1hr9P6GVk+py5O16wlCQ2XGA3/Cu9EKOL1/Cn8tmOLC/Vbi9mvFEGRTxNTDQS4
TN5ytBAB19VcusXUNT//ckNEmgb57C2FAHhooZxKFuZ1QUe31sze83+eVegbOKmZ
ChGxxwpyMKzYo1AiVWZUoKSYubXmOWXRaljIB4ZDArB2eKTucwm97PfG7/AwvKxP
8hQ/Niekt9w5F6Bg3zFI4s/wlggrx1JwaeFaEMzhg/pTqkoO8/IBeCyUMqAAG3ds
hSDLsBNjP78QbXNrKqktNd5gKT7YHWpsst9HXs0RdTQYzX8z/l52s/JK+v8iDtsD
CQjiBlcfVAEi4V4w+tGT5GtzK9AX2GNa5Yb4uUj79BHFyd6uqLPyz4Qby1uBilZr
M+YJAzEvOz+2R8X/wfPyWlrazD4ugtb9yXKtHas00oN5e2FO0U2mTxDt5aS+q7hB
x0stT9IunjVrF2zdxPPFNRwSo25PgjRAPWYi69Z2A7HOdzzzuGZit6rm33W4dcu5
FFVV4gvoV575ffpoXN3VuaEf5z/8poB9salUmgYjYosWjFWFbRp1K7pylSX/9gaB
dQa+NJvFJZ7KLGZYe/k3tcJs2yADMIV/UMTN8nrmBMJBusT1bb0OBlxST9diHV9g
sNIWieLA6/3CDd3JVVMkwa35/LzPl034tVBppKVnlosj1JtwUhGFpX9q9G0qAAvf
xcD3y5xd1Kqua5KAAipKOPreDcC4zPDKbZ07slLJ1EPppkSbF9E1FBzMfPhPfyxO
qbRz8ABHcTTK8taxuo8WvOg8tV/UVPCSwRSauehp2QS8+Ami4DFmF6E1imLvhPvo
8211T5YVf2AP+GUZca/wCdzbfj8vegq6EWcI/80D8PEw0SPz+DmkE3q35QrS7sh+
OVh1Gor1VvB9PQ4ZvpvydatoyivI3RM21412NX4m5BxSElvlf6n2P+Jmw9iycs6L
tXa9ayNEMOYyi3b0ojTpjbWkrphcvMqTlcMg9XcmUdsx4LXmqD5uhNaHGBj1AZzF
yX4M2Ve36LVbVM2Uyo8/rk75R2rgOG2t+m/mY4RF7oaKKeTewBSaC+YVL65Pe/PS
qJ7d54tIL0w4A8X7Yim06JShs1bwx4Jm3z/6YfmLit7f7Mev8jCtCyapFrm856d7
lT48X/jiCGfseRi5/oPYPh6jJlPagNIvErOs8azVa/STEG6Tfw1l6RznQNdB7XeC
J/OGehbri3ZEoi52v6tgXF4a7AWQgbxoe6a/Hp4Bvb1X2JmOWaKmHJTMPZ4Pxg7d
UhqGPfcObdafKxnUVKglN+2L/I63hApXt98WinmAlTfZabZ4gxyijRp3J2MY7ppP
LKb+oLXt3RhuV7HiedvLIx3VE5s/1BtNH6Mg89NmXgEMjVTDiDHVAcjhC4zDVlaj
x/TXa7BklMnfr4yr4xnm1twaW0EYk54d1UhQFgPxlyduqdWfKl59q6HIkD+nPrLw
xoB7p/MpVDtiZUL1fDXUNx6behmj4kTt+FfRWSdVQgZSettvHSC8vFSBT1QizQRR
0OsCS1PYanwdYaEQwTxZ3lRTGoQpPLwIOsVCztAliBNvwzOmrTR0yDY9HkGJSJO/
NqnGpv4jhL90dW+ObPkRaiojFRsaQyGedluKaJhiI3DtwpAaRN2+NNn4xWF5hM/X
05kOg3vuVYHdwy68rbYDHMNABo8wkJOv+gMmhZPDa56zbvfGwu62H25f3eHn2wlL
NQkS4JQQeH6qrRRR3mCAIPMVac8UUFmCWo0IUd67UHlE8cUUuX0MHwn7yb7CD8H/
Waztnx3xbAioz7k9h8nt5aQZxFC3l/Mb3Kgnhup5DGnH1NITUcWMMIWAWIeZs5um
3c+91awo6FgUeMeMy/rcLCW2g57dpmq97TQDxVpYcqlECEPw2eNFqv5FhfT6A6+M
2wa5wn84V79IsTVWp/aU7I33WwG/o51NKcF9M4V+EKuWhgXy4ksXDf89IZe8NPVQ
kk99D/cQDqg7PIILeVzbdOct4k4P+K3tHlEUAGou/FJAmZjDXqajvOxdY9Ui6wjR
j250uitsqFRURfbw/gigTucqw+PbvcZactAY9Xdv7sQ0hRic25oclicVcrCr52df
boXl/qmycl//A8NbXvqc9So+X9yclQ0yJeIPM+VKDkh9hZeYDXRw0LuIdm/Zf6CX
b1mNE9csxjlPjEAaNRNwvGat3yCEqZEEqQHxoruE8nOsH7R+/yqIhX0lM9T0gz7H
/bZQVQHHkAJ9T1pduxJVJwcevE0MIoh+UwLM/OkCVEGHT7b7jO7T5DY0UFZ2CDYj
JCv/157NnZRL6KsBliqmirG9l+a+90uGgS9q2ZHQEJnZbz1x2qQFcqvW2ZXeyZB7
i5UMYw670B1T2k0/dpq3CTKL8UKh4ULBSubIpLwz3DS4tls5uHBacs/+88qMbmIe
/Xt5DLWNtXXIZlJjB6VXNXxvC84NqQCVG7JeKZ+ydQYngVVo38S+w5arWmRpj5Fm
ux4Z5g6SMSGgft4YYwoaKKhu5DMsTeDEUk1Hdw7pTbqUb+pnd2tb/hfO9xuP0zJd
KNHdSw5qvsEgx8GI1OAmUcmEQFEnlE8IDcYewXFE8fXQEJPA2wdnaAyZu7dL22i1
shjGQ2ZNrLXFnefNmw7ybJpjJWkVf1vwHaOY+p86u/Xaj7LJNvbBsi6qSLHxjg/f
jLBT0n/8bLODf697Samsnxt65gpsa/VmtWK6ON+rnGRUtAd1VLF1LW0bG2ho0FjX
hTVvYgprXNQvkZ995CErgvXCcCumPFDGkaD2cNifQACoHWMmDyHt3XefRL6l7lJf
wePjipEQTRlhJ339tRzoLu4QHJI7dMnx/4LUuMy+WJNQrkcu6BwbrDjq5L/0SFxJ
RoZ+YPs9G7YXJrtEd6RnG0YQ+xwxBeMtXDhEB11Dp7trvnApY5XshTluq7W1aY1z
9qEty0vX8q9l4ervU57J7Bj96E1UawQw4CgAkvhNMPnEgCbQtygKgWs++QoZt5yA
jgfHFWSwGiI/OwzihjRFM9UKUxCz+MIa2K8j78IS5YPCtfQVMbo9JCIeZKnSXfVH
5SZpcZguTrGS0y4mXcjpduWTUpvsL9auvkGtn3jrRHHrGPdj6Xq7XPyAAqGOrSt1
EnjbQWqK+i+jzr6gJyp2fQdTJOq5xXOFlI+t0u4h8duxFj0yBN/fnVJJd20YzHuE
Tzh435hcMvSKPC8uhazvqlWYdBU8gJyF1sqcXcaauBHP1TFoF54Cu7tiWujWtjw+
E7NwAYEJuvLpQTbavwOHAldzwZ5m23gS+0ilouB1qMMkwWqpHo6lx4ElCTbPp+CF
eK4f2J/+Ba/HynkNJHx9IyEHMgC5uoFNf91UlKDBjLOcBd9Eg6rfLuceHMt5zwXc
2YTQ+VDth81WSWk9QY8QWWFYnAuOM0PeoAkwZ1kJHJvpiKOihs2EEtvxu4pP7hNr
mu9RecgPLZuoO6RpBIth1lAfi8tZA3LDvaCiXmFDQ4gcQ2WNSiZPHCN59jPpS2hQ
ln/vwmFz9UKT1B0xDoyRnui5MZUCl/x6RF+9OKpfSPEgRcABKG8/4J2CWHtHILf8
nUMkcuLVhs+5Rq//mTvoIxYR/KcbN8H31gJPsrl0ogMCs0+r+3nZzPBnuYbTtbJF
v0K/lyGWDKAWe6ikTNS9PZC2cKu4/q3mrlkzHQ+8CiRiWnFLHlcURHkNDZP+OP8m
JAGEj7CqCSGC65LSyvm2OqEtpikCFu45AM24e8f0f0ftXLM29tk+GivrYsGTEThV
GflxSL8s3sy7qSP53DnAzaNyrdjYdSJT1Ndt+bXm6FDW14D/c3ZfaDdmCyWWPhRd
ig5s5NUg2KambjpyhwCOQmcP32g+76/UNngY2N99bD/eRydkG3cINv12XGJs4RB8
5waMdPD5Hi/ddDoZKpxmWoRLGz2VbJjBCOWxaGw0ENTY3IMTOeWDryCHkMjlR4G3
Y0yUXdhdrX2AingyKkMKlfOMO2+3TQcW5/idHBFUHO0dI/TqOnzdcdiCiUjST33E
wy7JkPrJQKmwBQcMdjQEFE7xm03bsogZwZJJ4oJnr2URXyVv0292aC/smzADdpjH
1kltucK98XZuJXPuFPVTvjBih+zaxI5N/MiKQNUn3/iDYK9xggaeUaHopCv6JN21
h0kxbPrbuD/tRKtyV+HvQwqgXkMTIwRUNiNgrQZL/Vi3ylJ5M5ll9Gua/U6ViaEt
nbhFryd8bg8J9iYpzmLcEngT/Hu7HlktvGmzh/U8rxaZdnUP/iltzBC4I9MOjR38
T0o00N3LPf2pg7/BVkW826VCD8n6uT352MztX1hTcNJ9GNprHhqdSMog7KH9QnwU
N8f7ys9f+FqADTw0/08ID7VdlhnEjMdVkXHWXX8C9mcGfsq5HFGJ3TqaIfjDwMe6
LmpEM/KRWnq4BykNNj8uLMAaRd/8ZQu+Lvd6MSX94uENnUEV2EVRhKQkY5nScbMG
z9MGJ5voa/3blFcvHtDXiemk2eitqRKbk2iNySGTfjvjW65xHUuoxUXEn2uMSNs/
mCRIFPC2eEITIqJF8M87FTrpWqr6FxkMQz02hBzHTsNkLCZPtfHvBsnjpF9LRoj8
VIAVQRx4OFBJ33yxkC+H19egnAmvWd40z3WWiXVUrQV2YkZXLPvk+pC0vp+hqlY1
up8QjkkAOn78gGnIoE2M5XCL7GwOqSTQE9QWXSUTNPDNsXayOEUkIm4L67Y2iZam
6rcS2B6xP/JqxpaPN751xGhIk5vj/mLku9Btst0dzBvNMP5m5fN/B6n7R548Y2gF
PaPh7PJccoiMa31onjhUBudk2RiJ/Jrxe/gWwMIV6efQjEJT9S33APM5hF1emiEF
x7m0NkFri3wYVNF0yIQcbfk8hyxqQNd9yGg5CUTJTdvuXOuwb4RED/mC0CrCatDH
v4q4suS/hk5pZjkZ37V/wSP0LXIQolxF2tdC/U5E1TOJCUv79dQF2GdRCY0/QyYY
hEQ68ykUyePhMkeA1ZbAc0+0z3QAJZ+Y24F5EMq92dkXFzdSd8yjj2et2ZqQl7bG
iywLWabBjnkMGL7AKPw6LnnPxEM4Bsa/7tUx1oi6uPOjXe8Lpb8TYVqCIcSHOETN
GHwPSrndW5Ld0/jjGHW0wCsWHMBeN3m+XJ3GVWSUZuqIwI3pmYajhpXPdUI6za2g
+yovLXFSfZkQeo9PaZjIYTz/GsL1/Hd9LPFSdFFvcBymIHpG93AuqCW3Oy4EAF5w
ZtOQmbS/llsPHH/eNYKHqc+6QzlWsAy3okl8/yc82cYO/r89/v8CE7fD6dpMErRr
1nn8asCnFsk2ouSloddpM0IBi0vxI4MALeA+qRN9O6IZ8M7LVMYwDdgUVD2faRuH
o6X1bVSoz1Jtyac9AYAcR8rQxJuOvy20UeKrkUo9w3H6EFf2UjHtlm0ysExgVzUN
3Vh9DgnbJSJXBaEtzGPZCr1IjO/xAdl7ceiOnpJwhK6MrxfH41vrMaUwJbNcBgve
x3FOdjen4ydBLOmvrMyG8Rk0jRV1OSFl3wgRoQbjF4NXwyzH6ZB/6fWSfbhwAGql
vyy+lcXI5C/73D5ZRjSbqkkmefeNffPEot7qAi8mG3qmyRx2P+sOxGoIpAIP0a1K
u1+dOD13aFohFUw9OJ3hDV+81KrkrzJ5mPxFSHf/iVPqdaoe9KN6/59oRUUjbxPW
Ity2vJyMWwzNVPWafbbPY5HcWJvDOJvSJG1D1JxSNUqsx4OLip908SZIPm2kzBPn
KVP2ZxSII3GSre5YgB3QyTknbfiiTC8T+uz7+IqP9/QseH582tN7/7bbI9OWF8OX
Mo1Ytuk/N8kN9WDbgjxEqo6JVwxkRvH03KF2Hx6PfxmnZ1b/tQ8G1UG8yuOQvcNR
OKukUGnyyF5Kp3ga16YhDhMxnsYIuV2LgnfLBZhGB0YneiBfUJtT0rq7igVkKqGy
Tlf81/HsesY538xw3UnXRBSB82JsmHFhpyjtyWAeHeNLF5cd5ZMxSBDX73ezSDqG
oxa9WLgv3CIXuC2mLLVGiFApRLRm2yK2d5ZUxqM9G3GDh7QttO4MW1Eex4ENRrZn
974BhgMm4oPQU9DupAfJ2LFto2YvZ5V+u+FFjrIr0w1G8ALHeus4JecSKiqVzVUE
hNOx4Lvlq1ptqPPQPFJrqoNEEtXwUBCII9riG+Fp09i/jgaEzjseCrjW9dTf3EJq
cO1vqz2GuDf4xFznvj1WGYOu1D3vNldvMbaIsJZ2TBDCsgIqzLz74HwyqpNfscaG
lqOYwMp8DMSvoiEOtCCzJPRmzOUPQtkQG2j9PCvQd/otSbxgDJpGQT3eieQRBnAs
PQlnD5S/aERdD/tWKxzUIGRlLW7GVoRdrXyDTdllyKmEBc6HVzxhXPrmE6YaL+7D
vZOaZ1TmPCysRf96BJJvYgbeZkPp0YuTyV93wJ1sEslmsFiisea5Fa7UpctKBmIK
UndpqTZznA08JDaj0q6DW50XmfXJbNN9rQFL8zkzCud/WEetCbBzwZ2RDUWPG1Kw
44eyc2vT6wZ8/mvEpEv6gg1kLfcbo3jwrjmU6yd0YQXL2BbYNTAL4o9D+yAaSw6c
AmRj67+GTHY0mtWvSyuPTXhXStk3jyl13ika3GUDe3Gp60Mr3l3Etah6V9Knk+0U
raoUHVMT6w4BikRyStHeAMGz9KJrcSWMYkQLrUk5AsoXMhLr9y+KHnsJ3k5HjUCb
GVdHPup8Mulv92U4JAqHAayRghzDvgTb1KDF7zZg+7yr8NbGxM2T5jzjANNLEnsV
qHg8J2EixQgYjtc+4OdB+9BSmycovDvp3YKpbdoEN9wS5kEjGDaaeVntvZQgTLsG
P779K7FBUENDIykqfqjoJNST/J8gFL09mj9JDl/yJZQ90Yj6sapX6VdisdW7EHjg
wI8RPWn8ytu4FKyH+iMFwqi5vaH2cq1Stf2LlagdGJc12eomKFCZsgv2m/+a2DHG
OdoPLwmfkMyCEcRA7wexM/kVNefmKlmWDIYsTLYq3mvRd0FiNUGLActiUm7wyvP9
Cg720SP53cE51jgURkXNRSdEGJQQWmROLPfBQwqDPOWMxEdUBZ8d9+wYtqInZGum
Zauf+Hip7VuxUOL6zFzWfhJTUwIRRYt464ekKqAHfOFbd33eaNrmu44Lggr5JlE2
g9s+2ZNZfkHgFaNCpOktvcmza53Kmvv3rPww764gsDH/jYFQZd3Rare4JwflXO2F
Na6Pl+dg0uGRzKjZDW7nwNSxCQprqV5RQ5ilREQU/osY+dr4x1BaRo/QxKXna46i
2MBJT9NT6+BkdRG9AsyvQG3XDFYz1J2bs35soyoZOmtmPWL0U2F+DFe2ML7paSCU
ezYnkZeLaD9503J8VgbgxWhpiW9Ij6EiKj3aTFxKUKzZwFe/7My3nCPbom40jP5c
qVqwnME5vRKKlRUzi37OWaVIOAml8hfJduMf7k4Hp+GOS3YAOPlD7ni2MIupFOFM
UYgp+kRzZpMymkkn4l1+2DAAWDCHBbskYX0DrkY0P2BHTvsL/Sab9i2+SFZif9WU
mtJtTNnm0gclexZiSMHtEG+7p4v+PoZ6W4wpx6V0Si8oVS3awiWKI1i0/naWtiyp
P68t9D0iG6oI6caqwm0ckJguCpV4kpa5n0h8WKu+a771SjhmqNhnDSWu8AwOHYwW
Q40cizyiLtFDxFAP/QbM9CYMGgE2C6ovWzPhp68waC6/fHTKLLPL39+wfdjTaXk9
QE98b3T7WoiNRVQW7j5LONSiO+O7V0DKfa6qLExN207EZgDkK1GHR2gktdLbqZjG
R36a87DiHfJQuG7n9inU/lZESe9EhVXsncisHUpmI4IiFGviBAayy+b+cLB1ZcAx
XFi4WX2UrQzWLoz5lDt/cpDDXMl4qQWd5WmjEYg57Yef+X12du1MUde3Ra08s1kl
wN12CRRGrpPpY8XSJsAqAKDGO5cVMhkW98D7zcfnUg8YO4yrftrqRpIn9UOqd24d
3+4or37XJi6ZX25rSxsuCH0Q6oLrmAR2BqIDKQfGH46Tl8bQNQp/zfcLih2vKgta
oFAPH91MC5X2wxsZTuNmwKahsVqlmcJk94kdB029YZzZgawyl/+1vjVvwqknbeEu
TxATb9mbXc+DaIWBfIhg/0sNIAFRTu813flo9h3fRFQpxizkbZVO6xQA5ZTzZpj2
COWdNYAflK6uOcH45tSeQ2H+vpUzn/hGMHGefGbWUyJFEKYDQm9zSFG1llpm35T9
R+ZmlzbH0L+3Fx4SkGNgG/wdgwJOzaf96IJ82CUMUBOY0lsnmZy2HNtfTNsLWcRC
C/hpfskNoXPOQ7u6blBdgh5kAAz7q6g0vd8yTn6Ck7fgw4tl3GNr/Y7ktxpe+Tr2
bud7tMXAjs7b5joSb4XF+fqiAzvVtVvmCTcDB1k06lOnD5848HcJI1xi5stt1UO8
Hq1Ts9Lh18dpEtJDLQ/atde8pd1rtPhHPYl5ooCWCeKiICEa4vkpL7/1Jh7n1sDy
K4lDi/NwCuFtsUhsoTf93hBYI8Pj09tKhoBhrRkBtnTu+dEnj8l9NW7F53Ox9D/W
ZCIO2wEjW8v1XAGft3o67sOVHfCmD0dCR0LUq+mGTll1SO5dslxvFUkkhPmD/WH5
NmhXSPgwUTY37Yjuvb5Yxp6BEiez7XbFYBpHvbniFjHnXKIyq5KCo4KyTWcR7uco
oTkkfCaSR0oWhpPEpU7oTkX6UfFSFWcH1LOFufS1e+/vX06b/18KdjRfrynf8DF/
aiRIFWBSp6a9TlyxZcjqb/VzfTlhw2iCR4YkPFpTQnwaRU1A+14U4wYbXg4PyoCK
1tOojliQng/VCOYsby6tVSraULEUn6ASSajJ4dfUtdYCuE+rh1JoJi9vstrUnFnK
dIqDfe3HREhTsQ94v7z9KX4Iw6QIITJJs9H1L8ZeQK9JH9VxKIMfMkyU8UpJdrsd
IEUr9kHOqS48AGZ2DLe8p1c1SQE4OERPPPR8SZs//qn93MyE/+B7A2YgyIcA5waS
U0l/6cWlqsHTZIYBDMvhnAkF9aQ2ptmGePcvNcQHBJ9TYY2Wv+qC20+/n43QZGNJ
FJ3vs8iIpW3Wp0eOov21l7pwaMg1GzqGU3M4KCmr7Q5AhcF9sI79Jm+Im/JF5ZBZ
/Qx07sxTsepUIuIE3R8g5qlWzyLItWkK+NU4wAxhibA66rjizV1955n8KLXm/Naw
d4Pme1SqMk1T8PWvnf+FqLwTpf+g3AK6sJRB7XXZRe/OurIskOTbKRDfFVvehRMG
6YPkYh2tjNrw88YLJR5WrOWdOkiagmik1pLXmM63zEmFAj6k0kT7VrZkhzh2bfiC
nxec28wpqdWhf2bHFrGWBl9VD5hJLgdYh1NuDRMWRV/k4UDHtW9xjkpb4yGfWynJ
VMZ1iFW/MRUXbgVlyzt6CIQxfveFFsxsxBBNPh/u7Y5wKwWgUsHsiGQFR+O3qicb
MFc+UQUKNhS51OtIRbhmqJE2a/EK3KWMYuMr9J1YABCJPFisWLTJcWYNwKmZjMmj
MgWzv+0vxQErcnfLujmZXYw3d+3CW5G8VzKvOjCLK+OBzGLf+ansKMsDEEwOgxKR
4rZyIw35FgXOOhO0W9y5peZfGHg+pNTpfBxCP1yDRw5GraO4X+fUdvVkyuWlCpU7
H448pRqmltW1rqJl9In4oBjfFKbfT605vQytw2Johb2n652hMuLsfxS/0RdzOGb6
deQs4sU/K+CglOmaBjzT763kDcmcgOkXI41sCYHyTYb+pYFgeoTmARJKhV/laFV/
Qe/9COWzwYXmpvAwA++rUqih9/XdJ5sFBicRhgzL5CyiGjbe3B4cZjfl36p/CDD0
B28EMBrCYUPk+F4vcO9GWf6fQX22Dh2XQidML9Ev/CrSQj4NXkNB7QayrzYzzQOC
pcR/iwKhxOIXOs81BmNiHUeFOmYXHir+XKUtnhP6xt8eZRHr+Lsg+tzemBpyohxo
k1drdHKZvxlrI0ijKvjNC13pKD6OEzdtZbYxe0NvqUzICCrt3B5DTYAblwjoAxJN
Wox5TsF4IyhIWNrgZc4UY4wueF9Gpo25PmCXgV/EvM0m14+S16EGc37Kau+LvtXl
47Wi1JnaDhSRXZ1Rrw5QhB/dF1JmHnlHIkIYJAlqdFOPdQQrMzwGTjHl30Mmq5iI
pAlpr+xJ0R6ywEvG31LI2kV0ofYc5DSIaej0puxrlCib0721q4fVrcVFVbZ78Gg/
hOxaEWYmMUYIdXYydwfgtpMhjFNPcYRfk91qAIUMHUdpDd71j9KesyQVEKL7o+wT
iH0cBdc53Yt6RZgP+FiKyUTDobHIwsDXiXCyq8vSHptL8LUvrSyr70L8mZuizzFt
ApqMOxe2deZpLaECnW5PMEGG8Rc1rTYYwI+Q4+aAlpnDxJipUpXOiKcYH/C/u/uo
hPO9wjRFKdqvQtGohlwwuIU/eBaEgymsSg3DzmHPOqFsGB6NIIw12wlYo38NNHkQ
PlmR8JEVS0AAnr6VW/BXN4U8LLGUc/9diULcuEhhBg7S5zm2jbbHftP5nn0BnTrP
snESCS1qzae5CgSefo3hAkEOjd02mJo01oAKRbwhFnryvWcOYtuAlvPHMecSldIn
gxpHk1mvvvDLJFvnzPaYX0hM+rkoMgaFfuGIqRxg7tpPRAIVYnT1BofM//NkS5my
ImS+nAVXdnN4UDdZNrw7HIIkKZWKzf6IDlTMYe/mV5T6zBjqAxzAtWeZKebEkdIq
fOSy8smFKgmR/oUcgUUcFzqI/4cUOflCyEUhHAZHE7rIuXCrPSvoca5EFyf+sbRB
WLEufh69DuCoOARihzRMFlzJ5PXcckY45MQLNolmOL0iXFy186Z8N8RxigaXfoY4
7JQLrF5WsRgiOCjhKsLhFPJOIjYBcVVIWGtnUWqcpF+1yUWTlFEY29ye1EbqTf8e
yaGjasm49gQicb7ikCuAghHXmXtAueiF+WLgoYGK4zr8MS5npLMvrCvOwxN/LGf2
VXJN6sz+LkfQjqp2ROeJ6FOIkCAve7YxHgVDrnteTrqq2d9BbN3NLqIoZ02iKPCz
xQY/jF5ck01WKh0kcdhqmWSxvo5AAS03aMtsiBuyvfS71DdgE6J+3daatGM7ce6s
AimSVe1+L0Wn3MmLCMB7087hjOEMkvw9l+YEgHj9WJChRwiUMAj3shYAqQkECM0l
asuayIQI4sk0eMsW+4EBvfMdJs6mAZzVER5QGEtQUcrVO0A851PSjtp7RpSaD4Rn
uLXTmBs7DIAxtUladytDwxfcgEDdGXlituYL9Si5H2VmuhKKPafw+VPWw8MKO5ZS
iEOJX1RlHxGYE2iQWDUJAeHvpAt3QexuKz19fPfQo7XcDZBY3UcjQR9l8MOWDnfO
R53W3ZzF6cVzS8tYXa5KQfyCHOJwpRgDKcydUF8RlFbd6K522rbQDGNtsPFgH/JZ
Mp+y1dUdNSuiBrGihT9Ij3i9nSISIJ5m49sH+IpavGrRmA4RYM8ET8Opku8KBUWx
QteYo6iVLY86UMVMi6Cas4pJbXfdNwzHpxoiMLu1lSfABevnl62YagsXb2ZnO2Di
BcK854Nce6c/gLpqYosMMj5V4FFJvOfj5mdqzh6vP288iEkImDnMxFmUBvLH5NYx
z+cgJq6jV5EEYnvs8RfHQMX9fq3wY3Xly6XEAOWf01BBm/m7+rGKvY/rtfwio3Op
nn5oRPOGduYYon2aJBsn2ElEUHm7lJVIfJcdzdbBQxpdeGk23tndC9vHUXIy28Qp
ZC1LnNWTrY9G4sl+WIb8+y4qWUkxpb797LYm38pdKUBuVV0MSGUzHl+yhbwYqrrs
rZwltkN2qEMLMJy7q/DhzAe1jPgxOzlwXCDDkMn7rzRrgcgMPs7FoNC0hRtTIIOZ
n2yWvqJ8gG5xaKGAY0AIHofZl1mxLF010mPUqyRWIvTsWgL2zk4KO3B7DPxXxIdI
w73XVYup/99r41XCcprpPM5PDIyPYCImvXheMGG3VYUq0HagGwgxjtgKeti3pxKM
v0w9HhEFBGV0yNkSTSGcHS8P1m9HwhPUI10YoCXCbaOP2ITM0VP1XbAjarvpF32e
fkHxjuRoH0iAJdcYhvV5Rh9ogByC5cGtB5yc5caU8Dq5AxBboHwYuMJSvleoGuES
F97eUgAQBc+91QKUvCUBCoqE1IxcOSIdxjheY+fP+IAbQSW6lfBM4TM6oWUeZ5Q1
ZPF9zYamCk3eMIwBODFruotrxkFYqqgDReHUeRhSfOZEUn+4tZ7NAIuKnjKISV2h
hFbdl1sWOemzqybw9h3JpNktHvNYXsFQEqWh8A91tOhU79FGOeTmIisL6exPlzQo
WKihEeTvSmNy1NGMlVmEDkMr+jnSF/p/yvStN+x0DkKBNtRQt/bq2pHjXLzkI55J
obNKebM5YhNz+1nxl9Us6XbmKIpDskqOSk10YbWl0q6q46928sbAQxQmt+6zVBMn
YDaKqAy8anYgF4SAbnFoltgzwtfBtiChxZYbNXGbCJ58q4ES43kkZiilrC2YOdpT
mDF12zAEB0Y4VInXqEb3NN6UqcbEQXLVXi3haehiseUaifhju+uZyV9BBtrjHmxv
nS1Tv+pJHDNz+ZLa/cErlB7xB1qGxnKRRo24UCGyCeSiRe9jFhjukKsnaeFKwnbP
4dZtU+NhSoQX2jgDpxlBu3qWnMhFUBfZU2RufG0GnAcZOw9Ho4o68BAshUX5sIYj
BGiR18I1dIg2a7pgDwgWvRIxzWEmdP5JGchUt/+hi7aNcsyM1zX9hgmUJFZfQfBg
HfoFB5a1K0ioYllMZF55Fz8Ay/3T1rBNo07aWVhxFQiznFmf+ta1kp+hTdcFnHr9
KfFT4COtuJiumAXYUBnJtpA/JQb1kwADprcLY60p3K04AgVwv/xGdm9Ucz6ITw58
6RdYUzwv91c3tXniiih71K1OKksl3AupSnSCUJ8M5RvgAFYRqARGoL9PPyV1PGCc
RN5+uo/FmzMpU2HrQVORDZNRM4sVEY6BWvr2d9+rE1j1yqUkxSfER4s99rdnu/bD
4MTD0fNFbJ84WXXTFkMZFDVEtsYjuSCEi5S3O/kxW9MDghuBbgxAwQiGHfRmb/C4
T+/eWMHIPP9sQCLovzlMT5mujy18r50ifkQQcm9U9BjQfQ1CKklHQVKF0ygEj0TW
lj0CHiy63J2fTrf3UG7aw+6g5ZmUux7y2XhtgBs6BT58kQDoaVhGhSOnpp+o+VAB
g4GG47NOycbzxogEeJeGMNbc5Nq0BRzfKtW2ppTUP7r/Ve0CdLneMjaeZYE1GgAR
m7n9mjkMj0M+paopztjDug0luBQyIDbK8A3SlW8AfWrrRtA1GHRhjyDzqlxKZtQj
IVdtEc//Ole+l2WRXbruk2FyWoONblhTP5PNjiuQOrFD/7pSxu1EDH7Rintzqb+R
ZitMa9GGlr/hF/K8TMyk30QgcckJjS2+PPwsmI4mnHulQi2Iipi3Joe7jHYQpmEq
COfCYj+QmjLKq+y+aZkdKcOlQLlOfKiqv7cvFaA8ug3QKs+gH0XnTMkDzBaXMFmB
ziEbsaZxRAGPW9XpEuOMrWWAYY3jn0Lq+knlhj9afaGzICLjKHiUlejJkSyZET57
gPy0eoAn54V1Zvo/qyyfUSLaZrFE0ytOS49dkG7PK5u8y2x8JPsXJPjv2jtMonVT
m3wYASufWKVL4ePPxpcs+aDPN0jYJyTXIxwO+pjF3ehux5aX27W+zN4TVCm2+FnK
ZrHTJFYCpEX00D+WI7BkBEuhY0bLl82CZrWUxz2Ew5WYU+zFbP+jaqcoBW9ThbJK
5JRWKkm7F8LT/EcYJCBH4dJxgQH7ZTezqTBiyDuW1rx5C9TUrTp8bKTg9lHuy50D
Jf6+oi6bB60hCQ2je5u9FcPGUWOD3C3rldLIiOOCtisH2SHixjEirpIvFEJ+t25k
I70nxcHwdtTqsmGajJhAKZKc4/0HIf3ILUiC18KTbBaiTt+BUu6h0rWz8cMo0IjS
x7xmO5Xg6Go4wtfJi/fsVXLwCllagz9zADiHfq0rsn5VYRhn7lRYG+gE+UdYnXBW
XbTfL+EsyidQZGtx6MeZH5J2U95a4ZRU2MRTfcDfaCdmiuiLJlsTX08TNtO9/R7h
h3hA6TvXUkcBgy6BuFeLcGgZFYwykneahbk5QS7UOpRFoCs/YfKWVZq6/ZeMPzsh
tB6tcikN8VE7HyjP3YNkT3D2zo1yczIcyRVkPFtCxi4fqEqOd3VDr/XlPz8nbUV2
sQrUXHAWulenUAqPpcKWOsjaGKLNQweMuU3ysmaIRvnESrNUURHncTTYh3N8YsmV
ujF29vW+aWtxlLXmoLUJ+nuLHSmYeBrz6t4ZpVlBRotopqbYwCKC6ZKaKJe02kdp
eiX4wMNXCqhC2lIAw/+E2v4UZj2ZlNq3TFh8uS2H7tXtJbHLDngs0RJaZ++gv5Hz
iDESCbjgiQjxOJogrCBZ96lMuV9UR88Kpq00/s5Dw1m7UvBHyMNFs5u3pwh7/9Mt
13MbwUqENFrsxjABs1SC7z+u38wxn+KUhdb5l3LVWgxdaRg7n45TtgjCLw6xxzyQ
aWkC/vgird2ZaSXWNRcATripFjE6wUW54pfByt4zq7IcA/PLV8xtve2TJrlhdPPf
aWTVwaKzYuQUNKC6ck1xi+hnqcFbnUdcX24xxUSzTdZyPmTDBDQi7o+xdhZ2RkJT
wI3PQXwIbnU1/WVpcc8STd+nDyUfOlvcxPS4dZkGRrxeXdoUYNGu3WUrnzKHWoZ5
YCMy6c9VK691pZrnG9+ccrOwk9GGsPsMQqpJnMSSDOISg/+tZgaYyuQAZi3WVTSI
GXvueDasRsMh1/IQts+zpPZjnJ9MGdo36bEs1G0uqZVmL0IDsJ7ABUjjyqx1xR8k
JmIrtd38HVvfR1hqnVVkIvE5OWFT/ZPhXXvXtx7qz2jGtJmcd0ttEC/YX1uQWGAD
Ac4J4V3RRLO/ASu5At5VNyvZTFIlHGMIcVZAXbQz3TubR4yKreVv0jqq8L8zSLW/
E6ctY0+b+cNukT99qIP5sB47UFMGhJgwosN3nvVMQuyZNlDUSuJS8ruipmnxcQrd
NYBZQKw034j5AyKipkueeL9Woz+yGKwESq3qNGVtMDD3kYcKckunVOKowoQSuUnl
+ETvfOAVshHUO/ovvWtx3Hb3p1zy/rt23Kqv/BQ8aI8NUormbowONYJNJdtMoeNf
jxRvtAY2D30ImjFzfK6uPKnLMeT18OPDyOXDfGpUqwprRrVlLKPp/JXCPT3RetIO
X0xbJKdExuSs2P6JKahXSh7Dd2tQifJGcCNVCzuwlPkK64Dgr5RkCAZ1w5zaAZac
1VHJjvYPLZm0ewtNhdJOwyj/11Js6jh8nv9IZz0qrofY42boCm/T2rfO3hUUhH20
5kA2syBHnQ8SZ4DufkhXCrhQ31+k3OJKh0+ULS7Ku6UKjCv3/1I3iJmCvf78qsW5
3BTBdbttXSZUZF+WKBo376LiMWd300f8NoLaGkTN47D3AjWNq0Z9lnKaU6f1du3W
WFK3DrMxCcLEafmpy8N00tP2ThuHliD7qQWV3hOAL5uLO2SAcEv9pbJeMbeFUzH6
3KL+hPr7QVH08y75xXJeCuNlWaDHuT1nNqmPkJ1nXBJ0I0TNfBJKFDCekr5SIFnU
q1FT2dueyHKpLtBJfATsLdbo5rKm11lC2DS8GsGc398auTu7TR0TrjIVSiQyDFDQ
LtCSv1EPHKuTZ3NQEokQpSJ4HHACbtGOsguEiI/q8pGd3hKfOcFv1BPIURi2JrhX
j1xV+YdZpk+evGjasKPeoPBAZlUigZEWRR4MCYGR7MZB1tqwtJAYd+s7zqv9Caf5
b3IqZif9bhT4MRVZg/ZxvtgZosMvLJfmcfszRdHJ/xJGQzeueMqd1Fu/T++Bh30j
bqLLArhZUCHncMHD3DL1RHGHc5ldyY/FMVJjqHlbW6KaD0UxSaWuQtcjjv1/2R9a
9zxCKquZFlb8Lzoj8rpVgmxyleMbI34szCGBGPG1SqhYx9yxoc0/pPHfcmcRYwTi
8TuqB+1C7yUtJ/G67MwfJibpCpagsfQgOlDv/L9us+E9WmffHPa7mdQwDGLWLDfe
4IraHdPus//mnibhnqEig/S6WxY/jt0g0P3F1by4b3UKHurTbI9vEpGzlvCj5gFi
lm+sgYwiexUSkFH8/zHKRDdjMAR9ArkuDA5f5zwxiAqS3U/8gYAVsk6GwpYc/iQi
HNuQODszs3MQ2HXEeoD3iDtcfVJVxlV1zlk122whnvztktIKUsaSevjsGU+7IHQh
g3j4sPNW12lkXA/6Gm7jasgHhJsInJmK9n5NS29hdKKJa7JX/4rxJZvwgJk09V9w
hGY8x3ZlLmuiBXN/QPCC8TY81EmeRweVuRGbKwUI7izHNmw3NaJabpIbfkLF9JU3
U7h2/DQGN+UTogI4ynAfNCI4gzAVuRVXjRACZv080G19G0ttLPgecMwx3enbf4pI
bOYD1qRupYHsLZJF6uhKr0l7HoH25oSgWmxYO5l4w3EworknIF9/UciCOZBdXyub
U8PhcAMsw0ThLB1+HoQXpPjQSZifzn4+4t3vlJBDHOKgbTUqobMqV8yiuN7ypsj6
WSZXz4XTESxWwHCdof24U860r+Eo7g2/x/s/z4Gla0WbRN6YtigVH35iebDzjh42
BJz2uxIpl+RxeBWDKDfw0dSYJmuXUegmjGJhiLZ6R73A+m2f5f85ihGHFRb8BBWu
SQGC0+CdtzJA6nbRDndyi6X0r5HgWuVrGXgGC91ijnyxlHuXpoKhMUE0nFYlQDu8
a9bTa2IMKL6WeT+BSF07NlklcfL7tDs4uuxAtIteJjE3kQL9FS8HnJaGUnDwno0H
SFE7/ZY2ZFxbjAhrhq4eaV3GO1liGiZzFBvdF7dx3nBYPk7K6drfKl+fWlzQ3hd1
1LZPGDsc5WchUGVYOjA9XO998LfwSjahYkn4n59egzAidaEe0jJtsonQ5swqp0Ar
EDaitVjx9Cg6NlkJSyzJ1kwCRz/saEnQDgv0qkSY65JjAtmAa7sfUgEhSyLQkJtU
RiKBrJUAMgzyinc5Ns3GfWYBQ5/cHzYTe0v2yzyJdvfryAr2cFUXYYoEpt3z+x3S
erWVIkwyf+VsjZdJn40DbBpt+0P/6ucyc+m582C+10isFgqzKwT9AZqcmzOiWRop
tj/jDMOKrWaSIXIXE49VFgJ+DxT0h9dtZ4RRNv9VfmGED5Ka1ZUcpw8VYEoQrd4v
Um0khMW2Ly+9TU1Y9/OhIb3oQYHetM+wmIk7m43Ulrj8uip/kkLN/ARd3/Mtu0jG
tpSkZVh9BYhJ9eSqmj6cdaRQOGf5Q/hcosgCDiEF0K+Rm0nJ5eXdg/suq2ZinAA9
5b4NuYr+BHc+MtIvbYSxu4TdmicgzxbxO6ISvDMNRrZLhPfd1nW6voud17m8hNLJ
iQLUCJi4Lqu9TFlnERFSlHDVmYm5rPRKUvqv+Ivm4dhN9roDG7jXPZw4Tb8WDyCY
OVylL0ZUq8zrcpwi8zS/N5gfG6k2JySNSaNu2d+cUDxBcbHu25azS00nEkiJxH0A
J2l/9RKJa9dOTrOrWLwwLrK5SNGIzFh1aFtstl3Q72qLTGRTC+TtnlVO0cEATa+B
WaEc/eyUohfaA/2v71Vmop0F/liPUbTxM5uTqDKKMDUJcqJbUztJn+eIbPRI8EOB
2LXHIh/CzZoVOtw8UYeU6ON06V51PFRu2e4QjbKs+387bcnMwfJaQo/Kb1uDoryW
rLTRvjM+ZEZOM7ilDB09P31Sl4Z4pwlBjx4d6eLwvhiPAT53B618J1inTsLu2KD0
r89+U17bbxbMVznu+vEs6M/Z1YX5q0tABwVGFsnuUTthncmXVJWfkWLK7vYctBFB
4t0flIXG4IO4xCwQNXDvTOAfTenRmquz6xsj7pu4TAer9ypKAgWB7Xju9Nw0lGt+
4IMbNtkodlhBVocEEqBvZRmgLd6EcPDUaLWzM28Pf6CXZEoKwRUm4xY4aqpFp+s0
g2QPk8Lh9pAZuJbRE/S+hMf78U0V6jjmLMymapfa8L8F4y84EViKr6hgHqWf3VhW
P+3Ynl1lcGVzLzr7DIw8iazTETe82xPSqYnuf0T9zWsWc9Mf1VlUGhpcWSFo2lYC
x+WSW6ydI1fJzbAtzMbO5DLgplGymUjxF94F2zJxXNb1/wMZbKqIydIo/bgY6Xpw
NdoNfqiThkJqC7e4Fk3GnuxsmcR8munP8KNLrSYGIu2y4Hf+tYP1AoTfUxRTNvJO
Mlu3VnaB+tQfkxqmevbgf7FJJ/S1lezTHH4c65DZIrWiJ2Tp2nm8/Rg/2glo/m4q
AKmZv3Q+RxmXbtRljNzBAfIgbGOtcSY5etAiuRsd0ekUIiMmkcu3a7W5CfmKY6yk
8AjCyynSCSdwiGz0DQoufFfgya1UkOOw2FQWyfCXDRvfEue9Y93Pb6QT23LU5n63
RkWv/7jufIOHfRH5V46TONeAPH8TGvIxSahrj03pVGMujzfQz8YHt3W7NII3AsUJ
r8BD+lUG4dMoOqYNfbVlis8UBzn1Kl5fTMymN8lc3xfH4UETDrVsho9tQz8oaR5G
s1J5smHBbY1TZTMj04Tsdh9pWGMqgG5sDTqyrD8/eJjaDAYh/fbUbVwGRqBlV0gs
nfK7y9uMBzTDCZMYHAl9RTsESTFtbxH0iKrBNhLJEkBfjt6zy0z44QqKdl+5MMRz
ZUC1thnmuAv8WVXJP+q2zCmIUpzQIds/RqjEM8EdMFi2b78bo9d9b0hMTJdG3wQX
oNJcaG1hqfkF2EW5rcCXYWaJteSlbk53g4/E/D0PxLcQ4yq5S5zw/zC5O9emeQBj
zjMwr5JF0y7+Ksw/XsLbLaqtDGrIEulsEA3cPFWLpPaKkPtUdF4fx6b4SJvEzUk4
xSBlgVEsQBC6awCbag2iIc24/S9GWRWw++1ki2TMN4tI6FhnzSCkYaci9ckZZzRd
7efLa9JRqjuAWDWeXyHhLM3wov4AcGT7OQsrERFlOwc7NINz6x7FT7U5/aKVh2EX
lzsYkDCCvrxlvBtwRwgbPi+2qYgh71nEVpUDNa4D153MrO/A6XJXlV69ef/N+d3G
6VsadZIkAX94eYL209zRpIm21TnkQv/HDn8gU0UP3svIzdttK4IbQP/7qaZg4zBk
kykiNo9eZJzAum/Vs1SSdQNF81XlhIAKaR6DEMcvgbuSRuEO4dPPJWYdPXtCAwEP
RVKyA9xbyo+B4Eqb8uh9Z3eyv6LdoGBoiq8AnAfWf8E9icfsGxy7cna8MpBqinbD
r1xArvdXzn+7aQUmgqsd87aw1sv0Xjxl8prpNtYNwuZm/ZxuQSoWuozmTS1fe+Z3
QS1MWdfoc237Nn6JnVWrdOoOrB/uKtGVENPR9vcgQek6HVKQVpYrY6CKUjitZc47
vi+kLNyhHVeNQ5xq1aLUdZ+Xx93a5aLMIbUcSSmutCLsYSYHLnObhB4wr1CAPViG
1u97HO6EmPmum7HKdE14FjqptxcH1P8MOJ9WmIAdFCOjTZXPirrrzPqsVEHQ+t4p
Z2Siemw+nrmh+I6RLtKZaHH0BpHeeQVYqswMwqI2K3Aoyg80iWIV00v7ammKOTDE
winslajUX5QApTm5mgQN7JO9q204h8f4m4sTxCvdKoJToYRAi/zAzB1OkNc9qp0m
8vI+DyGeA1HjtcdcRfv3xRlC8IiVgcj5Vvl0KwxSD3Qnu0pigQi4UWkqhmFSLCNz
If2sJuXxPTbqa/rNjPA0S58nlLkfyZarfUr9j+6JgOwMOep9EcdLLJhcaY5GvBrc
AFXabyc6mjWl0Si8E1mxMlnXJClK1e/rmvFDQlZC5ZDs/P9wcNu+tmUWOiSqOJDZ
C+c97GFXYKP0zE2G2QkFCciejsi5lcjJ/VSDauZOf/R95a2TUrv6HUjPLXcB7rnJ
Vxk9FulvCf/Pgzp213XqPSqUwopZDevpywYYJCQWqEs7PpWKvXJKep8rx4WVvoBO
5Lh5lFHXeNWjPNHiqGj6kYcv2gKMQoA6GE7kz44jasbSnd8hceM7jcdALi4O1gq9
Dq2IHHBhGxc+beSA4znVBPT9I+tmCvo+eDE4/QP4WNjuI5qt+tr4Dopvh2lzQ8J+
5djFksEQXv5u8SO+VgHYjGvp+l4WriE1GqtYszJ6PIj8d1kCLdnouCCnNHzTgH/u
ocwy33dFMeDv99O2m+3COSOM2PTLPO7rwKdTSQIEbIPuk4fbeioTRrz1HjVPmHIu
/5jrG4pcWALPq52kdoQTNO1c/du4hXLEFR6nwkNPT/URQyTh7674ht+0ALcp7exc
BsibHWOTTvbJLlIhMjPEPEW+M23SljvX+LsIXED8K1kPSpBQ27hAz6nRquK8Oq8w
qFsAzASpicSL/rA8lhHxSN/UjdMCLx/leu1hJrl2wqW2AfXHtT/ZdGrXYLv1CMlz
ZPR8cwOBl4OkC5iWZ1xQL5PeAnMZRjV82ZbDeOCaqTRDa3fugLgbHzBQJgdMKx1V
O/OZ1Hny5inPtrGfvwWyLOpD6NYTBU/45bViR5UdEq+cumzBofW0Gk8VZhLo5Amx
XikvRymDUZkvloz3Yn6qQbe8/Zvw3iFjphvfwT3ROXdVS3JNayME3o0RYmiXSK0T
exw5AmUc0zayOtbZROZs2/uJqIylBF3CutvGkzI4Dz9LnUFO0ciKSy09yqVVerBa
DmSgqxQX2AAR9Lt3etA4onhCPCiB/gJcbdEoZ33WoGGYLLi1+boYbRIkcuE/Rive
rpbYWDU15C4zczvGV/zMFeZl5DL0HXp0GaZp94BYbYMYJ+qe3ZpJONq9q2BytC8z
ydJsx/HxerTnFCIbZwTphEeFp5HzW9d1EqzQFjxP3ElYpRO79MHuSnaGzPqtHpXK
1EPIVDnPjL52WHduLxgQaVqKs3cmEuivvc4Es62ch6VGR8Ssktcs6JqA9UacN9tN
i6dyIpJgYrMbmAvXAdNobImcMzRmutB+Of/IJqb+DwM9nmVvciQLXeyDhaJvajkE
hffL4MmABNa9HiZ4gr/zQpg4vIz375szVG7w63hrF5Ql+jrsK6bx0SpNzAzLbo6o
oqsRyXe+ImhSz4YKf+70qFA6zhYVR2zwBqE6P/w9MWhTcso+rSua4mfZ1buoYjOv
DUpGUpjVwtKFecLbkEQFbk78A3P2k/pTO+tb4wOsnZTwgEo7fu9RYxe70BO85DC6
d1AFE4fNEgzhz636TapYUtVagf1HKBEgvgr6wXsOqiIJz5dtpzYyObsS2/iK5DLm
Uu5IAoruWhCrlREETonCtnlaKODsjyudPGNGXYidganSaVvKjIbDko3yp0TnYFtj
93L4ThLKbY3uTx9aJxIcB746RMD7hCYhy7bnSGdKS7plvsf/cwez0g9vFU0ob3mS
RSUdCd3G81x7A3xpF/CRfNzGLmZTSuKfeA++/OERp27E1xsExRAolJ/tPAH3/qz9
Y7B3pgl2rmk/10rGm0gbSSbVQauQZyRGCDzFTuiKuk8I+Ypdtt6Ad3Dalbo4oiI8
BmZJ1Z13k78OelnHOaMqP0prtRUtlC2XwVXax9vwynD/6A0nk2JliVF5LwCqEbJH
pdv39lAj2YIvigoWIaDpMhpTdVOTBnaFPZEmEfnVt0C2NiL85TzjZ3VhKt6Hh01g
ECZvoPhsBgL+UpOhXVvt3+2p6ynVJgleqD9oy2Mgf5fGqxwdmehNRbHtrFDu+mnQ
JZ/po3QlZRgX2H4Itkz077nbhPzY2JNAM3/DARNZupetOC+FrqxZb3o9p1ZsonNk
WqLm7gHjt86Oos/ByZq1jGH6jSlDdttIIQ9i6k6tmywB3m+ZgQVY9b70LCTeJf8G
FPqmtjMk4FcDJXHTtrOmVMVs82a1G7zNnSTwL+XW8G6eue6vuQfeu6/L9GRhph3o
ooZJ88BHTE4SI1ELgFUbeLwoANSlEd+asOJYyqKlC32pl8IBXcRZ6VwKtEnGcHKB
4mgGAt1XfDLjPCTzFxsi9xyAoGV9YaVp/Qe42JKUuoyTPRPAYIL6AR4wsTHxSBWS
JZ0QJ0k594dKDA4fPj5XXF11fNo1YFaW2wXv5GPJea3n2KVUkPvLO9LvzuPzmy+A
qT2kBSUmgNCTvatYt4n78f6IyjFGNOJj2UZRoFqZbglKvKL32Aqjn4lxNaoHQLpT
KK3wjmiN8+346ILjfFQUuMFOhD7rpPtT2eDS34y4sLHF+dVPF1iWLJ+ZsDo9q50j
FrtlYXsGcW0coAvHN0J4kVoJwC5AoQAXgNfVeBWC8jqTP12ZqaZj+tDcQEX8jMsE
aTFFIix5TIfWj2NGf9Rr0LP+rRIIINmnP/1kGC1eXkBqvwsHvYsHy1tfXfAJdz9G
WvOMS2S3S0uJ/rfI8QkborSt+Rkvcfaznlwus8z7b6B4Eurk4HI0XnLmxyM01Fuo
+3jBns4WoiuInapOxnYIPdxPVv70M+IuD3Yd236WJLoTKg8pLYzXfHIQybfF/N6v
/y1EcGxcIJrvHsC0L5ZZcZVhJ7VwN6yEGO/NrCNoynKzCf1061mIhDLN+x3yd3M3
UVCzv34vPldTAkQ5WN0XQD6O0j+B/MVoKGQ//g5ad+4umtS/WtPWhG//EU7hsFMg
XWOj6mDTeGNN2O1HKc1zt82gJteCS8RpmTV9TMHlPbIn354/m8gvYJNH6EdNg/zt
c7C5WUb8d5ARsvO0Cg+Zvdk5mNMebHZh9k86BouodzCbXeJdlIJimCCnjI5A+BXe
cx0Hr66r0H57GHXvP83jjEzMYf2YU+upUOTS03fRsGLaozdo/RKKVgwRxaR8j9H2
3aatenGS+j/MUGPBTTI54dv7rVUfQGSNqgRHBK+McD4dlxSPtibjonB/Kdi2x+ro
u095SVB3VxNC5ZgHstnUDFYyH+W6FznaI/VrN7ZuWvYOJN2zoSaQrSELk44+Rn+r
VqZgsJwIvfylqS8o4nJ1hhOiZeOXzds/CfV6Z2RFVfnJW1JnV24iB2n/Yu5tKD8R
xvEps1mDpRP4MevwcJMSyb3twKS2OHb+xr6swSrSgmFOJ0Y6WiWbNQV3cjmnn1B1
q2bwD5bf9EcD3mHfHAsUk76BzRZ52xkE8rcACHY0npzubbey1bM5R0CvcpxWQrxS
HhoRchTv2Cs1qMkzbdoJML9TVeHntvj1/A5LgfXWfNb/hax7my1IS1Jez9MUV0OF
stlhw8CjCC/d7itHtykMEny7bn9UUVRn3F8hFxAr94pSEs92iQIfkiS6SWZSfKMf
8cZxsCWZUhwNi1gbzIodPgD5apHxy3aPe+DrsFMHWm7YlnCp6uXTW8IN/y2f/CSr
jW9vgfx8u5vmdHMG5SvNOcBAlZbs3bivYe5QkpNFAwsNyhKzlsOzNLEKq8UFvSAP
hsQEAeaKj7ue9spW2V6I9g/yDGwxsLngSsfKfRwJPQpWPAzCGWi+traYe1PTfu0m
uhGKgyOlKzr3DeuOPoW/tH4GvecHYdiWuOw0ELIvK8Yp46puW81ZlM516oCBB9PH
/PiGQ0C9pi4TNc3w8lcEXf7rpsnXt5gLSiGbkEqfj5CkUfaAa/lVuYcDonyOcw0B
DperNchFA+y6pzsrMSrCdsxNhu7gmBXMr427c9WiGrTjJZIaR9xnbs+iK/puAxRy
oyafKxBYEiwGmujzXV656K4qxfS8MNfvXEipZCA+Dszzii/H1NV7d6aelrpmr89Y
Z/divpJW4bbfwEUMV/OwoBcQ9zm2V0vweB5jOOl6dr9g2bMFOIeTcIP67c5ngX4E
RrVR+3INz63N4mtpXoDNU7AiZzC9V5QjrvcC1Ht+76j0CNwyntRwysV05uxja8Zw
ipgQID7M0vF/rtQ5LmDb0W3FyR04uCDkwWsVOBTqWYyDW8srFW/E4dAFyKFUb2EG
LnjFDtHwjT/gmSeoUqpEnIZQcOMHJe16SwEAoKcreJJiAnW6QxnlfMR5wVXN/6KR
Trd9bvRdkMdPVVrWmOJkAEkXQRU2VG2WhPsOIztXvrpyBi0ofzlAjvldTyFU/qoF
l0jqBtnexOqAa5Jzmq4cHboMmw9sikO00kpyDPRcXsR3CQk/wQyHF69ARcoYwLTU
i5/V5S+bTY3Iu6GdO05ORBMgTF2xDIGCxsffmss0YRoVsQfk9IfJvbuXqd5i2NWZ
LeptTsAAGELb/C246I4PyR9WWd3ZvXUgyzxYCHC2yCHya3Fv9ywQ98PHynyKzAcR
oZwUlhfRcu+n/3SzO7U7jf+PPwnM7E3Kbe9989+cBoWrySxnGKI0D49+hvDvoz7Z
C0qlb7i9dYRwZt8771K9OCQaxtcTqO2fVQQjnveDp/2oE9NOzJVS+l1Rs/DXTYG3
pvBEv/ys+lAfq7b70Q9a/9Xdq3vIG18s0YiKJk7PQHyiEo4ERATQFgK6i308hPPH
krL2+0UeIoikP3Fr2NpbFZtWtQeqTZq8JcvO3T2Z/0W+I+NmWdXmDAKJjCVQ8vje
hUHbL0Pql3TLHLKGgGEKtS89HjO1NWGaNuxIGw1SfBImYWzuVG4XOGF5dE6h3Z0y
4SNEeoYZ3ftBnYsstDAirnho/rQfKAhDWdbo7dFettrKCgKp/bK2Jpv3wI4NIWU/
bHlrzCYOlshIaotu13lg0o2uNJLTaSa9pHRl33OPa/+AKQcINe7Xa3j/+DxuyfWT
pe6CtADNkCXHohHXD3k+j2YGyjKzhu2Dwbqx0tk2iqNZnUOpwpFw0GLPPTTlPZCD
YrEHfUJm7s+VpvoJNiwKMsM2bZMnHNQ1wr49Fze+D8JLWOp9svsNP2Lgukt6AwKl
1slvQ/JoP9xkteH+v6Z6dXW3Rv5zwhks7ToFseG3G+VYrwGR0QYLLpvZZqdBQfLV
xGhMjN/8WSRvPfpNE/tInNZQ6I+B0JOInjjEwjFgQGUpSfYEgCXdclzReTpTQpqk
8P+8yZ7+mgMkB7fkJD9GK13Znrb0UEQb/3FQk1plZYAaielZiDv4vXlECcTW7pPD
bRYlw3h27oOjIzgfxAxZjp5I75C4CjNGHqt5/M/GltmZ51lxNXgeziGjK8XzGx1Q
J9mTpdC0Tv97MX2Xxcj5qXqjDTOOZZLAVrwhxqtIx5/WLeFjaZhGpXzNKnRSafAN
g2RNzjebr4tpyx8DMcwYBbTCV7ntw+qGvf/SbYYwxzAlmQkj6I/kLuhpii8B5oSE
muojrA3cEGmfTeIhCmqcBE6iQ8Th4tfuhx/fo14hLywUE+7zGpBjh4aFJ9ivo4f0
p+IxcudOQsykJ2aBnlWihjgXr/+hzfP/IokBFpfFagVfxi9jmESCFrCzluqiVJ66
blk37Uj5cmIPfsG+uezhCCGzBbUhSGJUoUkC2o1x4VAMCvfDHCB3RfPRKODYgb7k
XePPvHCqLLkZ0jm/75oTCbNziwmW/6B5jEQvaeuap9VQYX08pmCK94vdaQRAGqql
mv8OhRBkCPPd0OU6QT7xFvEDFZNJJSSkFB/5rwgLGOsktCOzfLr2XOV05Cy9gR9a
l/LGFtHmbk4NeArKJ6q06GgyrFEyANUbbwvnhelJFVJzoslnbMjt5FtMEMPQ8qR0
HV9K66N1cJCDBYdx6shL6koqDgX6t36mFBlrIUA9dJfCJeGpiPU1pQs3P5p3d98E
LwO2rkBHj7Sni15s/La17EEclayMkNztNoYJFuVtOQVwv24V/BVgGA1fkVqh7awT
7g6UpJLCxYR/L+IAb1iATyfKXA4HeTeojABBpYjNQ6WUC0BvESm9mPZQpMGE8eBg
tVTHaxojzCQKM+um0a1KoOTkFmDZ6ZIP4p1EIAEHC2I0aZKexVdSh2034vNms7Wk
smPAh4XRBjXiOHU/DjMfW41flH90nyhw+UG61j/Yaz14a2iG5nCFZGSdbMX1D1Sa
o+LoJtQ53dehNjFg5V1PoKoyK8KQtqObWqt1Wk0w8LWcehgvYwK6CBLtW1zprYmy
oPI2oCrSYmOmY9Pjbp+hiE81AVn23X8eTDigylE+ZhDWMx91Ji3E+55MGd20qboH
RFIgXdxYQRQxQjY+XeKYzrM6m1k7tay22YJ7t1U/aT7XDSU+46i1l8baygHCZz+p
43Mv9yrELBJPoVCj8uGLjI0Z3VrBnFKpLWL3I9iUzr3PaNCeRBZcV+C+msIpX1FD
ORpOkNqJPD+N8+wuYxs/hCv0nFPT1EoNwitybu54IOl8FkHQlXr7dpdAIUdOqDbN
WBnRp7mRjDB5rz9QKTjKNPGl4KDQGbC+9aroFmWdSnYSMMTCRluL3eIAnHPWkw4n
ETWnsOcM7TS4Eo1pcSJwGI80S/qWpXpFEtW5/HF6ANYa5q8fGKX8pg9d8711/RCe
dAyQvRkAWQGnFHwoWQ1QQYJ2RUs6YJwo1wnGCq+EBnQgWL441CqhWzFVsmIIWMw3
zGI7ikdmxOIrXFCoVBYbiZqe/ZEhhpjcNGXF1mVF4yFdMa+77QeL/3KvWziYYaHN
6V+5UZUaKNN7Ze9uFqN31XHsH3MAlsshTbHEZoLwDq7ZYv90V3l7/oc9Mglm/5mt
O9JlLEV6Wub2VMH3XWNO9wKL7q+yHOBBxEEiMJ7dGuKZ9JWCMvWPqRmP4y0gNQjC
3E7dVhBHam2TT7Mt12DERFhOGZcTrvKPX9W6SIDPBWPyw/6SM84RE+V1EpO3wdqM
B88iE4juYH9onfaFOOcRj0eiRlToO9p89OfchXu2/X7Fh6eOXKD8qljpkEpBv0Mq
C1vv/TCjE8vrjWgh8o+NvB6oHJGEdAahWuzIWVjrD9xguKA4/YFmnkqVP4xp78Z1
g+xQjrHD6cuLaQmO0d7Z/tjI7uzvobSrIiTw4f/mbP7wLxBLQmUc14+GlAncOMsU
woPhVJrCulUXPIgR1bpNXNRXoTjzTHlPOt7991bxrXPYadIecvejDO13h5F8MuSi
4+/2JxkADJjSDaeo0m2rOkJHoEw/msVqkbyLge/Pwta7c+mkc07646q2uKW4V/hR
WsDMZDi0Eo9jgaRhvTNAO4XhmM2eQBooRg6x0g9T+sRMeEpZ3/Tvcrrr+9gB4e23
DsZF5KKRPNoc/PZyTasOmfaqV16694VgcpGxOixM0upQyOE7OVtaPY3eXUh6vzbG
IAvOR6vD3dtOVQKjBtjOD376nnWkhL/5tJwUIvTmq0uDVC2mrC8BtZy7+LxZt9vF
NbJa/giblnAk9CA83B0hIa/di1cCLi9REXlJn/nmyecH48VJ/9Hb3KxI29YwTIzu
+AFC1mcbosQLrxJZ4Rm8q5gqWV6HDOYRMqNk14BQO9Wr1JfsA8FCkA7yGDonosmV
5FVIU4fpwrUXkQsy9C8hBz2vGbfQTl4QHHyaupFBxKq5wFgLVRoJnWOCxgFIKAlL
fNdvjfxFStoyqyhrjbLygEbcKsf9XuYlgH8kP8Od1g5iqQIpT1FBwVENk2Md+ld5
kqcACG8rEg1H8rSh0c7oOcVP07eO3KFj+r3VMKR3Ml3/vRXRLI8D3t16pMrGNcL7
FAh5Epz0DX/BQfinDWhMiGGsuyfnuOPUUGQdM5U4KqebdOnYDAiTOkHfU5ugPO9y
vvIBuAJErp3H1PGhDY2DJeMlrhEe2c34640QI/cOR2kEd8QB2UU4t1ls8kpw2ZfC
5YFOCA5O1ueA3YrTvIHmvGnWukcUP1FpTmP2awEg0/JwoLku3K4xaC7tTcG/xVu8
CsV1xiQ2qw8B5OCHqypCo2RyFya5ixf8fYoSxfE2DDVAq071bQnqmpZFh7cgNKa4
69jOJUx5sLqFodchSa+G5iMDq19XPkL63e55h1ToG8KW42ZoOhSyOlJ35PFhe5Qe
ZQc60t7DY0SgTnJNbRw9+JL3VCZZEgSdGzu1hWhYOuyzjpHOtrbN14lP9omxLcuG
L2fHwDeH1JkSMO4Yhei2PYhNWFXZrvUWLb15anUNvuQddKfIBQI4y+5MprbAjfNS
TDois/+TWmwjvvdsUnB1B/wR0QlPDo4QerBathS3uRVB76iPJXG8r7DbuuZ+oY7v
qynGeb8HJBeryyBNgbHI1vbGnbBlHgB9IaQznQDRw/zZWGGCJUpPeqYAjTFzKJC/
y7VrLTTbq3YrjhWfiQghhJAZUgcO40EZ/yVRMnityzvOXyvpaD+7BMTtYmneu1QN
fbGmUxoMeXVkTqJbaUnguB4rM0g5mKdnM0Pje86iK7/Fa6KG8T8cr2Mdir+eXRkX
LNwZkU7k8Kb60FlsWaL2P+TN9kUIp5xLfFfe5HFbjz9RmCroQtyXtBSI0y8CyXIZ
ycjtWU2XxUY9oqn8peO9VXfUZg4EFB5SVjK8gBZSjU7Gs/51Wpcjq6nNzP6n1a/T
KnyFhC7Ke68VI65diPud7yLD33Lt72rF7xdS4d2rIlZsgsYqwxWhabD+XODdS+rQ
//NVPVMvCPoMXjjQuY09qKLVWYgi6YXVR/RGPL01yjtUqe0/o9Mt+qmCJfLnw85C
MyldB9b/V4AePqRNgFYWpKam6N7E02WAcdGjk1N9frCogiCVDr2BkHXRQDLWBlts
Otdthkdgp2eUlTHrt4rNbT+wYRBE/eic2g5NGTMdWEw6nSRqK+TR4lDjOOkxQHc2
QVsUESMg+fTgoUO8+CsDWLo05bAjW3MvFbq7nq4YJGETSFUBVbOuI+uCHgu9QaCb
rpsfEnNb5g3TDCV/7rDi/3ZLRUcspy1u4DMqhfiDUNB4lzWk/fDkHSiFaXbkX6ZM
u7sdCWAJsnkxITFSZ6mUJhOmPvEZfILh2bHxb+ZXnVDT7c/6PMM/HWJmBjbdpn4G
nHI7kgR0hENwgqGK4t+EfhoJXA6ghm+l6NLei3+rSNiHzL/Z0T8mEurbAmgMbROR
OV3Ycs9u6Jv+xXFTJXhr/fWdHWFg7Ja9A9rsqPJ7R59Pmu3U5RlyhfQ8E+V53Dge
3rqkDdRJQMAWNfOacTTQ+v7yd47G/MI+5x4CnT8Efou06BUqp7H5jCm5yifVia4+
g6XJeSFJXxEnwTF9SEIwNPwv2rT4hU0A6hmS9Qe36m3rX3oeik6vbQKm3AqSznk3
ab7Q/ur4/SIDbm91NR/vI5c7DJi61Vz0oke2s2/2FaYfrFAcYBHMyJBapKaMEaei
hiuR8X3iDuDhiBt59oSUxC4TNo8FKkuZgY9Vt3NsWJ7IYTwWYaRgkcbAsPt+GjiF
rplAstalJepCf+uD8qmQQiheqCWnOdQi4tc4R25c6aejlUX6h1wLn63vWBOHugVR
VUpefBHTYprKcRQHVCcYkpFV1kKZCAranu1jIHKEZl+uddBNndJIYLCKDQ/itKFI
9vigCFin5x/6HVrI+e++wtZ57i6InxjFMRURSqsamEv0ZJH29HXByIz7VCJp6Dki
0m7E1Wck44913jTU/W0QIB19iOtmgxIr+yFDu9282adzFulaFxgDl2bImvZOdnpM
mp95KLU109ToNxdlBv6Bt7CaBtEqEDzeA68utQ+T9u6DpGT0XRVR4pEbOyLjHdSa
v9NdVA+chyq1oa/niOzlSyqc88hnHY13ZYu5tkM3Yh4okq76KTfwJETUzRy/sVWt
ltVoInE8fmsmgR8DuRfH4bM+Jn9qfbYe2YCbLvCho1jP6TiHwn1Ji0s//u511t99
Rjm47esJ5NEl1PyEqz/JHbcM3edsO1WeAQcqoETGWEpbcGsXKAEU5VtZ1qxnhS3h
VROS8s9fOKdu+n1+Y/MqsbmDHpe9D1Vx/yA8WzlnUZOEt/dJI4+I+WLjbZaB/6pa
tTXb01pumAEo0M/Zg3FmjC1h/ytl6tvU3CmvSO4efLLAXyhzk+oCW4xUaFGl0tOh
KfVqnK0A3BH7tTJJR9rNKR8GdedF2gIwAnW0W5DrbTlrPFMEiqY6Yea3vpDiE5UD
1XZ4GdYZ8S0Em65KMgXQZUn3Hg2+DLOJ2MCmfQjUCxUbdXCwsdh4PVB/jAYttvZA
LQbQNzfutTqsZM5z4AP6rHb8SXOH5Vc0G+yI+PV7FQkKavrn+wYJTndxZBwjOX0y
PChwNs5ndc2rCtlNk8eSm14cYogYfonCwFQG/x25P8Li10lKIx8C1gUtnPVXCRWW
zu2TrqXInwqYjGb0vCVS4dQ/NpeW3ymly/ikqEif3Mu6PGz2P5ot87usnbgEHi8U
WMy9SE2ZWx23vX3NgVznM+51ZJbX7hc4mmgDWwTjoggS2XJ9kpn+PxZ0cDC3In/t
Xo2vcj8HDBzG7rK7qjWduf9BUcuIHjP+bNTuCN49h7MavC/yuZuGMNI0QJ6y1lxg
2ICVxbun75UdLFq5tCq7O4Zrm9eBFTVRxgPFyNaNokBOTI0bag/e8UPA7btaXhzv
TFQQpXGM72vN5M+x1Iz05sxz3va1MvxMBfi1Vb5puGpHwGARRzeVAGd4o71nchRo
orSmNlRXkbaIJXAWPdWvgLIGLyOOS0Naa3PnWAxIYyA6UY8flRik0H2zNibRMfBT
nllfzV63sRtS7rphiL6XVkl231jsrSIAT8yfM4DkuEenik9F+CfoU5xiPCJ42bkb
Nvn+PYGaONu9LUnEjKGTL9YIO1zkHYkMEW1U8PsmZvG4SWRvy3118SCLSd73gJVW
/dmwStpQU87UufzHRWMHOBZb4KtFfA6r9jZdduOOf0rsayaqxPsaOeDyjnT3pbSX
/rarx3jW56WVJXpxulqswaFGP4guS1eIo35F8GuJoTLs2feC86ow1cuGnRWIST5g
89Qaqdh5BIuPKe2A4jFI3f62IM1/g3qLq00eqM20gPdBjSEi68/f2yt5IExu2P/x
vS5QkINrXO/Bp8MWbkLTkMpfstmXdZLC7/XW5XJrEJVGZ4pHUYotMSROM3lURZJv
WmUe9NFHEy2LHowS2kj05sq14PEz5HfRyxhTnrt08IRQw7yhyp3yD43/ctWLw4Bi
zNOxLidGozCoiD0yH8KQUan/vZlUO5KxH39SArhMgQDG2EuX1x6kaKxurCySfKjQ
t0yC96QZyz3+MS5cjquqZas+wW5BcKDPYS7QSwFK0GsUEohmLSMTK5zW5zBj2pbN
edlN3JRzMotncr13ii4fc2A1H0gFcyCt0kewvYVneMD+5zp9LSfIKAca31rQ+SCh
ooLgd7Exzv07XF5haTHRLYQxCnAd+fDw382JkllP7PAXu2GxdF+TcZ368CzQuUY7
aiEoEGyMi0K0V2M6wQp3ML8HVzDtFAR3uW7XMzxMIQCULSQp0y1E3MJMzRRFFCkD
stwOocGAZ0rrL7H0J3j861WfC7w0+i/SgUSTsk7kaJm8EcFgZGcEOEBYZjP6E+lZ
p9DKZ2aaarWEe4t1MXmCi9GbChv0rPHuAFXf0xMO/lts/KarL0pHJy3MyRZvpL3a
u/pPgGv+t/oTyrojEwbvOl6awAPGWPtxzs7ICI1v8u+BDpp7ZvTMewDEulz8PyF9
c/BFB9XhmHajVaiVc7ddBQNABgn4ukOQGmzVscgcZMK4B1LfkSq5b/O7Bti/7Cn8
oWhU3VWXt4+xjGkZld1CAcw/eT6Jif6iQAVB6HdLP5x4yXCV4uPlNI/7xho0xhjs
5yBMb3E6ozjAMX8069MiBgNy6htwB1xemcu16F1UikLzD7UxZtu/F+nX9aYTuhVH
U6M2WPs6wjnhK95lsJ5wJ+lplicsdAnFce+qGoIRQzdN/ibCo2aX07fcMVmO/Ff4
eqbNk75VT6lSDbDp6vdyObUYPGg5LocA1jJTqhVqQl1sOW0/cJoM1Jk4PF5LcTBK
cuP1TZt5GXdnRo5PvZZ5OT7jMPZcGEJcf2NfYLqAD3qvnNvdziYw/6fZAbpPibuK
u6ljMy4uL+7lguxkzA7X0aI58g4b4EMRSiHGwYZjMhdQ33pYuOD5wgAuX0NPQ8i+
3BmQXE9FDs1JyNIZQWJh6r1zLkTplm2lWbE1eAExi2CG5EEwsHPfC7HBc83GEVj6
IgpxhdWH5UgoXoVkWHWQMgodWaz4aXp1hkOYtB9CsDVR+Py3kC6r+GA6xgtRk90L
u9alE+b1T1HSEbpO7tRk1c4siGa1SQz9tKrtiv+me3mWoI9cy4WejRGCQimyBeRu
/Fb61mjcNKPWOBUotZatzabCtUZbfB9RIEQxipWSorUnsGiUdp4WYp3cgf8zh84u
E5gdylm9vqfvebA57UBzEvWC/hMhGHRuuMTp5La3Wtx+odP+wr1wuPeBqzF2+eua
R8I4tPZ9jSmKo6mMuSBVcEvAb8g1f/lDxtVtqnRry02KVy2B5Qz1benr2XhnohGC
V9uBkZw7PjK6Wl0twKmvgXFGmZM8s1AMvlTvJBHqCM+WHzLeOCWY7XfNeZKTyAuY
guBFYCItwP3TvJg4P/8qPabLfFJdn25IoYEZ76N0IZP5bZbIPOGUYhGfthekqSfu
GVPK5WXPT8LED5OR4Y60lILbOpeDFb2Q1iPJGajC1c7xbCE1w/qU31uaEvMDv9ip
XXdZUVgzXis6KTi1dsHv7zJCInUgvwG/dNdnu4N9HkO8Z6HUC5LC5/JV7BhZB8Jr
fuhVtvYxdpU6I3TFpBNie2FcgvjgbMTeWeOeo6cUmWIwGmSa09QFMauQzBsuIFrg
SrouEYsFL8R7/3ry8L4Liq/wLtkGhPsxiSplcFD8g7ivibsZEMYAfnlJKLpr/en/
CHWG6QtDv+XjB5dTtqEbtPUejMSmWApQdX+Tc/ygOZwObbfEUkRUsVbsFEAsx4aU
HJT0YhBYreaJX2UhoK0+fYu7Cb77dyVlzNcRbtouuZgCo6X+wHm1Ptw6ZHg+h91b
vczlHIxykB1FlxZXmCo86lbH5+ZB2FZODfOblQayKt916AfnQ7GX8YxK1SpUPex/
YNo7PeZS3hei0gfKklz5q784njSaxBV3sQvUry31Nmn+M6S5O8gwyqEyf6SAlXLC
J/p01XUVTx7Mdjp3PyWV7edlHGSGwXMt9f3POfxLLR6g88JGQ/L5srXpqc+73FBL
v+xxOTCOtODVgei6nExho3d1+uMJeeiUtvXsY8lB+oZpPeZA7sbmMttGsDn1944H
3cgSLyZ/AyTEsquJIqXM3FGdDvAlxeUD8oQn7+/C9XuGvSYZ6+7hhQK6eWBgxGfY
3roqzA/cApkwAErmFIvgdMKec28qfZzpxE7SMLjWYYg7FuGjdvIoc4ZJ4aUmzTr/
NpNuPCRgfojFgzel594lzOQeyFATXB0t5icC97BfoUU8htPRGlnn4Ik9UKMlU+rM
6uNrp4cHJeMhaedAY2Fnmn5j+nUIOJKJaKU/v+W6I6Zuu0okEga9fAyp/omK8J9Z
+zSoXKbBK16bEQebRKoZghrf/n3ZyyZy72pVxawo90JgP4KJAHtXuEGKRdKBJOwY
bOx34D373ICteRgRoAfDYL29YEUbAISM1y12tX2GtCinzaA9wNr4Tw1duNGnKIbz
ylAKca7C2+hl6DFwx9HQ3W2mGwXOA3FrzkAgilGiTehRKUACeFmQMwts6fymBzYw
0AcjOvYzWU6gEIGkOjUQOvYk11gxHJligqCdUZ0sbaA7mMqpmqY+iZ4sTxPbYTs4
4wpv1H1nKYoqWye7jiPjGUjLtrYToiyNHfFFVX+ixqsvDHhOewUbAXVW5GpMoJ2K
VHBtaaxgNTiG64S3Dm8SMe9uKCH9uyfQktKXC0ogEiUxoCA6coSCiXupwN9VdYt/
lAvSsPyoYYgCX9TBxIHRlOa2opyMhMctoNLod+ZtSjqEz0yCE/0gGWNshzBTqRqB
lM7UL9wbUZvtXo08tJKUkYNr/wKU6E25fOj3UhfzzPDlhFAhCqNTMszpVulYTEKW
uU8gOL0pYpaRk0RqqN94GqpvIC9Qj8irfZFh2M4jzGLGPLMi8CCWSlOsuCOzook/
Cgz+8z6pU9rQWNkFT2DMwRUYlpd9i5w61MMlB6NI57lvIBLkvc7y083K2HU4B7I8
t6LOekeZ/wHnLNngAle7mbPk57BNgTJNVkbAU0xMzrUG4nU4Y2UcRrPIKaqMZlUj
+4HQGfrTsKLByyDIGwQIRjfznDo5+kDRXuXUUqRxS6UOClncts6jw4BVavUSGnC0
8QjhmxLcgvTUoBlt3PZvJukQK2SXDx6XuVCSnz5G3zrAZwrU0Wd0nccO/NUuF45J
yUbbj8Z6yCoGrJHbLGFhKWjhniNYpzg4DK3R36EJYf9QFswhDtrXc3/pwhk29iGh
AK0v9BYkfd15zDE/ZfkdDc0xdM5h6vmQ0y7MDQps+cAvkBRdLxe817aQRPkrjnbg
7UNav14NUIizBFdD9NHUpJvrggLsz7kP2hdnKkcyy1h7zxw1K26T4pXFuGxUJ/3m
g7lacCUBP25H1J6ZJnR5N1ensBQstRs8Og3y7ONdN+KTpgjOY07KCfX/QBE1LLGK
hECeGE+lmisPTgjFe6mVT2HYoHgnXvwhPlx7Lpln9yozAzYzE5ckq8vmvNvf21DT
cBzNN5wO7bZvCCTI9zV12aYRn359ykxMjq019BNjOWmUNyipdJuT8sarjRxN2NLl
92OZPS3a39XZL3fr995EuEoVPu1a6XbHbATE3THJsr3isvW+fUUjB+J7PwZzOnKV
IjB5hbd9PgrTYwaR8aAqzaLdVq2v1kv73Zh3Q6F/ynMfy5BSe+kAT/hZCvxtYCZu
Sit+YAG8ATXq/3s/4VKFg70EsoGMSvb+gjWIx0vxl/NckQchpR8NsPrC+EdSB3CB
vU3jgrsHgjqThROsU9GvRIozwVq99AckbJKgR4TiAKT3H1l4D+ZOs4EUH49d3ODV
eOnACvrDn7cbevmsZT3u0V4lvGvS1a048io/1o6SzKHcIJeKSgHrHcDhOT56zsLG
RRQVAfr80S2baRmkdzCrFm6NYx5eP5kzBJWyRyR0D6HInL7GPJlYA9ZPSfwnqEP6
6rWxbm7UMPEEs+rXyIAwrjmLbqBaOXO8HRQ0i9rn8qwdl3V+Vao5T5enUVsU0J1H
M0unkRZdj3M54ZpxsCT5sV5JZkhPg8COdSTaY+tMWjG5QqszfIj29OtakMo/nhuS
VMq8uNFtqRe/7Y5lrGqR+IQkFDEd+D26/ZcyNPkCramc0bi2nWTvVgIoDwrnBVon
flqX33AfPh5Ljr827aio9Yqxfk5j4wn61GVZ6fw09nTE6WCrZmC8H54fpkAtUpx0
5eZvtl2nNP9l9rpF0blwW0vC8bEve2dcdMXMBIfruTSk0ewO+9YVjHPkimuDawgn
su9pytX0AMS7prFD7MpNTbZ6gOY9g70d+ttWug0z8ykiJrQVkIGSHTciEIiRDN+M
83/d8ORpMvYpPg/rQmNYlSKCjQ+mO4lD0PRiUM1/oh8DdKIDxpwNJpn27ZaXgxET
ZtgAtU8PeD1d5W79K+Mt+F5say39y3uS/RoXYV2m8twRcluuPYOn9cxuOt9awIw8
if2x89lq3EJdmRW/qGFfiyGWNR8r+3Xxrc2R413IUPZ+98i48lP2saFV8xB3gB1t
6VedSBxatS9/uZXYqvb5j3RJ52OaJHs4hFTphY9XXAEyZ2TRxBFQW6fqQJD+SdiN
ZpQIhvE8fLSV/iLYTzCrToIqG3/aOswXkQ08adTEH9sVpQtnzFeQeRW0ULQb+wGw
nQSVTuZHJrh9L7RK8/Bx9ZOpj8Bb9U3/B2iKBfiXwYfqsSeVkaAbwJgMFl4DtaUN
Dw6yIb+rNWXAhAMp8MdgauArdK1NdADNVymjcuM2XL2PK2ABj+8N6otHLvJyDAIP
2DGQwrzFFmdMTDCAL34OKiT5RfJAlj6XR0UtbXdHpnRa8lTLhziKOU/kH6OsA+VG
HxJ+7SOfZQYxFLJsfiTp1qJD7mWJZog0edSvzvibXaytoDFlenYD2YAvGxFtNd3A
sj1HZOgrLdIdgORjMb6tFSQq1ObGvnUmOiA7xRwl9HNqu3e47KK7j+AS7ZoJvCJi
2i7+ihCYa7Zg+uj0CikCsVqWv53thak14g46MoWLCUDfObBygVW/Dr31n1/6YpvH
xlnHbSXdPZZkkX309i2kcrNlfFS4/aS6KiPMNgzDw9vS9cLpLZWMFbztzOofppNG
st1fxaFrWYq/qHwOeSf951kuKtQ2q/vZlTQ2oiuWRyTHNATVFNjd/87KfsRWvFGB
dbrvLJsyIINkJw+rAQ/KOmx9thEW17UaNLLRnMrtsHcHc29Sq8G2shzV3Px56csV
4P4/dLnFzJMc1P1aWj0VGp26jsAfRe6Hr0lhYK78qWEMCmtp1iyS07U88face1Qn
aZVAra0okn4WdOnOlXayk6sXtf+4AJDPJsdaISrDOfBW/3IrKkiief4WogayypPX
lxVPhwKmenSX2uH2IoLmLlpu0pqJp6dq2KJvkRUytZlUDBWb08u1R/Ab9qT/oApE
C0vm2ZPfnObCozMJgxm5uMU/gA7oyCg9PYJkPeaDXLYy3Vospd6RuVO+ogjd5YRb
z9NZDRxY5dhY8AN5dKThB4AYsCuMu9nbS1h5oQTZNOgxxEvVXfTWvcj8v12OvJVV
Qj/RBeoK03kN5c0JFTyDQcfkBJgToNnTCm5WwbU4u1Hf/oc71fXoJ6YHSz8U6+ox
eJpIX/xMi9eMkM7AJmHd3e6FGJp3w6KlDKwDv/ENBr3baQaXXKlEzDbIG97BAOS3
/D0FE4L1Nfb/Zl9wz4nFCkEC3kzQgMXjKim+201CyWT6MxyZ4cNVmNWVVwZ3YQPm
8GwmEZdXoo9sJ9XLCygXvCLoycZRXoaMptUjvW+aOvQmkSWV+LP0ZyulV/tKc/OC
Yiu3GxSQ74MkzLPI41MVVb9VuFk5fpfF9wK6oCQ8GGm/UdP/qotQZKg6z1xeZOHI
ZVHyFkS/npkIA1TmI1P/GtPg9GkrLcxAs0IcBEqtfCOJyu0HIeBroWZkGYlbSu+x
nU7a4w5hppzKvEouH+cYa3UUcGf9ym7x4TY7KbfOLBjSneBp8+lD5YRDJJY6Gujo
f3awLUOk3upfKQCSombJJOQvAjDaVmZw4ThqWtFcAXaVZtpcZHW7HlDHY3+tGEbt
UZTG8CtVCUIL/DgNoeqsb0DvXLAncCXwbyuQ4bYpd+SwzNfrbhCPqBEmQOFyTVu8
UK6d0EPubhtBIHHv5wblJLhVwkePDdvwh8JBSLOAfrTAAd4V46v8H18EqlhlUvPh
odtyeTGUmyT1MjOQmXdn+1+63SeeU2qJd0/nNclzIkaANu828IK2y4DHTjpXMO+2
Hjf8TSmNNOpSPyCDc02vZPmJ1pI1CdzZWWUCb+oo4PMoVBDVOUyzJqc0kBv5V7PT
J6A6AU0FolbcCc17e4SFgtIDuMe+F+PLNjFhjH2ZKGHo2uCLuoEHu8Cmf+82YaX5
FozKxCepygMbIc2Lsbfp05jPfetBGDz8/p/R6XHI/1gs1rTvqWDbZwtquGFYNjpu
Il/21PZJrFU9DmipWGxMxfYzOdvbv1cVPTZYe7l1O5SEVEY9onvyodLYzR4Fqm/P
oMmr0y7WVODETwd+T1jfY0DyuF/Q0dZE2UIDq/ueOlx1ACQ9wLgKhsgzEPa+jNDJ
F+wzfz8QPKFWTDLzS9BBWnlllukNEKg/fzIxMn2FXN57HsKNyynQdPncQ6UJPIGl
Hdzbk/Hr5eGg/JTwrD2c7VtsAYR9qxZwxJegVA1kK/BmOj6JcgBvmpyWS3TU4+cO
8zhfnWcWBdlqNQCQ75VRACBANfCFd2T+wmBpC/mmcE3oktaCZwu2/k9UWtnmWCwP
eHzqYi3Rxvtswu0paLeVOEpcCVlxn+PvWnHds2wKgy8sjA59jcZxbPE3YWCFnDnd
K09OrRbby46+fwAQ0afsi2oXFSO4xdEfIGXGHgbKAXocjmGtiVPYrAmAnj3o8C9S
qMHdGEZZhXuvly/kYvdzjkNOQKJCeF1/9bxSTSg/rNwCgk2t71cbm13hOKBsQnp9
g8Zir2vdCcJRGl3hS1Ftzim7Mxnpx7CW8EBs2LsLdhEbiaMGGodewbWkLKAmWgeT
3T2Eeumrbm5/YyXYV/Y5kvuHjRcoPK+Xj+h9zHxl69CMhN0PmIUyQ79plhQdQeqI
Y0WubYY18F7NcKUF8jpgb9rXA2mQtDuXB6dwhnNweO/xBjKqWpZt7CQv50dGYsyp
foU409b3Z5A6KXI5v0EhiLODsdcapnZZxohkUMp7Ale35G4VFccOPdVJGXPtQymv
YIcMAxnPJYDdvybBFtykufeNG0HaKm4H7owx9OP7gEdSXAK6aBnHxb0YhVSHFtGa
tiPVnXbhH9NfnC/t4/eoO3CL/Y8FnpUY35lzX91/wdpqfhgk4BpgB0RZkBeQfL4U
UJpw6Xo1RNvl8CtYCmKr0flMcuMCHO1MSPo7MYOU0aeDwMulb6y8S8GyBIFgR/Lm
ECXFiszbRAsZdcZliQVHd7N1dpJbaB6kr/LS2JSfavCZsHEKI4LnM63v6VpX2vD1
qm3TA4k4zL9C3V7zGde6NENgUeyaDYzaqe2HrhTLPwzwndJZh2fKxZypm2aoeM/D
i/YT+JjbOsnlTrLn8212JQSsOnZPEo/b2h3m/6wnKJVwfJPZiOSt6MjyN9LjJ/8u
vLBLtxi2x+S/2Te5qJcN6pbxN81PZbjghG8U4tzyVpAaVeXKRP8sB9+wDmBawhi7
4s40pBFr9MqaxIkBU2Wa0J3h6WfnzZ2GjtozCel/PxEbVNBSlU5zJoikOX5cVJ4a
NSoPOZczdqEGJwIeBCYNk9rIJIVg5z8dA1bDLzpEZCHCw3ENsvZ4pGZ0gyZrrJ6k
aNR9NG3B0bDXgjDkk972l919O/3R6AEIn2jzP+10nMT/2noDpW/yY5TXDwIH+KI7
5MvJE3uSJuCDmKUvDHTDGoXGAVUuD0nx5KBg7X3moLqPttQmuuUAHKYWuxFt5etN
wGQlpMcKye6lFP2EL60+TgC06yVIdLMV654/A/bf9UsMGF1YUp/OOV541Kya7CpI
qgCsn7FfMK/mBsY+eYuKqSFlWyMDXL1e3UqL7zblOgQmeK5H86yylIJKyM8tc/+i
WB+/Qd4pguJUN7wjABqUX9Rh8waLs2c8+UAx2R9AEGekpsjYn896eH/RZkRIKxtc
JOlgnFTPdrYMmyYhWHfk8ea5Qn4IpRkKdS0sJT16CRhrzjS9u7Bn8MObnp+aNEei
e49EkXjDDqHy2TglKw5nGtB3t8Ivbwk0D63snN5LxKYcognTdbsRfZKYJRYaLc7D
oMw08/ABf+D/AiceHDnYcKwwdS7UmDynFoYz7aUkqstZBycFle2qmJ4T4v+RZjjS
EYUqmDQecQ1YhUZYoPihPav+R3whqrJptQBxwxVp6hTqk63tmhxUm8JkgYMu02fh
eN4/3HI2o2umyWDHoM7ax2AZuMNc8fQm6LvxKQW72k0xm37sc8lFB8lVi6KzPCKN
6Otj0PGwyl/5Fs4vkEG4MLSnkBj9rz7OY3l2pOZmXTG49V/wY7sciNftCaclGBb3
G+KFayRifIfNxXU1CPIdAZZNlawQqSbAkATwSs9/HNE7kra/FtejUtJvmzqQNFAb
DxHFxd3RC+1BkP7nB5rWUjruKYz4wQHeeWDvjqfe92MRzIkv05QoaLMWC9zLMjAd
nlhjX7rTzngxn898WN/lJxeowO3sc5SslB7Lol74OSJDKboWjz3ZTybLsDavUZ3y
uSnekW/bkBuLF4UF7BDOe6gYtNN1BvyRQOnXGfoxNwwqGHeHN1Br+z2rFfK9GQ2i
sgdf9/mJl8ciXhL+Q2BM2AOQKeu+k9ukgEMklNjOz1nAhoO4DiXeMAqxExvuC8CL
ccLAUXYTiHwrOAah+z1FeyMTaCnq0oVlCjo2/3Y9VYpOcLrIQaX8Gjc9IoW42hXL
fTtqXcIXvIng+ZGn8w9HAM2fB86TAY9SuHSUge5Bg/+mkQjgOUxtkys0dZyzbKo9
QZNlifRiixNZ+rpxQ+dPY7pyU+9Pf8vEgLGaDbq6h9D41HsoLeYdtcDplWbsHpjG
bqTAnGO+Q/7JEtX4I4JMg3Z8cWeU/Kq6gnBPrGKtmTfHwaU6IDB0XqwSiD4xl4+b
Nre2Bbt5KVjPKqhcBgDkdgUU+pz2yrqYKWg1ujXxS+Iq7w1yTf7tW9EPbWHUxigt
pj68p0XWAzKWxsqJb3nKX1cjVAY7+gaK46yVv9LpKqhjbxQPKudYo2DHaN+bvgXv
wafQaZPakn7ZQ3zqcVNUQvVP+073u1GWAOuc1tEJbC/K75ZuopDzF5r6GPQJO7aG
uFI7NawRC5Yzbkr36bpX55tVtSW60Gt4xiz2ON1zPOzsNt9fbbj9BhzJITdWZhgX
vAtr8z0megVFzjaP9YZy17G5+ZfIksIm4UXWDgeaf+lrLm/9N+USxGCGi160pEcX
6UcUfiR4/KBTC+bqjAba0+go6zQ6dYdyuDa7FztFtXhxsD7OiFtJB7lAV/arMCFU
TeY5v6kiyyqIB2dHUhduX6gP1zx4/Xmnvo66Wg7ZVgajrwqfpvhko1+5c+lLhnQv
5mjvhBP2VKWFIviUQrfb4c63ZLWL++2+HRsSmBoFqqwdiiudqZhJyvnjki7rrBEt
UzRCRgO+/nfYm4E891P/8HlpFWFrnC3pQw4upKrgeN4u3Lx0PUbNFpMnMPeTzShO
o0Z1vRZQ0TOzFkswGBGdN+a5DB6dLtj07+eRxPXEKkO9Fsk2fmWb/7UjFYBeZgYE
VoHqp5jvred9XS7vxX24bUjJfvjbBGMjzygX56y4Vqg6pSvzY2VdTfcgJdcw0o/3
+PR3q7iYMNYbfUtmr1BLmDygWAd+6KKdl+Z+Xb4KcDm0oolVd2JGzafswUeSdJ2v
BpswIu8lK5nGUt1j7acJdRdx+BTKBaW3DT5dQvZ9XUtVgHqMrbELrDAaB9RWLNCi
eeYVVV3z7gFGP+sQo8ynXemN3SIIp6ahg/6yfEqoRCpTIXPNqxi0jNvv1ONLvuWi
uZVSyEMNN0a+GP/8QdknKQPm+yJ/CH0+gtOM9AHqeyOq4YXuHjaCcw2VMRI6qtId
WvRS453swv/MYjnRsykddZqjT2ypGM9kI6miUaR8EcTu13dV+d2a6FcJMU3lAmcQ
0C/Lt4DiLB6+l/1r1RqL6U9CazgpVvgJR5EBwyY09OJV8VhZOWkF3TsM0+vOam6W
LZJDc2ikXvQKwBa2NmHowH0khYOOBaSn/lHhMBTqh2VqExGkvykCk2IIu0NnK+fR
rR35AfepSsCAv+a9ntSikgCqBesuCopJqb+87eprOKlPUnZZqy0dREVRDIk3VxXl
blfc/Hq1BMAjjSXu5dzbu0XNxI2L/3AgmmcEkBYSj2okFybQR51VNs+VbOyejtqJ
FEYO6cNCJntdVPt2uE71ADtDdnoZYA64Op726VEUCRgvkinoUegyQ1wM0cBg75jW
5u7MYZD0gq4LYfk7crckABmeXJxh+VWpy1eXEGkjQzmgEY2Ssyf8naTUNQL6u+XQ
UWXOYP9ADmg/rvgl9h39jDNBHNsEId4waI258QtcEju/bekqliaoAxSTvZjiHAvg
oA9bK30Ym7ecQQjR4uWlxu5vTOCMCffHIek3Fd2Q8OEM4YpmVbHoURmzXipzzX7m
fqgW8VljnXe3ErG+LZcRfU0JdruOBKuFwolFym9hLzQogGe/UzLdjpC0i0nuTDlO
CIQ+3UA/dS6Vq7AFaMTVAlyU4x2FXc31dzfLRwVYeEHfVaLUSFLfM76w/WBHe2/h
/nHD7enfblFbNA7eZXWi6Uz9/7rYeIFu71wemTrW8P9NW1mZy3ujLU1xY9X9u29A
B9nA9LtZKceqt/vcGidhVkL40PPRUaIY5IjhNkf/avyjSxnSKzhUP5lTXEjG7Kyy
2j/S1KDW0X7RIDGBdwzFnPdIsTS+LjqQH0NT5hW3xjPu1jeym6cZUXh21pmbYeve
j59TlEo50hYCCDp7PEozKHlTNTs2/Qu8t2dLNhmISjOrVbF8oGW1RzQZjOuua5PU
y204MTCUIzsfyhpezLITGje4i9lZRHxpN4hF2QBV51/+KcWKBiyH2BsQ1uhZd/vf
gQqSapAfj3h62dRwk+1JWJJ64KlkzteN6omRCKwermG9rLc9Iocw3tVS6MmksP0V
KS/g53gVyT9YERvRL79sSnjRtZsBlt2TKeno/5rt9N4jCmHV2k54+R3lAFNcA2w2
I3jHoyz1ja51Yv2QaxvY26AWIuwwH2IrmiIix0s3f0ojGg1i3UOmRVGmokhMjoM+
xw+FXDJX4zX4cYLQ82/TMK89xsNH3rBnQGW7PVzyntM2Lqt8vObH3+1LVMEglzA+
Jkmd2q8T5lR2be47tIwzjffijKGwMqIncgeOD0DV29c+dQS7Cyf5zSO83tuyDgAk
Nni7GnOy8pL/INJUfHa3Kzlgr2nDjp6r7kGgl8uDowBcr53l4u96KR9IgEtDqkuK
01UxL9ouU8TT4AP8cIE0Zr5BVJnv0VWNYdlQou1c0z+bvGEg2ZMlJBkJnLy9sPHO
UkWj9FS7PN0EhUehKpcUMogXKhuXhfav3trEjx3DuaUzMvEm2qxd5Srb/qzENryO
uoGSaMXej6/jJ33wuPpgl3187cU4dwhJMa7hvl/Ymaaz4BJMPooP1Bx+6JjRNFeF
o4vUdsk/r/zPN5+uVh5xtketvMeNgLSFwOIjGMc+HgzyO9Z42TgIMju7EOjlhjXs
l/Li0W0+2aFcsa1mtY5cQwPBAPayXwMh/e3+7CrejFfSxT65ncwGljU4vC+oANtR
TQ8hzS3EyAm+6H7x+1ZB3JfrYlVkObBE9cs97ZkXG1z/uVFtsDyHIYOgINOWs2Rn
BOydjv4vBTUYOBF1TXq7XfJMCFY8fq+f5K98PDfCpiPkSv/2cdqspr6CtOF6shfH
htJpc+bN6G04YH6ex4F6cTRGyVB5VJ1MAwvx8DsapYErx/vSEk187jyyUfQMhWqv
0iaH8JVjW+UxKqHrnKr8lS9i3ooqMfRG9WmnTWAxLTzPAxN1NUmg7D/lIiv/DTXB
E1YqXjWWlPd+fM3ZMWV2b+X9MIayKd8JbfgIHNoiUNRNKwwyiaPRDeyS7gcqsorl
fGtJzUPvwHbcnoHaypIObIldx94xmCy3vHy8od8o7fWWVhB1i+VyjYkOBAc+he7c
Tct8Frlmbn+pFFOhnORwH4F6yHzkmUqlPpyBToiWtbb8l9Vl4RiwXmCR+tZ4ghdS
cNimo3xPja/r1AzS5eK3sKxLSU1dXfE+Hx1J1uD8P2UzvoDcxUWE3YDXx+fucRhi
KuKLWT+FcdXZA5Ze5gqNs2eY76x0r8TKYaqBT31rDHbVYEJRiia3HjQg2tCgxw0f
emBFmOyozW8ljIiRKIYnLUcVlAD2X/JQhxWQD/4PCFn4gEmDv82Cn/FVai87F3Vj
P5X+a2HAL9qZf2ImXsFEa6XyOsmmafQBEYK25UA4SQKj4CtJFS06TZ/3h0MmYrab
xmc53HvO8LBLcI6GZb/d0GHDYUKnCfEkm9+ICZyF/y/rYkuD0T6cxj89Jw7128Gr
ZsYJJBfeTMNkpC4aRYVSNH+SsjszBIewKK8NAASLuX80+QtB29EwXUGeD3d96UXm
Y3iionO59ODJx0QS9WuW2Un8M2inc5JVfUiaDEqXZiRyAyz9R0MB+1DLfA5dwGEl
ZdbcHDPhA6LcHe/GJ5SNiG32t9yveeXjjdWIpVRRa34lTa/xSUb319GLfu9iylFg
P/toTd04+VjuvNX0GXPTjtUPgW6gCkKN/4qidQuX+F+1eAYrVUH24aryun7kgtsB
0MquzUfMjOoSV2z3rF9n8TFqk4eSGoTKlCHqeqH5ZVn4W3ruynHuXXLp89nRM5rH
i4PDcpAy7pQCVrn2EJh2DHgZZOZNuG1imSyUshmyoQCCTAgaqaDTHP8L7nk1BXLx
6pNWsZ4Xk769YzKvvyfbOuHTaasRrPz2WDcesotG3+HTqZsFB5XrK8mVEIPB13Y+
0V9XBFwJow9RNwvWPzIiJjayasgIiQ9VLEa5oEVeDza6tnUmpT9ikoHMOblgB52o
Q4C+i2121IJpA1u3aoF8/4czYKGXqhK+cuhylT0Z3MkQKSZPKSndfYylRo/eyPfM
s2gvDWunluL9sU8HQMjn/soN3rxaKR/RL/A41sTY+Bzqd0MuESVosAtCYDcT4K6D
Ns+wUCGySKwbDOPW9G6Pjb0neGdHbyLgxp39ee7DrPe1jr8SozHJucl2NqIGzvoM
eoXCUlsHGOfSPVBMjuqdJlZ1+9WHmungeSyZ6uSMuxc7mTfOzu5x5Dq81fflDXF2
wK5OrrIhmafcRQaWPQ2PI6TpuFYKFrYMkF303xyoreDIfk0rP/7LMXIZB0pkgEiH
h9eWH39lcpNiDwz9gLSMjKDpnRWmnsI4eaF5gg++kDlYQOX/1I+f9qs2h/6rKblq
DPL/5DRrx1VbIzC737ukAztSxj9ahUwHSp+TFqcyei5ah4z0Jw2xWRG+ktfL2l/4
X7JaH21Zt4ciudbggkMqWiGNcqcJtzviBBfV8S3g6JcaTM4aa2WmwGdgoVAK0+HE
cE0y1n7QiVwMMkAeFDonkOg/N9uduVP6ao6GtZ82ARO3WB/Y9KwyEhCD4HnonCDO
T/DO+wIeITcE5cp4HIDTSANbjZDDTx+7A2fYgItvhoQWS0/9kMMBna5vDH0MPd8z
ut8fYU98PQiReexkFzVwDilad1K+Njkk3jmwWe63Y+p9888hzOmY0R5wxwM+PmzF
lIcPyEB6icQ0taJhfs48cVQX8ApGbUxeXvl3SAP0TO0q297jsyrI4ob3yf/BXOhm
CiyYZY6Ta0QWXP0MM+7F0l7Od40WPoCPVios04/FNiG96xZe530wlKCG7oApdAhk
8NOgepB5TtIb+18zFW1QLRJEIPuCTyhTkd+onVGHtqHY9cx8YWzlH0EGgTqqZHu1
qmV3kBcsjRZB3Kx6+LmBQrGknjK9vhIXNf6TXCxlEy7ll+jB7hbi7r824TxPoLqV
wlsTQY8JMd7if/cZ6kM0IiU0SfUSxRt2julv//lAaj1J/dgRN6knJIQl5q+fCK0z
dVXp2tzg9PwmAal95j7FfOMKAHVFFunNBQeybAhHzEBVxGy/AamgtBPzAJ2KvNtv
sobmmq5SsvPTD8uDze7wsBTggMAZjNN9So3tfPMi4n4Z9EJvn41oLTN3NVmLG56u
+FrI3Ckm3q+D/WE+6+AKkqZws/ZX/DYZv+j/ITMmqRQ2Z4grx1eeIv4NKqCWpUbD
JYGfVfZwlgphND4pc0u96qFZXhdndDhKjKSlH0+hqHCjJhVamvjnTk5jNMDcYJZs
DKW7TsUPcYdMKCDFln9QvU2c3vJ3vzbCSr3Fo+6SoXLFWkTKTkzT6y38rKxVw4/y
8u1nRgqoLrlV/VERGULSKhV5J1W1fpo56iGn+0SAiiWj4AkosKv45Vf9RZ3bo2Y9
966MTTHo5i0acYpJxnOTwWigJqtKww1MGe/jrSLlw0yLlQCvN3HhZHUkM+d3f1oa
xm/TX2GNgp23zVdh9sk5oS0KoZqRZBKxVKU4nWP3jOr43pV88fA/pHGSTSkusbWe
dCx7BfrYDLCSfSHxlmy7X2TX7/TdD9odzQ7T/XXbixeY/pgZUSjlC9DeH+1HI740
7m+Iu29gu9BaH/BOrh7/5GqFflLYYO4avDXrJXNUGGPVOsKp97TpyoO4K1CywOsB
GKenZUo6faqy4IxKx1p8/3ivB1tohDgEv4dvvBuV29gDruVR0/BQrgUo9DmSEaEv
jemLNQshe5DFDIeppGpE0N8F5le4gNogKXR6LwBpQSASJLW5YnT8VirZqiQ15oOD
5lH3Eboxtv7MZTM+WHXUVuQSEEMj1+LfWKK2U9MQPICX/eYPlsCzNOsgzYJTz3r4
cxk0M+qZm/Mo1wYaEge5jrSRoFnYRjpZKFJahh1DmnLwKdLGlRJuyYrvjdFDd5za
qbV/Pk7Wg3lTpk3IGkepQnHgmeocFA8jYcqh3Pd+Q72bOMPionxqwVYIcuncEb6t
3LybgIGtiRgEcJ5bGFy83FEPzvngvOeNtohyKrQikTW7jVTuwpwEtamFWsMGaM+u
mYy4JM9nv7HYv60D2XxZkL0Q7UcmkwT3jjBqVYckcxXuFSM6jaLkwDQtc0ix8PIq
yDFHOcPU/8MVd4tBQX8K8AXxT62c7pogMONmCrlYCRz/GCnPalnK2iz6xkKgSxbK
W157OGOwoNJrMwUGHtUmFjMc6ks48GYJEZbfgRhFGAX3rwaej1MSK4RVrLTeSSAP
Er7gWzXZt2UmmQYEiI2yxWKJtySpkya+rGgiOI/5sTo9Suc4fHQwAGPo1b4c3Hdw
tE/nUZMH7MzrC73995VgKC5sFO081XIr5K8uacgDOTBQhHj333Vxxn0B8/MPgNQs
oSMbr2eXUAoZnTTwDsxAbbROfsgz1odQvaVH8x7ifSEk56LlXN65DkGrkLUYM0bb
+LbezXeK6zXrQ+AHyJuHXL0g2GxeZY6bxl2IX/maUKWgynHOrHOYrh8pK0hrE5ZB
F9AwVZbU7Umhe6WtDAjU2Aw1JoqcMabfsUNdQM5Cw0o7eLGRsCkeDXTQNYRli0wD
DjjyQxrw7wVlg5PaL3X+b3uVaEJQrq61w/86Ilg+plTM/khg5drx8gmQCTdMxnRn
PGbSEV/PND25XAoC8Src/YX4W7BlfNs+5qes4KnNVLbh1Q3luIwTnw0s2X6nXhJY
AcL27lVTfLxaLiTgZ5l10js1dB2M99cTxlISYi9kJ27z/srwPyjluqs4sdsvBAxF
EmdiTEA75e1LgA13oAdd71VHgAEkBnANRd3pbXMc2XYqLqAVTiX6OGqlNIpOvlCA
J8Btqq+kvYiL7/1I6gxupcXZY/Ky3vSUdDHeMnbI7sdD0s2Loe8nMP/quWNI5MER
miR2ACLIesVqp8mVjkCaykmIVLN+LI6v8OKNTSotROCLX2DNUzB89O+ZIuPQpFEZ
HckMZv4qNDv9PyOhuPjgYEPs6JTY7NXPx5f+asxMrS1+MzijK9BudGvjA0IPP3PL
iFdNSEniKgWPh+9XZR6RlPIWpJEBY9muPLKgTkM+FHGdM+Kb2lW6WrnxhxLGKj/+
SQnJ8OPtnTRZix2LAd3auKGA7Km/JTrJjU/BxTUwuRCHRDyLWbHjTiFIc2a1j8Hx
+vIIxfg9P0WOZ6j+LXVxsKoIkh+AhsHbpnqjB8tF/PdVn5IJhBFQ6+H4bX6cQjpb
r5la2qxwtyiTXyMMjFC/nkK5XCWIDAgIDaHZNFGygMc424QIFfcGsOhce/tn6PYG
5njOjdumJ8IcZ/eqeqmLm9XdN267nPojAd4cV9gvDgE757P9+fy+TqiC0mBXVUyg
k2ZLH3ga/spq6OE4rKG0LcBOT4bmNam7/RzzSlNLjjeCOwbLg3DOhfzq1cyO0p5p
0S8CgN75QUc7r4MO+aFJPnUO3Ad6mje2MBCOs8hLc/BNq47QZIeHks04P7psBp+3
7S97728p1S2aI2qzlRFMOSvMe8fos2mz0xwdNfVfBCBv3NRRUQfQsXAkE4S+pd1W
XyrFVvntZvL0TyUfSr9gESElSQS2kgMrkX+tKZ9RL0ZQe+D160NU16+DrNBsOiYn
BjakdvuHttQ56eVCh5EIvR32RpclontdwmrA+GVrjbrk67BjuMIkAYLK38nsI6qt
S+K8mbFSFNE5EgGr31umEPJV+wbuabed/jbpPvHb7TJi2td+a2IBwYZWet2xM7xJ
f28VbFBerdXHhWvb8ivqsUketlEb1KjOQxKG1r8wmxNyE/51ltwkqzpuoE7kRnYf
mmAWRSxiP/32G7LeMOCg257j3C15xskJ2WQFXBYK9brp/sozmDxe/obCn2M3qyVX
H/jw4MgbtBtyFgvTCzNrsoCdhZbfMP++frn1erSd2lJWxeWMJ9qB+TKAqJlLT7+P
t1VK1WQJy/yjX33iNvSVU0oZNn40KmbeqLDei/2QpnFHA+5pf6WkHkArMCJ87hXQ
WMwnJh3v8+ITDkMSnhMFxYtl7Sr/N7Kt/LoARe5riqQaONJFwECT7x18gqQqcjJE
6d2GIgut8t9gcMKNlNepkbYfeRagVi4/HgNHKUO5os2nqdBmPeN9ddByXA289a3l
gS3JBydA+vam5COfZzht0+7PV06YX7vOOo3lkHyzK8ZcwWQI4VCcmSW1gSd2Awpz
RJTecL0lNkc7u6gzTBiLhsdpMSQfYb4MdtCFU/r100+3Z2A/uKd2hhRzrymRtSDO
520SkZSoa7V8jCH4vKW206MuOHhDDzuW5mnrRtVGjr8rXanjq8EPr2uK7yri4wb6
xUPMThrIDQBMx4i7ueseATA7w8/5hIT3Lp7VSTPrsWhRiNM9OGt9NhLOTsuta9p5
0jyvmWItWwOSI420Xp52ySZ25hhUvWUjJaavcb3yNscZPMhDx7d6HKVoK7dvBKhM
NbwNtW+yzvKE5A9wP/PDG27E875Z0NGtu79Kd8JqbqAnPbB8QpMotmOx/2bFC0R3
kSfSAvxg21xOc4Rc6JrvckVAuxF0yNWqvOJE3A8EdI/71qJo6viREiwQo3SFY3Lu
r8OeOKf86+axCJultJnX5zCng/5r1PbD+xafLRoZz8kJ5bxNahqVIydijIvNUurm
Z0X/SRaeJxX3yRQKULprIwtl3MmmN/O7q+3FlDwCtd4wVXS58cvgc+YInR+Vy89U
rzYp6ZvGg3AN4GMq2WhY2RMk5nMTCr1doP/aYs/QNFH+8QooQ7EZp5PhgFKhHjd3
MLo8PV4lJRn0xMH2M61t+chfOILOFu/cpfsMoFVcfACW8HUwNSwCOpPrPBjOuf/Y
XNvU/iJvPJZzPAP0OamlnTacmj9iXS30ezTQ95nzrs5j/wx7dVlfyeonvdKe6kGf
Ib0+aJKK/M2/moG8bPUhfmj0iG74Uj85/jk7l79bkKq45u4mLgojuR4+KcXTtM+d
4k/iFNpEQ82ydog/OsTefmZHj2K5zlVzIOnyFMF1xrulxPNCSG2xARl/Su1gxZ4x
D6uX5ZdqUzSLNIKSjgFgfWbBvs8S3QNvNjFNPuxT7GSL8DHRbVuLwkGWifAWuhPW
vLYs3RWSXtv2pHsKQDGJ8O7wB0rhfVePiaGinsr7HSd6U2Hj9QqMZumUTpiMbfD3
R7/j77bljJSdy/RVeyJfLufrrpdiXVWCaXF3Z2VGA3yt3ykxls3AT1SuvySQGgFq
d3JhoRvzZFggRjygVYN1O/et7FTjtHod5YQ/KYL33rFTyWyHeSQlBNBzS5vlWhFn
ijhjG6dZsz+y2LOJsWMmHNOZX4TrsQ4R1eCbABul7vJslzSi1aFvhhKlLxsuwRLf
eavkuY9qJMn6zX0lzLdASylfjMPVNELdAYz95Hs01uVYspUF5Cv/0/PvHqJhIJtU
lzrMMwLZrj2/5V61c/aWA/F7tnHPrll9krh9Fh9I3bWOPBtHRqRVTBiqYZ+ACvJT
OWbo+Qo2b0JHkRAPEvGvoocqZ28mlxR7PFb9ulkyhYyNyICSGFLX/wv1QccJ3Noo
gLhri1AGSVnTLVm94/ap4e/Laww5VzcoMzN9X9hOtm8tjoDR50irAnOg3W8pmpLN
u+SfaQLU1tQ4qFJ40NSfAiITeUnHjN2uAD+TvqcXdIFrl/GazlbIqUsHbnXhsLYe
t4RdgjaRsK6jlu8eizSEkALLJSCaiv8/PXLw21xlvW6jfMiCXYd6yvpP3ZXNyj/u
FDgErch2LdFJt6iYteDrfuwq/fCpDxgBe8NgZiAiPthYKQtCwFhnvWIoJAWM6Xtt
wexnHXW4cWFS9f1TAPsYfyxxnzH1r0iBik0Nn8VLqy58yd1YEkAnytkVlYKiFi1b
zvmOa/JGddevh7wbffm73OHbnLhTwOt3JekANBDaIf4HRWz+c0Viidcq48EjHw4F
1n5FOU/uIQOHZZNgRj3nzB+iZ1ftm4D7vMva7GTOASnj8qVYU+pW5LqpmS/wJTV+
LkMyqb1VqNtmiPZkauav0J6EQFInsqTXfE32Ji+LM7BbgW2XcjeoL3yF/TfdQvpO
5+EboyPZzG6oEHl3UbLohHQsAgTsZXXDBOPlZaiJcVC3xoXSZi6vS6pftNuBTF6F
YfIZqFWN9TTyxhQaLtP6pJtieLjhUTXEtgEz4CNLj+S2yCBmwh9WzgGfaqi9D5Bk
E2DJK2mS50gxGkR65hPnR1ITYxSOWDwHYp/WLV2t575pvPR3dUlbeKzqwEs/W3up
JA1ifFpTUYOchjN9InegN+WD7ODqSdBF+qNMpu5wXnWnBPgQb9nnO1i+vnA8cV3N
LpAxlTfQczaMX/geYcnYc7G9OhaGwYi0jLSZYMENPQ1GTZ1UfDot7ZTBOj3ix+Gr
8U9m46Izp7lgEv9N2sNryld3R3fiVseBD7wy1c+CuZTOAgvqOCM4sZXXugBEU2BE
gVcopzTzQKTEMaduk6F5XLBkTld5Th2IHlQJ+m2BMQ+3p4ADcz1NyxvC15o5s9lj
L4srNu8jhSf1t0D41RJR9Wo7YPE3m0k2fgonYSAT87qKodm3CiePVcIeNtDtYk6s
UInCPVmXPt4eizARV1P+hmCcooaiIjmAkDsvasubnd2djSepQclWb1DvfXyR04Lz
yIVLS/6ZQv7r6QWW6OmCpp2M5Wt7z6JCAiXGY/RgGbbPRTElsjM5sLYqXXo6qzVw
PC+RGLBhEoIomJ7lfmoykSU31UzfvJrAxKfXYqCB21hlM1PXN1/Ajok0gLsRtwdX
ejQQPOgHGDx10octUh/wABPJrTcH8BiRz44xlYPUjk2VRjLZ6o8P6KS3+1D4xnhJ
ysFUYOvmr0yanFPXdIA1YAIFyNcATpm+gzy06Wo5HW1WZr6msBhiZ/MybcJnAGOd
lfb8k95252ZeT/vNOywBQduJs+8nhC78e0pfCbWxsvNoDN+qaYNOfG5hpkHxl91F
yzxrvsxzsxJzCYnYKcsxtzjIbbXrADg/pqOgTBL4PpJeWZqlmxhwjxWUSFZ/i0ws
fbgUdnue5Xuizzym5hnb5vNX6nqTdNHCQZwkg9AwedbQEp2Xn4QVDc3H6Gy+i7ts
4BjXJyH0W04DqrkVU/BMen75BSHAYg7pw6RsfyVmh2R/kzacXLINi4d/2f9lyzCQ
O8FDGuX7B5XT0rhXq0GDaUXZUDOy1hkCVOpnOrc3s/ddZ7wA6KeYu+r76v563U6Z
NbKDKCuyBv2DYIEoYHMWXfYC+L7uH53Gy8zO2wCy/BxBQE2V2jDobtWC8v0gSFRL
Rn+JsfaZQmxY/WVi/ZFPU319Z0AZZLeS+EmK4WwJ6pYCMbiBYzZMKFCpEFu6Tyf6
P/3XMBsMDqYdagIKZa1rHX+0cBsXDoekAMf1XmQ6mcK+LWx8kUiHra5HiVJHvLp/
5G79iMLWwOKrugz2IjSl6luslry2V5m2XIZQZddhmq+hYDOA9crNkE5aWhEuqUOk
k+jZ+MYZKbRyxYkUdy+gafozVquJ7DQowsxxe+SpOBBQ4uOPUJ2iesT4O70LPtMO
D+7AcLMIL7RhvdTQkfr9MPznqwmWcSyn45UWt/xWldI1INELCu991vfmO/i5ISVp
M38aXOuT4yGnyyQjyclYKoeyq+l/LM7WFx7FbsWmDpF4OipxXhJaes9B1lDP7/R6
08Xc1FYoNdvwD1eHV1oWGMtu8eYbNZKIh3cp6NSmVJyjApbpXXJ6SOMa3n0TSZhL
nfvlKoMq/T33NjO54Q3srGhqXAapjc86KtrDg5rDL8tZdlXhPYml+YjFBAczFYhP
pARxZj4X+PoiJqaoXoXMa+dyyZyIZY/Dlj/qyNtl0ZG2Ek6KYjsBneRMKhvMFrS7
GNUd11An5MUfQV7gjPf4mTeXhPrc6UR+oqjWeyyH3s33EpOOSn6dkHJlxcahW8Ke
6e2jbF7dsMnRzsTaVus+RzuTUdfMUfTKNupyGiRBA/TwikI1vJiPT2x7KYES0tzV
DKjpIb25LWBqZB38gp8VHGyrCjFBNyz0Gr6CCFpSwAfQ4wSLIQy7zOsJxFk4FFNq
b8fhhVnqnGtIrvf5rDJVq7hLwrIu1LJu0siQ+w6Yt7hFjVhbvRa+7BVEzTvj6n5U
9MWjMhyIyIG0KB67Kibg88UQlVBXxfVlJJIYj4dgDkY9FLh9x+6N91KkDPPyYx2t
nskcxdqg1Rkg9AD1DfeEfB/6+k18S7m82aXmwx7dPJDWJLKiH4T16OEPU4OYhYBY
9vjQQ8ROqY3T3ulNFFOcwNZTN4sVBdSSlO0UoyrE+pf3tQ+YnS/BPFQAagsos6Jg
N0wHI97FS1BzHg4n6642xaPcmJRu3j9TCdKfTYKOTq6hZlIFM/eudBnaJ/Uhb00p
AxrauVSFbJLREL7P8nF6+5cxDPYSpKYz6ZHO5P0aVJvaAvqX9MRC2fTL60g5b+N/
qxwrVYVWUbalYoCbxx4enS5sqQOkBRd6frvNyrpXwQToSOY3R5gMHoCJzlbfk/An
MDK1A20rKmktQH6K6q+yg1Cmmr5fyi0FDqiL5DVe6fAaiPlM39DWiM1FQo3U4P0Z
76QV0HlOE/+jKVN7ygr8CB+X4AHj0oWhKuoXq9gPFJQ9LhpuFVbscosPZvoC7pFG
os36H3jsgxu6BJ3qGtfMA4YBv3EBdnLztZzUpfgEX7IzDBvKfFHSCW2uwepPEjtF
GjxHIC2Q5klrDrIcfI7P4rOcdM/58pmBzL7qbSm8YEXOU4yuZm5hWRxFZKVXFg0y
4dBMugTG98FkKBIWLBbJUx2fAohDjCJajrtFqdrKrnJQ/85LRmnP1w4yH1dtLzpX
Rk4tb0nL0Cq4Bt9H/urreQi4iWzN7amrH+YBP+1Bb5yckj3W7yfweoDa0KTSrjl9
sb0K6VyPOmp553SL4WD/fMDS+T/50DGFkkwPzv959ZaIFONDIk2sxycuY9G1z0Ym
lMPj/kPi9BRqI4WMCq3ryAPzir+OUjt0GcDFjfyQVzWcC6gsr9AoL6O/lfEOIVYa
XvGd1XzIw7xEAmCC2w3v1K9mx2LlwPNkKY/khkLydahRACojdsau5jBu8v0+l2lV
bHMaaSY0Mh1vMAvkpg3r3bxYHFHv1ZYWCE4WhPoRuskjl3DIOd7EMZm5ocSCzt8S
GQDEIzLaUr9SXSuc+Tsy7FjTr4U1j1EWPDeMdVEBBAOejamrPtJhXRqNICBOiySq
gWIS8ahpUusw6+91bbarmvuRr7DGKjJlxUZrqi9RdIhV/9kG35+IAmpWXb0nnuT4
47JOZyaSYIBEQLFgXvEi/Hu/uexUOcqV4ApueCpWqCt/Y0/nWBXHTAnB5qVJgkvc
bp2KT0DFFdmZV7cSPgYCo68EsiMrWkIRO1Oqz+xE3LAU5/y56dRpmN5ZWSahMiHA
0+h7VBaOQm7kPbBtDwgIhyh5OK8UR0lmbeQXRiDUDUKjsk4NFP5SscdNHk6AmQy+
RzntXydncx8zEyQJPiz1tNTeb1EgYMS1zcqLDYlnK1f7EUg0Iy40bu2LQHrVm57Y
F84/Rj273bnbFOc/Q05ZLT7rneEIwwQjafMMUY42ecpLGMLMIahXwmhH2eHmZ66V
xtKYXbZ7cqxAzgMnZ83aca7oZY+zH9xRVTBMDGYIOAnCl+QnO0Zo1CzNV5viC14t
LLvHVik2uDFqF/zSglOGdVHwlYU1YALttFH5+HaXVbHoOK6cgkzRwVur6AZEWqC6
PWO2/oxUDrhMUMToEBGAqsVlnSdAneOBmt8KgdCb0KAm3eXu5DL6SVO3mJSatTBc
1ZVVptrnkhMI/LeSdSUB36avcR4cl/subZfRVTdNr6sVyIwIAQVFtQFKcAbR+sW0
KZ3jKBuKrsE+nb8VNBx7u7njoDXcVYGjMXpK82PGibZPkvo67FijocRSDg34KMs2
NDbXt92uhUYhUgYwY4YjHdQJW1cQg1m7jnAGH1/w/LrMtvhwSx+6EjUq0kKSNpU2
xLUDLMBWsTFWbFlozimyG256RCDtVux1gudbwWqNrx9/GueU0HcSbn3drDXQhzQq
LvHVp3kOZwY9BVIS5JY3O877SoO8+W0G0mclP3Nl2DwFZLuy0x73vhJiAuFFIuJV
OHoMilgsYhEIPAjRJy9qYFeWkzwR3thKXLO4Q9OR2jXMEh4whYsJ98CGddURTW1B
dvln1U8FRF0mihjDnQV9c7Ti2BqpUhG10T5RlEjSSbG3taV3P3vZjXHaBskUFdXO
IfsTgn70kYX7GNSBDRvuoXPxKqVSZUaFNnUWGDjm1eJW8/L3xc/4X7j76sipp2bx
A4KEd5X3RUDhXq7a6mY7V9+lNS8DC6ZKYCp+0qCjudR/GkM/4ilBC8J1AZxLhd5c
IpQgFvXbCZd/iKGjvasAo1VZNNhFGUPhVXJkvFRcbl3nFRokIf930x8+KEP4vLcD
aXr7iNBJlrrL4KtKy7std+enzPHGkW/uwUnJXoFmPCCnTuyif/tU8xwwy11erTP4
Ao/RZcMLbun8F0uRqUIgpplimOyld8tnxPCYdyICAyOWqIpx8kuAdM0vGOBcK++Q
rYtLEJ1pkEa0r08al/1PmKqYbtjwgLFrE4MIQh41D1RHPyWMoLpoIyHQ8bOJMYqO
nxsntrm9cd3P4pb1qhx51l6fHUprqvbTHntFp6I+bYCOJ6JQStKrvZiFiwcw5nmT
zjHUUVxNWhPUTtxlant7cKkKVoFwhe5swdDyEBQp+OqTlAEeMsxkIESdZat9GO+X
1kKno9mHZX1aXlQS0MC5f/wEK/nBb5A0kXfyVH+CODG4Ko+NJbGKvJYGZy2XOmsb
E8ljzGJb8YmGTYKz+/McELeSopR2kq/tyz0oH2P5dyrUFigift/vF3vYAfIfVbPj
sRROf50KViqUnaE21Jn9JZ6rSDEfU0m+c30Lwl6Nf//rpjv4EOsBVjTBfz43H/tc
8XdEqOJ09h3g/5b+GeeBt5XbBdrQmjZrsazT2XdU8DMJsokt0IbIc33ddmMMTI7r
VYTkKHq4xlYeKy3Ur8nZtYoUjcEgxeBcZKKYulSQhUSIprk8KBrshA3Lzs0o7dbt
jlIE5rOBMDbyPiqAzwNwM83QXbJvXFJcn3BxRpShBiRBGGlT9+cVcyJhxgbuh5Ef
TE/JmUScNnCrOLfiqh3CCQrad4nGbsSQxMOaHkWYTiywrxD34J60NWacMx/VSX/m
2Vz6HyjW8HRCxIFfo+VWRz8Fe2bS4BvxJUXoWBfx781qGw9ayAbfbYeuB2/m+11Q
lyp2fMukR9WhzoMuVGA0cnpXQVqUiSE2kDlFk8eKLOO1aSra/lANoluvlz6MzUxN
DXhHi725YQORD8KlIprr/7c5Ea/QEzMf9FxWXwkuFeWI3MxddreaX1rskxkQapx4
fXLxgRGqscEmvleQm/MrbJHVFry1O+VPikblDEKoFXhjukFtKRfgqCB4E4R0Bc24
hPj9HvpbQlaQzPrsPATQsd4kXxHcUcwON0VoxraNl5ygy/v28A4ce/jCHwIEd7Xr
jkHA0FBpZ18b4Ww4B/wnzCUQVhIxwENe9se9BfxYHBG85+FzUVYQsd30zdpv+SXK
k1SOswaANTIpHT/5r2qYrf+J6y3NaGqS/EayfmjCUhakd/cbfqiy3WS4jrM3bxeV
lVSZTMHWgRpixXpi/a5esv5nGxlgituRwyjxGfBxJ2LM+Q9gSukGMp6gavsU4DoR
8S9S0oc6/yo1zsi71RfsFsxB0sHuoJYPh0ti2K6qZylFlmtxZ8L27WewdiuaUF8V
7OL8Qjqzixn8ttpgPVvuICTA/ezgWNKn/VTgRnjd+TcQAKnv02AAvZKRapyvirUa
V6g1AiqUlJyCOfIZJp5la3MZyVABKVI/MnPuRLBPDAdlYfhcVncUmwa/PKlfhDnG
CL415Gw41/WdJ2+YuJ1Tt1nkFdKYgvbTUS8ZhlJLUk16kFzrnXb41NptXAGisTze
zpdc/GEa02aEx1vL9f2014ael1L+Wv3Z6zTqtvlKnC8KDfQfngW4Mys4y7WmJUjM
6aap2nUw+n6sCRUFKLwf0f+rvjlwhWR7At5eQbJSDsYO5xRFTwPBPbHDUe8mIWUA
aHbjY1AQGyqiF8JWq7hxh3BzEasa9VXjKusA4CdD25Xfy4vzm9Hwcp3v2dmjZ4Ck
YEG9+5e48bNsnzKLF2z5ADq2eLmTV5dkUyhN2YANYh/UzLmnWPGdnxyZcNh4dF+e
ldWbVzbMgC4sd2BYaAkepD/9F5WJF8CLHMkIwl6KmSmS6+layDQJ4CDr9cq32p/y
D6iyfwZ5O8VEyVdRftaBRSBPZuxZOpwuTIHNfpep9R2fyO/kTIVSL20K6zcoI0Lu
up6k/HIlPZQwbEF0m1OtZSJSmBY2DlEe6np8qv0V5NaBBzW7b6ldzwxET7soL7KT
46DKtACEqOYRXB+wJ6xsCgNgpXyDmtzwuVVq4Rl4iOeHmKQi77hMaFeJXmgfXIsV
kl/Ucjk5dtV4KC4UrssVXiK2IN/AWByihXSwjgwRilpWrDmTfWP8BTvAqT/876s4
1kCVHCjrl0RTV253KMaxgIJMWFt60PZX3BjkbmJ9HhcAW/Qpf6tnSGr22kWPwkzI
jRS1sYp044qd3MZjhTn4PSqjuWTR9hD9tSQ2BQ9R3RpEg9nlaoa3RROZHOA2sWYT
LjjdnNLEQo8ZqHx9OPMPZnXjZUJfcQyAOSyDm+ykLsBUt7tRbBCrzYXFa+WHx65+
/SPVJCUeB38xAmKyv5Z3FfBypX/Spn1le6034Q603yBa2Po4sOEmepDF4oBeQCYl
dTAlOn1LbBS0N1yNKJMpEpPz/oJopICwBHOdgcTrdICi+NQpkY04NsE8gHKjjJgz
RGPXYeyC32ExZ+o2vI1eIvLbFUjWKVT4YpDnJEI5Q4vLRh3Rn+4Y706AWz2We/Xo
Y3CAyrw/f3aQcnQ3cpNNixibc+bWnALWUtoXcpMixydegKuBTNwJwyt/J8TAMBGR
o8ch2kaqaIeWRkhjljKDUu5xlVERGXEDxI4d7egUSziNnxDCT2jvfWDetDhtFc2G
ECDr7C0t97Nayeq9+zUp4l365qBGn6Lp0kvxUXsZ86TvwZygch9Z4G+gJA2XHh3m
d5dAmrIUeOYeohWpATVLZ7JcZnzaBul+c0t303phUm0BG0UN8LoUT7XO1PEpHEGf
YkTHgKqA64TCkAvwj8F1gKOYg6S7sGdRSaTf5nrspkdTuNWuZTxxOx82Nlakrx2h
lT9PvSdL3uS8Cltfv/7crKNKBqeJorIK2XbfEo/XMjuIRFshHo+FuOs33dLKu5mQ
EvVLv3ptMQt6mbYL9+nljBSs/QfQCub9uP0CDSEWIjFtv+hCX5DriUtSy56+CuBM
8CG2CS0OBTn2uka9PR+rq2aasJ6F6w4E5PSylrXI590fjDvY0TplO5U3Q5bQs7ih
ErKPdFPq9K7xARNepMCw0RibKZ6JZjyHW0eI7MWcP/sEbn+JpBULyKX5UleJAcX/
EcOtNUN8J3IWZWM+REuxqz09YJXGMOb3HPngi6x2sWlZs/5aHq9+zbWykc6qdwKS
lbkDL0HxtSK1PfNjmXQkIxMkLoSzG8jinDO0Xw7iEeuSUp21APS66igSCqadkjwS
G4+bwFcPRgXlOQaRGooMTREznrwGVhXAj6MO/MswNzt4hYKL8Yt87+9IfWKI+QIy
LfyKGHSyw2gY26sLfd/wdhUZDLPirPM7SwQ+YhwCxh55e9BTxtti7FHeytiR03dd
oHEnTF4y3AhFmoWzt4A6irlIjKGjzGXcqJJAyaczsjaXIwupzzZzNBP50lkOMojO
IiwRlu7MN95XTDdoQwGFk+mg/j5DuLS5hI/i480ccsyvle4juZAmyPl4R9Ok3QBY
w1unPKz1WH6iwvXM0odHEUYP0HhTCK+mMbnrAEPk14T+CwJ9KbfXOZcWRGW/KcSD
6+DplUoBOEkcjU+QxNEtTT8oDjZF1cNQCIIYGDUx/Ia6iV92CEqbBwmJPQB+hMKy
8u5rXpmrHnVhg8/4VBlaIljcAzgpWVjEBlNegTiO5x5AfxBS0PwVrtCn2Ln8iPfP
XX2zFt70O6BKA+1oVa3Gp7tFnrpgjYL3bkFVrp45/VtlunHsodrUVtTFTbduclbD
n/dPrqze2lYWKM27sWGp9r7yDFd3Ky6V2UFb38OtXsOXqYt+4NvlHKi2X4TKBIpB
zrccXDxrMD6uHU85rXnZeAMfO1pWgGKE2qcwV0lDUgF+evxzg06xczYn75SiCnl0
LXlWakagm98Y+C1cZlfaGXkiPkyJ/rQUZvmY+bjKWVvIgWBr/RchbgVFrW6vgqXx
qtl1XwqLp/si2SvXQQauUOlBcFBI/4plmndd2vEyHl9JWQzwu6c2zcfOOJ8yzoMW
mvwaTvDy8gpd2lxZWYtitEi8HXEMlhsV96OZX+JMbwsSaWbobx+21P700WZlBpa1
zn5bxfYWpuyxNCvwZ+1lmjktZerZyKZ5sqGYoRwF+SlA+HFHQUECkaw/xzZNw5Xk
D8WieRZ/WC3ELeLwMIhPb5lB4JujmmK3fw7wJFeWI3O2qVFS7k8GaiCm3KchFCha
16INQb+wv2yKlFPjcnQPzilA1zJ4r6jmOm7L8K0ljXvQk5YpC5/g5q2fo55LOViZ
JdutlFtRRZf5nmHxaoguOKWXUqD1DmF0xowjhbdBOyqw1yqiI36N/aG7B6QLfWO+
SUKXMS0aSFkIaQfe7k2QlbJVWHhBm58KPH/LbcC6HPfUTfnBSFIKk5kpxpMV8/7R
Lq0fw9Z4APlLOR1RkXmzDxB+dtjV3Pm9jTBfqMYmb9KOARELy9/0TVC6KzUxKdHP
vb8ygrkN0B8JtDp7MOTvCmJcAveE3QRoq0Vv9r1yQR/y0vwWzcpURAlpWQTL7fxr
kCl1O0qA1qIQhdA0ua1f6mGK+wjrrjKiWqHZ+2cfQ/mQJk7dfMlW2ik7c5KNadVu
jGH9epRXwxebXRPODn3Km3JsGUqq2HDgtffdZxomKcMwS7tiazYhVxO2YWfVoT10
ohK5VKP/Er0AWI4kTQWEyJnTywpMSVKgse8yV8PDf/6z5aWhAqw18NE2TfFZem9q
wIteytpBMZ+WpaRsEGdnffvSnqY/Dh5xnT9OaR2Qil7yytJs3y9qxN7dJ2Z3Dhaf
F5Kb196qBc5fi+0MyVkX0xRln7ADHranYDIiW9cpu183VXtiP/SxyiZzlCdecpro
I6SvQprzuaXHLyIqlYEHLkIQlO4qB8wDm7y+J2Jemg6btnjkzs7n/cDN/vcuSFZf
rgwy5wQIeextdCUi2l8RLEjgiK+64X4eMgB9ISoWG5qja4hef/HosxUzQk3b+XlO
XgFjf9lObTCZCmcm0xYp9gvyHpLIRO21UXf8OUtk7Ddop92Wl+kHakfV5nJ/MGQd
x+ixiiZ0QiCwbmZ1cmhRNtu6NEwFkP+kVdEStqWNKpoSy4TuP0PBn4fkd/ZXWzwD
HEjmXfbB5z522ysiI7xTEjzfnebNlY3RY5QAUMaMVDHBqXuUA+PjHJwHyeudb3O5
5NSinCpPgo4W1IrqCOlzHDICy8IDISpkOORfEdu9Fqf77E/CYklzWPlt6wXCCxIL
wpxw4t5HBE60lDz5wyHVPfsshmDzGcTmOKufjOO8arJRqMTrwGphfq+BlG3Fzu40
gV+iNkhT7g69nLsXGOvVPHmAWb5AWVeIHBXrIyJ7Ss27EwVdCSOxtmE2GwCrgXEG
ZOtKnU+lDh8lmI6JfU6HgXQLTk0TZ+DDhkm9mBHfKP6+fz0afdxsi+EYNy2A4AcT
LcB94SZi/Zo7iztJPdrOaFks4r+A65vs7ciPDENZl+RKM/odkfjqvSJK9MLgoGGq
Wao/HH3/mDRQW/Sui+/Hg2wcGnZ6LhhtxIbtBh7q1b5LSLbHXk6z2vLLMO7rNfAz
kWDi+MHkYMdIXQQ8po4pToFZYAUHBKRSA/zsd28GeqIGkcsrlGF2hBIqQCAngOSJ
x3EorB1egIhFHk29gj/Hz1Vnar2FUJsCmNnBqgjurrV5w6RK0WUsp6rk2TcgWQP/
UZyrFOKCbDyr0MsdwUMmcNYgobT3HXiBUNnsSP3bPdA1lRso89f5/oK4/aaGKLyi
SCvX9VSZGXzpPTegPEiQ1fNWKLOYMrxF6+upwS4JpbGnwErsFuQKo/Grj6I82/vk
rgDuK+N8XyOOlf4EyElanQUk//gfyMifn6P9mrYU0h7CZSCBVNsgxpOkxgp00qrR
2dsHtQje3BK3y9aTVHjS8safZU7+uNg/SOsCrqF5t8CoUuQoZtuTAvMJYqOZhzeI
c0hGm3XgrEY2mD+mfe/3X+1Z/fpDMO2Hxemg1Bc6L1e0ARgHtoPlUyW1u7Zo9g8o
g+rhVP/STaD7ijQ6oDxya7wttiHekQrc7Z1pPwYJtb1pvUOOeqSyPIAHh9T+7Zzf
tPfORJSuI7Jxin+fzp3Je161otS3zkYpbreHRFEU0GzmqvIjYtO5BTNcmoPBMt8E
xEXb4SQoLJspV9QqNbqvrQ1xFm2e7Wmki0K/xPKu11yurlxq6hYu8GhOnnPHD04O
7H7BiV1eFhMrLplb/20JGDN6ufBotVlKyzz4OwBijU4Lr/8v7KA67bypGiMT5teB
RnyGTgxcBdoBmBfMk/MGOY1cSmfs8iCzYhM+bN/+RZuWHgOGf3uJuIQdbAAejF59
OUKrxByh79nTZKBIjQDXF5drcHObsg69f6xZNNe3dNjROnqGIn+wuoOr/yKoPv1r
tnND21j2gsNkkzuAZXhagUj48SwR+p0RXb/+wJOPLcwB4Z5GJ4Ucj+TO1fEJUyVH
H0xbfKYfwfKA3bAbSsjI4oIgyLOh0yzNNUtnXYdoeI1AojieGH1FLvQmDpUQ5VJl
NaZa3mvBagMiMqIe0llVP5U4FAz3EkfMOVPh0fUOgovVqoKNtPGqFRacxBKeSn1P
X+uqVgi+lWGdsDgl7hA8qji3K/BjdSw3/CTtqNziPZHOj+szHEOEJ09u5/iIJorL
xOnTqr+15KCQddzGSxKa9y0MJ5QYXVjqA5qQmyZxVjhUohs+7D/6Y0RRBxkJJyaj
OMeBo504K2JxnOJnUnM/n476Kybtuj+knrBoATJk42+1l5jivg74Y05wGn0Vmveg
rVsD/Hsf/hNpo1L630je9093H/0geo1lu2tZrlkMFNTw8ZbVkIvIrz7V+9DUOlug
WX+i8pRAZatE3G00+6jmRpMwG9/sfPZr8Q6GAMtUgkF96/SP63HwHbVw5xlKB3X4
WFlefes/uL58GTa9Cflq4opg7RMcaSzK7LtT0vQUSp+eXodEfUhie3XOdiSYdwJH
ZZNhfvGjGbQZ1w8YVZZbfzkusCtqO+30n/6y4o2x9u+AOXePqSbm95Pi98D6Wdfg
cPvH3PeVCJ194lUHW6FQiOa7ong+Z6xlw457t00H3JzPO6fHaoHbpFBoUVQqnix8
NrKo6Ka8T+x1Qw0Hv66aM5W6RRQf4/U2UYjLs1dg8u6z7iHy5st6BVAYXrosAMXT
i9YI9tWmvkDD9shRw49bG5RaHsG+aHs4qsU6bPfNGLItJC9khJO4bzQkoCd00c+L
b1Un1s8cjxXPx+xQI4kH7KuDwk8vqI4iRI3I0NXt79mfTYoe6DYK5TOJvba8I/Rj
iEbUeKI/JQmzNRkGO+GeKF6naJlwzRarh/si/I+7r7byk19SU3d46KgHFqTEoQv6
K4gcs8A2+VrtrRz1smVfosTy3y34p5TA4W/1rvqRYnmBU79wgMZCC2iq+gA+6l/x
2CPbYOxb01aAchI0FpqJ7jtrERvBaEU+fFspP8UwiO7s8yh/k/FhGnjkJUXxvDjH
o83OBKW8tDXtRVtDaMwFozuW5rZYcrDrxembd17DTSi7ayASB4MfYhth9w3YQGF+
wt3W/VuaGN8d4pNo/2HdyqC882n7gEJXW0m7pFwogu9bP4ulXEyTWppYyXwbJXpD
hCHU8CeTSoLOChZvniaCkniKOZRhYnWSabuLBO65mz/fr5CydeWfED7DqT8Y4Rtg
Sg6Uan8z7KC9As/g9O4B2LlNMpvZbTn1UbWZoYa/1d+071dDLWecVJCrvW4Sd5XL
rNCD02w8tp3goxmeBy8Ztzok987pUeC5q/ox8WWTfY560tovCpgIsSGcJNBvR9u9
HhTLYFHTOZa3eSGW4F9lO4RJOvktELfo2czczbp53nEL7W799+zOr22x0jyIHPab
/HCW0Jq3mNoBJsXNp0AkHzYUQdK5L/6xjJakFbyWKX1xxdUMEaSZKD6SdaKym1H6
79aO6K8VQbDbotfRWI+Y/woahzDhSjKtjfFoS+T9pBNchrjy50SDZsRptKjPiXlE
BH5Q9ihRsEFHpqFiREWE31yt4hzW0kZvip+xpFDoyBL/OJMM/iCG+jC1DLAg1iCh
/XgsqLsqP6Q8J5EaSI7aWZkDUO20tXV4Z7yPMx3FrqcNBdGJ55TtU2ZCTaNWN2gd
g9mi/v08p2h0GfcSh8I70mWU+XbMn1NzNVrIJbGOVpiDwFarmofbuWPcpBWrCl95
WW7H9lGghgFSQPQVz7f6MT+JtntEt8r3UbMTab41Jms1yoni0k33N6ShTbh/tGeg
jJ7zEJTBxIYmcggRZIpjDQVW5wcU9Kt3DkTAjMzavUAua73FgCIM9tblKoe0bQea
PPuQjgoUv64lnFNzkDrNts9NtMpCrAkeWnnuwHjk4jme6NGEFl3y7VZXo/OHmAMZ
9rsnn85ggiVdcuxvM//cofa+KnyzAcEFljinMT0sdnP1IXnW2+d7oWsQCIjnVg05
KS/NrrRYsHzvZS2UJFPqa4wULwZdbjfGlyHiL+qCU4l3BygwoEnbXsXGhATYb0GF
3zKzlistFpwiP+U9hMPC6k4I8IfMdrhLW0TQfS3QA9Sh+aaTXl5Da5vtvPFVwNex
QkVlfra1r8nGDPFjMVQlCvk9yj75aHUtNpkWGyvBjfzNcYBa1tyR/5OmlNaDpa7Q
W3q3M37VyHz+PmezwVNAVBHnOyAQ4e/dDZS42XsfZK7Qa63p/sfD9QAPOLbWfTXk
n7IYmHXUuHk50atuWsKFlWAauotM+x/+4DZ0uZTj/oQSir/Sp0UR6mp2lyol+qcM
K5YUZuts9NYF8t8BF0ZJ8MRjbasjG8lRqY8ZfuGVJqw4X6DEbhKST+bZBXCuSLPB
PZ0CUv+1MoLB+9yg80Tru4+DXYsbEqnPQM73PEp90TR96J49B5JduLqb5j0FkvIp
l7UzXox1LijrqczooKFE2HP9WExRC0P5bevi+h8wzyVOlhoC60cQdPZg0xehEloD
k42Kt1xmcuWHZsnGVIQB6E5ZAV41enLW/G6hAYJq4Qm+XH0iWeyQDjmy5yxn4Gf+
0xPHeAPfhOosXV5Ww4d9UsJZOwGtCw3G6jhvNswfgxCY90/RRDius51JYKe/J7op
aDaVxcEIGSeM4/GRQxEcnMepOj6bIb9SnJ2DWdlZOiLGvogpocQVC6QcrlGLmPUo
tSCvIWLcIFmXjx2DmWvWSbu4scthzXzfE/mMHeWM6abynP5g7j36FiFKX4jSxFJ3
wjfidL2eSkVLwWfkBO0iOZhKE3A5E298W3XRGd0/Lss5wznEvGM+JMlm1qjdGAjS
p+AN+sIKqX69JkYn2fAq+GhVBBy7D/g9FsiahgNld7OGdx1ap1g0KsBnFmtB4LQY
9v3oYWJF7Bx9Pb+ETHsukzEEpIhgP9ddMJux9/BTUFkukPqrCnaUU4DWKZGwsCvn
m2An4nhfswe7YIOka7zB/2xsCgLosZvlWH3i5lxV/nW/vdRZL2uNoZsPb7Dq7yrR
G3Jql2dqy4csq6khAUrthq+5P6VgjhFObANJ4sJr3TLt2v/SULHYuP2mkHSH5r9i
nuJtruxABjzy33tGuSWt4mu8PzbeIkqlBAwf6ybgc7WPtgI1n0/JU9g1l6KJlCQE
KvPntV+h2m2hBqZRrVjzBMS8ad2BCpAYLKfw0iwE6GAmibUWDci4m1J9Vpj+d2jm
wf04XeRSFLJ2j4sxJxowyz7/PKgJeI2CwO4gfQ8F2mhwoza1F+TQW0L3pDh8IOwW
F5t/1IKgFOA/eUehr+lgTFrriKTjL4wRHCsR5JvUrKNCTVnDP2TQs+JoW572n5d5
1LseS78Xr9JA7gcm6b7/p+mByYpDta/EtabiItjginnVRFbXkmPj5G0nYlwuJbg1
ApSvMRt5XncU6E8A2eOS4c8h/10S3xlHsRyIlX2NfSMkYJpD1hJwfg3jRswe9zPe
UDKXPsVUmFAp4aNZXjglbMPt08HgPzmyGf5abBduclJFovDa8Vv54guDO4HfkoUL
nqJH8J+maGwmJ02zjcwBZy1Z/bvvZ4l6PdU9jzN5X985BRkC1Utb9RY4aBb8Y0u7
j0WvtM3zKxK7l0x+NT2rIDD31C9GTDoXx4ecqKcHtCVA8RwahriYbT9QpS2VtM1n
cPPn32S4SDnzb/W3NRngB6glK9O0iDeACOWDTR5dhthRt7OhYrkWJq6oYHYeUfiO
DfWRV5l6N7absX/No1oVjmw6o0sx2McHD4IcxLZiM+PKtNX9NSQ8dCAk7m5Ohjwt
kzhNW1HVW5FB1I9kbFDqn05mDsuMjvln/JYzaj1JMmPEtqjo/8PClO8elSNOinj/
gPqTNxHadWd0AsvJUSjLT3lM0zyNFHe/ph8PQSjeD/uNCc6NLDGZl+FeBXMdBAYw
5ZBd0nkrfmAAYS+fKvCsbNjGvUDojzEPZb6aWEyje+uqmMtpPkfKUcHSNZoLQEQc
iUwX+H5LOX79m4TK4suiCUyBgi9xjOu+0OJ3VFibpsSkRuyjbLoRHNXsXWUX6pJ6
SPmFgsKz2BbKD8Ap2Ii0j5DRJ9X8Gmzo6yUdEO26GRWeWju9zC/PuunNa67Vk/ND
eodfpEweAjnzRgvw69WxnibUabVXhinJdXzQjLHRiPSSW7GGSNwyP+SIlguET1L8
uarebpzp40LZoOWNetb2CToKW9vrKO9I/sY7PG+FnAjf1K/Al36vEWf7c959n7gb
xNcY39dbKupf0mfdvLm+dfiWbEtDflOgj8hpK0Q01CfgOjKgC90etWo03OvlnTE+
/0LUN/v5VPkjPlbKU2h0LmA8SSOsexvjjqwiNDBxsLjfBTtdOWcM6c94GGxdJWXv
P28KmZSWvGbZNrG2wjY0i0F0SXCPaPMoSMIIs71dmZFWvKzaKfs26odwvwnRXLY0
MjY2NGJScbuc8AkFbRFAvVzK/IzKTUeSLlSTU+OTPNXUWrheas5opLAU2d0DTe9m
qEZvFAstChehwQ9ft6MCiNyjK5dB1qB2CUKLTIYczLeEfr/lTgaU2hvNI0U4h4MU
ahUIUnWlq4UsHLUTNg96cBTq29Yy19qSpP+diERwVj0TyyTj1LSraxeuHA/5GFTu
D3QCJIEQ3kEcjKUA1XiuFagg57Cfwuu24m0UcXxOxRObkcDVZ4sOdg5RCmFGHOYV
vLl/+WVK/QOlzkV6ieyWCFnSJrzmTillXxW1W/+WWDz4OYeCU4i9yjnkHLNJJDMt
5/sb3E/J94gKjRR8Kj7vx67/+MpbZRFzD+ye8LOPOgaMolKVkNOy2T7f46mQhFdz
AkUI3+d3jQi3wBJzoMGWu/ZoLX5bTPHalF3RSYprWErngFC8uoZqGQ01pPVTtlNm
K8Cz7kW+doEYlhEtFAjXZT1WB522ioE5ZykkJnJSig8ZYKg4cIJ/BiRbdEEiR9Ft
6iA6hNABlStvFS5dMIKfRlwb/TDC2Tkou8Lh1iMLXNwffLsUEQZa0HZgNZe24KZ5
pgDd2BBBLo7y2heFVajNDvTyqEZC7WXFiHXIrGNQBoLe3uUKLkYfTRCSieEGZp0I
FHyxLbUPgM742rY5D/T6CHkh6tP8UdwZ0jYoab06ychJqn1pwr3hZVdX39P+VwNR
GwwTDCXN0Uusq1PbInd1OKxWYKO0YEE/7gMF9AxURGV5PcINfkyEGKx8arVbu7c8
FCsX8p21CyROqXVsSwbzwB7/KwWYmOLLCKY0LLwPwZef/Dbf7OpfVx02z3NPy9GW
RER2EcHqYdSBr1keQVd0vvARmLPD52g+x+OnyhKbDII8/IjyrVR9FQ7BAOuwrVrj
nKDo9yQ9zWLo6RQ0magqaIoHyOTMzxNfzGhjeWLL/EW7yLjBY/iidFMuCJfTSNrk
PAQRLjSxGLev7XxZ5VDWTmWPzKbjUuyBeOU0Zc4daaRHvmj4zJ27nEByiDm+vyb+
LPHbycti3VB+SH4GgOUDCc3qUgV8RXZpp2HxB4GA0ujEYx3OeyM1xbugjIOeJ8Y1
c2QXJmHWsD++g5ALtVhAY+O31ffiL+yX97vKhfptj4clZINqnkS+Y8Bbn970uqAv
vkXGny7XdX+DhpbH7WVRgtpix37UcraKPXP1ALERRt3Me+E+Zjlh/Ed35CYajIA+
Aml3TxoNtFZDCoLsleGgtO7TmZ9vn7zSvz56NjVCOnRw47ymKmnFthAtHcwKvTC9
oEY7AblHrPlGymKBC3LnSXcUUUfp9lrH750ZYOwNv1V/KLvvrjXzlujLXfXfzEHA
Dayjsm4g/vxGAn8PcDqoHf/pDqTg7zzcyV3vV8GtoDv5mRyM7VpgnKH7gbEaW2/O
rYAwZvwqO7STr2HktDtXSR4QViUuCvjB8GSRqfBLz0Q5LVUCeyJsY/5X3BeH3erI
5X+86OS+gAxiwHjGvnE/hXwOIMsiGDXscCB3LG2g+7Gte4olrBMKBZ7gmB8CI6Kc
oRYjyXAwPRYPIRbGCU73jvWok74GTGkVriuwDlZwGGXEZZMz/IyUXjDFKDlwa9Y0
8xsXEy9b1VhaHtPB1g9KKYL6XdYidvMB/kW2Z+RJs1fjl5MUwTH3qS8MoHno5oED
Jqb8UEvuSoquVbMQ6qPquhjDPLr9gJgx7FeMaqnH2MGfmKrwGiK5xtuXvqVqUX89
NvezrYYe0dYjneH7Z3kRJsXXZrmQyOTe8hei2G1921dtt4F0ykQbc1KLeKY0m0WI
xTf1YEb6XPITAsw4l5CHU5c4ZAasHFNoA6VlB0lvrbZzBp7aXIQMHendEeq6We3F
4dFyWE1INqe9n0KpedQOjaAD0ObWT3zZCUi2jaaCC7oI2c6JW6sGP1CXbyScaRIf
FhG+t3vDBGn7gep/5bF23wEAFlPSHD4ixyHxNXWcNYHsnvLAmqGKYDC/qSa3RVft
BEpFlXwXQNYYb2G9AxFk0PZlBm+2UcBD6gLFxgdiXKIDs2pQv9bh+v8kVa0x5kMK
vc0spXwxHl3hDrod8YdxARouQd4MkJnmWAiKblCoDXxLAcx9fQ90TPzskiP7QBRE
+yM/Ue0hwdknRhnEyjfTKEjvGaMv+O0pt2Xmhv0Xr6YmiMu4eEnC1PqeDIfL++v/
BgoaqbU6q99Ym7QtfixvRcJh7nYqai2KKe2dRvDViqUorBf9yu/tXKbG3YwDnCwI
mSRY/yo1jjYuyEnbr6xcTzrF1lu2nknfSf8yh/KtIquQde9wmWUx5eyLANr/UT1U
NUwjauWaenNNKQr7oOVRIgnPBSx+ROyzypDcjDDYXjU2SAOtQZHtpjNrbIpKVkSY
4GL9Mrsbpe31Zos4PohpNm5zhJ1Rz0DNecmj6PYkDV995CMc8Wa/hoSSgPAJYnQp
d18NyKxfgUEoWXSbpSURbL2PGc/dzaMLCbyavygBUOe+qhTOWqMXPui15WK4DPt3
iCdzcWQsng/ADedF9h/LyZcpawAw6+PU0CJGhKuwwtY4Sl/hRnHCeRsnmFSyKEQn
FEOpBzh8wRMmraLhMm4guOnkccskjSpdaVD+8gUbcYYip/ELFAcdaQXf81Xzxxmi
Nz4fo9THQlr2ykQ33akdzQ7wZKLoImjbTlS2F7D6dePWpYCWmoa0fFxChicbZdOB
93W37J2nMh2fg09MmgHwkBhY0K668KFEH5Lv8V0fz6bVjftC1sWpQ7Km18x+5A/Q
DECRPI4V/EJRomTb7kQD7QW6/h6g3urh4XW88b7ajhVozqLYhU/prux3Bn2lrdLB
tJG65haTVoJuhmgDHclOt44UDr3aI71jrGiAf60MjJeAysFdS6tt+VVH+sxIWB7d
cdppR9LLFpTP7hpZQsDc1ugKSAdWNJPoK/0w/QDw9ND7/koH//0ZEnn5AUDMQXuo
8OTjSAO52P/XH2+fDxeaK+anuPD/DwK7H5cjgyP5GzV4VSt3KB5Z2CVirGD14BSa
gFEYEtCD5IENBFFYW+MClX6QyIIOaUFDFQYeg5xhPQ8sVCKuhugfCiOeKEeDbtRi
ieKMPSD4X2nvW9EtA8VLFDmZl1FRAjzzJXRWSNoDZgGi69TRSirBVq8t2ojsOS1z
J0b4tGWpSEkGwzPKRZFIJEYqUKTiNNZfLNLdXPj6BC11tuTaBFFr6Jrjcr1eJEkO
xU1bcf+K70SOpMLBIjw74awJ4XpW3FQORrUrA/h0gASZ4RapeP+lEf7W2SfHi1WT
FW/4zcWssQtgke+eNHsgyYUnMaSijVahR1Nm/9ZqBe7uZRfPMXCUVLCTmFYv8F3Q
NzVFgYpPncseeVeppb56YI1GSwj2dDklDeTRxxsNrszd5Hke0ziolMcd3gd8l73D
mSEav37OExIM7Gtov3SeZbllQryVg9XmN77v1W0MmV1Kn9XeQXz2wWen+memnvcQ
+NMj/t0rbsLz7G+c4clfo45GGq6M1d2YfNwFK+gfSLW68B3lT7xxI2kCXyaIx5VF
i1cNc3voO76vjmB2IjoBQpvxAryd+BFLJ0KSSkFUYs6md8Ug1a9cxCVMrlbYoISJ
u19merCempiqgnp8O9LLIe7KrUomhoSbOzKi+4BWtGMlFVY5FVxieoCg4cc1mRPB
MiUh8IB9SdTS8CnoXzG7vCLqT8WjT8n4qVjB4wW98XIYfOvvYiYXBoLn+kZ08O05
Qb6oxXnHx+PWWIaFpO82Ndf7QtsZqm58WF2WxvcxIuaYj2Ok66oeeIoFJhs5NqGn
tfy/FOyrt3TxHkdKAZpudfvcck95ODpDHUB5puuPMkJ39xhSHmvA9D1wT7BHUVgp
W6GmrOPurKetaYBnCAd0djIvJ0qD9MgLzp4Wb9UVFQVgDtNlMAKGBP5YNFpXKA2j
M/26QU+9ymcXZvj3DXXRXL+TsZXLBM1ArpRVeDay8WZSMrU2zQGg13xsbHbNsuCe
Odp1ulv5z88/oqQzaGgxOe2J3a8vHgP8PEhgUGzHZ10CwFdycBSjH49UVnqaoRvo
sef0nQ6mVc/U6cOOoRgRoDr5TlwY496UR/w5ywLUVfvq5sC+VpMKjGaezjGRC1Sd
2hzXoeJUB4BFV5FlrAzmfB1uNvF2yKr7S9JYiXlEVJ/CAYUKXk6lver/XOnEYkBe
7fw0yfOrFRwv1I3cRpQFZ9fs4AaeixcwR+MpINL7bCZdvHW1NITkKftO4XK8vWaJ
Q9cVUe0psFueFUGwWtsxbjYoBxdv4R0L2rZiTaAU2HS85Nc6eYUM+PZcNsps4Y1z
85QkIc9IGj9VTgZVAlpZPPPs1d7GAZAfAzhrDr9LlEFW03f+luaclfkUaKrJ0S5r
T2NNSRhPQaW/uvtavqotPU6biXBwU4cfYKiLvACz3eM70L4hnqU7MRFZm+zE/VAa
QLRABqaYzv3QNJG6OA/+A+HQmtdQ55ApWY+nJT9tZzE7ACxjjLpGaFb2irXlZmQV
cnU7NlirqqEnz+8yyEvfDUOMId2+ahZr9/N6AI1S06P7yhLD/qGrz/HQ9hhf0xDf
ZkgJiTuKLNDRmS+krU9avRuhVWKvxZmlHDV0fthcoYJaprBhpB8KaKist/hNrEFm
CAf2UfeHSLwrTxBhORQQ43MIIJcwOgCgQRSzoSGVYDBzCntgSGi9TuPQuFuwT8w1
8S6D6XqwpTjMrn7SGBxfOw7litMbMIr3+/ydBaoZyXXGxuasmsl3nutthyYiXf4Y
T+U+V4hVv9humWeAG68DQzqT2+Wf/1YnV5hgaORhcFNIUe46wH361/dEv5I/KYgH
Sw2ZRpPrH861KZ5yda3QEUvq21t0mgp/NsgUTMu98qdVQ8NAaR1VWmfv+UFkw8H1
R7VyBHvpR6W7ptDSWwUZRRJyGdUPGD/Xam+PcDjiACDY9NhHSqFM+Dwwx4lGa9ao
Lp6T8SWNSeshOTG5WucAnchj2LoGoV5iOhML2iVOC9q3VVOcdIBuB4L3Kus1sXBg
F46DhBhnhBS4u7SvE+pGfI11VnTAicm3IjDpWnwXyneSa0aricYKafvnBAZb7/Tr
i+jZhcUOgiRiyN4w9vza2lgvulBh92tsOIdybOaPlz/njzDWbuY9xVHyn2lxaso6
psqXt4XjZyvonDeijP0BHgrsebY+IKNgRGy0VWsvO8uHgpB+j+yHYGNlAT9mGeKq
a0viv13WZrgQ1IjGhNFL+MDn3gXa3v5flX/+A4y+GEZmIGC345qYAkQXye1qYb7G
JdAW4pirXF6KSX5TIS/e+ks0VOnWDOIpRne+WgSktP8FVdszKCmv7XsMulqcwgZA
8Jfu7N5uQtR5BFh+ncjCZciKtuV5ibjMTUeKTKyf/SK5h7oDskoDDpdNkD93N1tE
X5qitnh8Gw7RJTtgRYb8t9TPWruwqWSvfgwpjpnwcQGMueugJCvgzzxkP2a5C9O6
hcDh/fJv4nEC9SfH17BBkygrnBu9FoT9r7rAXIXBAIpZsEI/MR+JIEfOAHX1+Ldi
5jb7uiRVGewz0ubMfBAQ2XS9xS6Sd9BzLg+5EotJvEs0pFZnQH3s8SZX8QLjtwOE
qca0zpOS+CNMBGZQa9pjcPPGIXnNYeIqNaj/x5czw+ve64lTJQmJ2f3KjktYFJgR
Q0DTj/c7JiBxBSzB78d/D6nNqhmyMbdn+kmQYpJFcSTVH4R5OamvSVWAkrDWTakG
rDczYLat7lmBYuGj4DV2zhdz/WHMUGbtS0zbvdBAzacRH+xJE9SHA9RYPSLRqIEr
RnMeHK8GgCXO2GtMpUuxQSdHysNutyRckRHZslfFgIraSTkoUWOplLQbOhQmx6gf
QBpRrRzNvhhLWxM6+JKngv6rd8SwLyeleV0lhel7mL9D5aaHtKBPPGKnWWMjmeQY
3t+ZJpDF+i5IJsiOALRGuwDKrZlZBAnSoadc5yxRX4NeAN2lmL8585x6wcT/mATh
I6IJoBznrMP9yIsPfxyVInREiEd8e2aGsbjdRBTv7H6stF3wMlJDZWRc0WgD0hdE
k5dYy8hDKNr0IsOJO30si24FjgrY3XaQXZ5NlPSYXjrdZ50Q1zz4tXFuDh0ioj7o
MaHwEVDVHu+XggD2NECHrTcmbzX8u4d/ASXUz36X+FnhsZDQ0mzaYJUH5sYgTSLB
ZgIYKu5560RxZtAK78F+GNhAaLlmKGd+UiPZMGxTAYWWUuvUET2ikltWpg1xEaux
dy4W+j9Mfr9Zx6wl8a2uat7T2ZP29FWy9ZVZPt2vBnWa70lupCHUisnh/K/BURLs
b9sUY22CBQbVuv0FRHY5/+lHloFQ+X2Tr9Lhjcb0zOYYnROoQYVYuKiYaK9AheGR
fxkvXGzf9gSATJsonykSH4qN8m9mu8MWbBvAwGyNBt0KpYUhv4q92phwmfnXolN0
0PnMOmt06uh7lpXJKm1OEhN/EC4Vt5+dpbh/cYxCp2rBDb+GDtkJgTqccAGfVE09
8U4WIyREGZPZgomNByG/RsQ7Qxgk6xCzkh9WAe4g/9fRpLqfv8odlpNes5WG4pjD
Z8/3Asiur22xJ3R7w+TWqLXBslNlEjqm6e066iVwLS1S5t4MOjedLSVdsdNMlNpj
zYmXzPSrUGSNFjj43IbQYmSIxQuEp5YC7ECML6by4BiyBXZ6XZ4SK/aC3jSPpDYx
xOm+iL+iYXeid9Efa47zK7M1/VoLvwFgdnzI4uEiEXRxYu7FhOaL7ZhCDembO990
TO5J6epD/ZTdFxp5qHLV6fgLew0PczmjH68KldCKCY0uZ+fusKyGbbVE9pG94DVf
CVdTF+VeUlq9RKF9a6PExlZOmIXN1UT1MGhbQAq5ud5/nwxHd0wb48NXXsNI+QJJ
JcJa5DVIFjEwbvJECvIaymyA//QCQ481HhIl3+sealLgdAM9GVpgo5suHkLZ5ZNo
VXRr/mnF1XkkXXMawePUShn9eRhCKIc/jUB9YRHf5arK+gnLqaekzebmurV+loIY
k1bVLu/2snFLbRGQbEm3xhsD+8x+yYa489eIykB6Z4zs3K7Qm6EMWSPVf3CZItFp
xkEibAB0XM6pjNQIGXouZ1/tF8SbColgSQtBCZ7YPB+dYlFQLS/1m1K1uw9A/x1w
Tw1T515MuNRb/V4Xe38Ox8s8ieGHn46KwZa1SzWSaM3HMP64Vg9VyLGRqUpBUaAy
ufKxdJMrX+si4DgQM0fbKs535IIzNLvc47lEri65Tolo9UDhvU8IFehwXrUsgwjp
bqnqEp5Kt5MVgJbLc2XxVGIay9XtM5NsOdv9aS/LGLXzol/GWC6cERpQpqaV8xo4
BeOM228bPh2j2gdiof+W3an5Z3iN/MBNC5PZWNltPnDON3XuHtQupt8epdgqu2Ew
vTZdyuxgl29ZoH+hygW5OYDMpM5Yfgjd+jTG/jM9QKyWcH84EmBdhgTVR5LcB46w
9MDsIktkMRbeoTKH3bBGZQU2jmpMWJT8+naf/RGfzY2rkRapixRBCjTSlbgrt+r7
yMilnqIBIjhTQV5R+778/46C8KJlqXFcXf2348MimHLLt8rZTMXJKSfMGYWwv4N4
OpmssVTTmMluj+sVLHqHOZNCefSROAr6Lds+Clq8UAqeUqAxglqQThL6iJoFvPgC
d75rjKmUMPz4G+xeMk6+vuO/lR5qo4dKbr9UWqN+9VIW7x2BN+73jiMmpT9SzzzP
JxEMHCAWg+DE7FPjTZvjSj+UqGrEFd9UJ9FEKs7RHLQJUpWV6Aeq+ihka0G5JIuK
I/lyD1eg7427Q6Df4SPgObN50QZrvki6MoZiaG/A41qfaa/8rq+UEAnDmEQA6wAT
9QW8iacAFIdeEpqSXKOiVD0JB4DVfBAsW4FoydfA00+VrDP8e4Jko9kw3OG2DxVN
7F3aAFOVk4W37q9puOQx/5tuqnp5B1369CXyZfdzdF63YZNlfVh48rpszGo1HWUS
inXGbJQbHvgRlQvoTGzNMD5EB+K39FdevegHWQBKlPfVVtnRUQ+/C0fvjUUqe4K+
kfe5yABwMuPzT9F1hjIsnhXjJ8tfqTP2PGIkt++JlVUGFK/WgUg2pYemurIprf9z
8lTeqkAVJNmN2YxLzMhM7hyphyKrL70sqtzzVZ/pQXzPK5L3GWKfccPXmSgX+owM
abtl3molpuBejMmTHCe+pJPz54Im3TTD0l6ugZgy8/bhsY8hi7mWhd1VGkd9kT8J
Io0urATmuiHhp0dQu+z61Y5P7qoFeqyrLfKTXSgHeBGCRooy99Wn77tvvixYMU2F
A3pHcNQA/z4Arcw62PPmDO48XoRaUklUXCGCRH1d/9p74cFIA5NPLHM+5+7xOOLZ
ljblu7CO6bdkXahiXfrP7pasp1QA0PdaxluGP8dwgYpUqNhIlUyc53JUFin/HTGg
uz/RhFUDkQqv2hk4ifqQFYv5efCHW7r5JE8Y3ijcHtKCpPC/ZqdAkmKc4iEj7sMC
iXW5x2kKCMOkMbWTAFlEWa344n0JZ4wi3SsEqVFxddSFZT1yrxQ5EAUE9LTM5RiD
dZTVJRxZkmgjCFSyjff+nCIZoYaKqKM6AJe1uws5cCjcw88VpL9lgSLA2x4ohW7b
bKOFv2bw4Rc5a9dDDnvYy5IRvEi/FalS9IEVqMHwZzf0888j4vJ2ZPA2AoqjhLZw
cTwT7ggAGq2gS54yPSJTSgw+rhErcwWDZJXpvYKDCDa6T09tkvRqVLA1pMQ1H20h
cOaHoAi/rVPMmwbylyxQk6mLg81klypwNLTSaT2NX41USEJXhxrKDZXsksVOh+zS
7evIA2rTm5kqd5h1kNRewSslnuhLb+jg294WvaXsgZSgZjcmKPZ8rPMS7LNLUA+r
9sFVeGvoadqjsUtb7qOvKKHjac1QR66BBzPcx/7K4HFg2pWTq8RHUAaudCXGIvxN
FfzFZTCIWHN2Jmck1siVQFGTEMBrxRvgq4VLFU/4YEq+83o0canLjjlC+tZQvC2d
N9OWx2IZHEz/O3L8Ju1m3BfwobkTxMRks1MT4B0cMZyiAcEipMSJGjlC4Fjmv+tP
DWp8A9o5jzb1iF+KXJQ0EKyqYxSCWV0rrHN8fOrh7iHH8v8ug2ljAmDGEWkZ6yqU
TKXtxqOAqiXXMSczPNkpOlHs9cy+WfL000Bd7Gc3OCmTqdDwcuuK2fGnkWyLjrbO
oVgGrHAN1NtH7TwEOegJN64UiC7eYozVF8WnoW06Vmk2o1q5rKFRTuJQpjXWFr81
HfdSZdLS99czaTr9r1vQd137QQo5XPTZfynV2V2Ub1Ltxl+OdhOU/4EDPrP3ZRow
qeb7v8ANt7irpE7VXAnX9VCwEoTuu/bi2Ze+zoqUo5IoZF5/3Yys7GlG6bE591q0
NvkdJwZhNHvLW8FlR5u5ZwXgCnuB+ZL9pOX/Ne8FpeGb7sFyUvXy7mMIxvNQvrEj
K50SUoitHRdwkZilnAncygeYzprXzzMQJXQLDzf5e9M89YCL8/+ylW0sYshz6Q3Z
gGQhzgS7jg1SGfPv60flHbDv0ofTAUERIsA6xduTbf8zM2U+R6ljS/mQHmGPCB3u
mLAAwRfsPIkjUQEYJeSCAmtvlzbRPH/BlsKCMsh3OUpMouK6BPEG6vCGzzeXmp1J
N4BSgwrX4xviGoKI+ru3w6CeAonQoCV6xXDMgdZoUodtSLwRSJZXB2h9q1eqx2M3
GJc9rOGjqqxXOmqJ2NKafTFIcKMHOOYXlI5Vb38SouOMH5X9q05H1fPkUQw1ZWai
+i0ugaRZKW82l1zSodEv+stYHtcNapp6uQ/Eo2RucGa2qhuzGp71O0LaTJug8J2M
ogP2XKH67PEwFP/W3cqvDzBXQXnb5A1d015A0iJEQibRdw3aTmktIWTwJVv05kjQ
3MXKbHA4mt1YXNm8iPkMEkkvXmxm0gZl7WTpbAAIsAFXtum85p5DjxcP/5AlDbql
+hGgXnb86yeHtsgABEYDAaO74qT2PLUmXl3+k547x57iqTicwQc/Ef7JvNoSM1sc
SiXHPrbi19wxbJqTKryx9miMqXUMU5XWWpTvVZbO5I4zNWwXt8EAr/FwqgRYYkUa
+NyEPFgkIvCBl+xeuv9mJSh5kG/AIi9O4pU+TpPpZcNW10NHH3Pm1lcLpjAKRThC
IGtpKLMTKE8KMONj4DHo1eP8kUVzcBfx6b9P4zgF/5pxEslIOapcVRRwoXtaYpWJ
AIQe8QqcatYSZn1EPCPwnCO+4ttG6Ky/DjSSjGomysEN8Ep5I3w2JY8ZBsGI5JYg
AYxqXrL/D81CLD99at/iDm3NJP8ZLoyD5Cne+5/ECvOKleVvsOM+zgt4qIvG+8KV
diI9cgFi4hLcCg21vBsfiim5XdANa7VGcECBtXtV6cWulU7THKfOlW9R1vL1S4w7
CKoJkXoyOldjrxMmclUXKMxToiZuZ9Gi7cMG527+DpxavikrK7ZZ348Z+LX1Ui4M
k25b9A4z/luc3kcTduWlo1lMedF8KFKttIdYuEdLJwHfF9mEKsQFKuJsH/JVoUBA
PMbdBYRiO+t5n+uhx6PRTshN1yNhtLqVxhagvxr7NhIJpa2C96RaF+Qke8ZNrZr9
vvMU1iIIqa7VRpUSBZW5jXvraI1Hk1T/bySyG0CWCMEqxzMEQJiNMx18QisI72Gn
zHrK3AbcqP5dtd730SwRynVZD8rtw5Wp+4lzTec8PrfAZQDqS5EXcPRzfgQrmvvA
V2kMmGSK7RMU/q3Z/qnuljC3nzPrGUD15b2L1pcqRXRLwpznHCgIIP9XofB6nwSb
dNoTN8W0z+/TlXp8ut6piV/eIj4ONNLU2b8eu03X3FCTx3/FOW787Y/PmNV0AwES
Blgj8hq++PXtCQdHJ/5YKDueORNtX75PXYwu7SQK8otmx/xiRtWv1N6W83NeW2gE
PAwQFWDmIuS7quUDRv1cXpK/rt31xMGwBsTEMDIHO+cM7JXFuQsbvBFiOe1Sn2Xz
7z6kXQv7+gHwocZCGVc9jU0byA6VbaNcvPf1c0YxYfJ1Izhln5q9sfrXa6ifsusZ
bpE3wun7SalaqhiaYyf8V4mnR8TaxUMHurF7v/qM1Vun/f9FQF2PWRwfdry4Kvnq
RqQzp0cI4+cSgXH0QTf3rHylLabIsyMGiF+QP3njUzjG/UgxRuRsSyTvWJrNgajh
Jh3W4dGrpMgKdFZm+7u/ZzcfI+p8Niir0lxh2mwqu0/igmU6L+8JPNrirpyVIevf
oze+BdXaYvP0tT/U9ST8+d/OCymCOY3lgpaj0HVt5UN9vGSAsCdwJSZXjKf9I8Uk
7xDuxk79zbU78N3HbASermlzpFe4E4XWj/q1VZ17gwnaNjSqlPeo1M7GUJNnS0a3
uqGQxAHA37N6isucvXZBFQt1+MpRmYqWv7gHJPRyBsXV2KLj7kMzD+OQ/7I08ya2
mBZkyn04GX91JG8ap1g8FAV6Plzz5k2JaKK/87brtQws7Msl6+Ffv1ZPE8cJbUMZ
S2hPGzrM8WIrELldQu3cZdvwe5gWYxOXw5T4opTTOgVADu50IKy4ADPOyAf5hv8S
4mQSqrbhjXQ27PTFOVtJmNe9tVDsLUYJTZUd+AsG5JwPZD6dQIvFJSgyIZaHYt86
70qAb7ArIIJpJTVa1zB8sCaKurflANBvqQDfVqwPMEHYLhzl/Bn/mB39P6wdWDgM
+ml3AatU6r0f1iOPyHuM21/CxoIWnOtXnk++BghyZ3yrlHCTaDieEHiuW0jD6B8S
352XSt7riqOuEqsA6g8FB81CB1Ki0nPP9Mg9cDXScMjREE+1UaSnc9HRzRRUiF7A
I62Hts8IO+v1gQkex5DRrJjhmYy52tbNbVArEh79zvruY9PSVM2UP7FKMHIrI9VS
HK9OIkDfffzUHv1tJJhrG4SN+7MKJhIiQB9GtzPoAaqZWSipjJV7ByIK9xkOXGxm
x2Ch22o2DkEPwBRTeo6+r6mAVfhaRkJxoJSRaDko1pfJCNHrS++pK4acxPAHT8pe
lYZj27CAD1K2j3FQ6kal+bYU1/HxJpB+5XNpR0B2mDPcm3KFhpYXakU5NF9gklG6
86vpMSOuAs70y4kdLFVPjcCcCq3ymDp7YM7I424EBD2IYGVEb4WlnYJi7dzbfFHb
pghPiy9IW6EGvC9L6FFfqLqKlL40sBY2o2DBKzZdte+8imZCT3xrt/d243HoNsu9
55C/vzLxfki/ZZDMP8aP+ugxOHWQFAa03M2VFs0FK1tfVyIyYujNOGkqAqVaGHiM
iGlQFCi7/Kl7tM/0aVyHxmHJ3RsHvj5M2mIRasl5uJ670ZWo1qWSpLA87kEktz8t
uQevFNFmJtErNAX7Tpk3NYDMfQnJfcs6B5ctl+mdIUT1/08V5el35iGMh8X+6Hsi
mos2oaIC6IQTF/CXTHsWPVT2t8uPCXs2Q4EtouQshy878uNIiL/fIA+HHqRq6MWO
5mEOmM9Q39IRyw7ej+rXCiHLArAGX2tgXMiN9RmhoMmnF9v/q7IeMDnzZ7woYQo4
vThaEE//nWcWEteM1qOTxR75XBTCsJChfC9dI3F2NTrVHN/IHXexRWqvcROa3oMm
/jrbSweFDnZmAgNmHiEwniIYmRJmTnDOiKUzD23ZV2lztEHpgQ0EubXeBlXskktA
L0B5foVF7Knxqf26G4c4hsJDLYrUfTFE3Zg9VJXViuVuGt0adbys/IZv9tkwxl8n
5SVTcun/yy/nZ2gRSvP7ufiNwCJ13Uk07RVhkywwvYdCu3i8sn96ieM/faYKGb8c
AL9Kni7JGGVWuDi3NzHb1FiOK8sfPR2a/Oueg8JPKBhwe8Fn6lI305SztYEZPhPg
ytmLyyOCdiZY9sxaPYXrkwt8jmyGp34ZskOL8x7CtjN8/rHs/h2Sbw73eFIGr81z
Oxz0PGxBWwnhuaSqoV2bYU2jWDN+OaAKAIVZIZsr1V+f8lEoDia8ojh4rDXert//
eOFKXUUi7jZDeV8uXmfwWVSgCdi3yWq3Ylgr2IPQuN1KenHAegvM66w4+FOMpIPE
ryEGPbjMwWfmtXOyri/F0VxMinlPKAu6CCXVo27bbXtcMJ4LNy7H/6ci+tZOZ/nJ
dRikEZxibHV/LUIDgB+iE69yGFQ0uivjcBq1yd+tRWuFDTmzFr7XfJBxzY4wNod7
ik+ep7Ir8aZUdaqboxCrRoPUEqzpval1HLLRRu0YqemOHMS5GJCRelD+6fs11+Hs
ySS6aewCmbQ2XBgrkppYRSnFI9C2Qq/QcAXoouuppARtsERyS3YVaLqYljm1JHpS
ph31CL64tQnqTo7DLcZSydy8QwhYT2CdfW6WQMNIKcLJEQ7ojj62GXvA5Bbfs9Uo
YTWHvkJ0EeGYOqZbOPOQxoHP3KC2mJXitGEcmrtFIaM8F0oJ178gkiJrg8qyPeIY
azQyEBjG5yvMB1qsXxQ12/M2+WW9f1KXofDC3JTl5hkAgZLUWn33jpwWrWNOuQvZ
AZFsEoFitUOLO1ti+Mnb9xQ+k1LIvXS3czU8K1IaF4MYKXJe0vdLGXM0ZqH3PokY
k//4gbJPXMLRLoB6+tK/9GbLNKdcYTqWxkV6YofoFisjawnoj1pzgkXz+GEcHKFY
SbsGZy9eQe0hFspiwGgL9GPocBaCMZyCucoD55BTtvXmb+n5lD/4afMKqDF4SCtP
hI9yZvr8iovXeu8x1J6B9ttk+6iCR0rXroWSk6I5KxCep491KUk1bhOD9pTVTpPM
tphanjqJDoSW8mlbsl5koWN7OgVDB7uIcNEIlRGXwble18gl2qer2p7LjowXnNTl
2ngoOrttoGW7PGDp5RtPhclCNivX8MkEK/zh6LPsIzbCobLIgEzWFwMl/nde9vAI
lonA0YEzYxm7UJF9WHUVM7wdvo51dAtFGTlxWvo9T79KZg6CTpp7fK9ta9tWxMDR
czN/ZlJMGNGxl8yMnWYak1Us9yoJ3BVzfi0tsoBZ8IphcSnklf6JiqpwlceMVEqH
7mQuD8/J4+oKcyuzuHQsR9rdin8NIcgLss5o2RVUCmcHKuMNqbRkP1QYRkOzSRW0
gmNjAjLngS9qSqKoNYWze3fEjRUD7pfvm1h9l5oGHOwjueQL8biwJM/iy2XhL5j5
h3JnvKD4eVUxCR1Ngs3BFtNu+gYTLUDZng+tVO7Mr1NWoNr6fU+U3oBzQwyn/c5F
o/emPKziCpmAqXn30v1liAtPpdyabWV992fyciEjkeFUIIpIYhqQNz3/KxqC2Lwg
mFcuyk8j7CZ3OVMH4S24BnBpQz0IGjiY0lFSueXer4/DgC2HI2E1ERRPL6S92K+J
CxVlorsyoIxlTJ+dF5aQ61PNN1qjSNk+sm9dmCUXz8dwN/EOkOPh+ODtznvdEJ0A
lqq8t/D1yMICqCbf6oUXyqCMYAVBv2qi683XPvHS6oPyB3a8VLPGKe+KgDp1KKcR
PEQHMjuBAO1O8eMi8eAvI3mhNewPRgQewafvUyTvuEhN1p7ThBD57zSIbO1muJKS
0GalqP0AmRAa6NPnvQE9vAlFK4mKEktlYCQUUWzcZXY6LQpeP9Fh8pz49HlyJrcy
BdKh10ijztL1TCw4s5FazcYmRpSdZ/0L1yBMdwnxSf5I3RF0ZOgbTYxXgRcyacy2
CGQ9UndnYhD3Ro1tXAUwgOWrba9fUEoQHasou0D9rbSvd5VQ+Gxo8FKykwQrTgYm
u26DSAj3nIHc4/Hwab0sQ8cJ2Ug1YupyNCWKZbffn2fPfIt9eTvDOxytvTXnZH0L
CCjPTgB5+rS1gMYrf5LcXq/UOz/HJqJCt6nuG/rWtgWcpJPI9WNTWaHJ8vVtojkH
UBG4dgZjvOJH98eAO6TVClqYrnOL59bjtr0iR6YC3Fchi2jfzmCk63jqw8pXCFgo
YGg6rRjjFrzUZerFzrdEPgFS2hDnItsF9o59SbY/UNMDDkbvT3Nbyideq3cCVSz6
D3nn6rE5X96oDnhqvTIn3R5LhdoJT7hblcixvD2wlkK/vJfzkXzSsEm88F+Y3lIL
fnf0xtBsJafXudArRqHVkkcJCFe6Y0ORcrSomRO9BuA/ZYAoo3/Y2Wg/39w5nl/f
ha9gqqJ2iE5eKTlNhntY5Rr66TFD5fxMTab9JTutJtQg4bAIMF17Uy6ftyHbqy+x
JdzicEnyFtrHvm4CBbKZCmQT4HxvU/OBDcYcdXJxBaeYG8nwPRUHSKIItvSMITYB
jGJO6WTq0W3MZyqWo0L/MHG9tQ2Dgt64k9RRBqoqQX95+OcD+/C0vRzqMgBitQ4w
PYBI/ddeMnN5PolQM584DcezO4IFV1RWAhNBfqIsLCxBbrtzXbHhM2RM0vTpzoJK
xSriQEFEIF2AnRJLKCtm8Y70Hvx5+bMZ/JZ6IVpLqu0gCMXWIF55E6e49GdDndkp
gOVOvZOdAvkEsno3zdJoA8og+l6abQ8tRpaDngV+O1cYH8CyLp8k+JOBtVPO+8df
GEcX0K4SjFq+q4Qk09NBLzgmMRTyR/HB15rlmOaseFBCWLjFPXFfJJgRl+j1tt8y
lnY+Jm/z199u84DzOzFz81yP2DmKDpllUDPL/340o+HULa1MwdFxry3sC06tO9Vp
nSgAjb59upamvfuyHe9/63kJko8bRO/XYdlfp48H7p6KKFTevDZPVIqS17/RzCpE
odQ5hdspxwumPV2m+/F4rMjd0EuLeeV4ElaWP5+hGDkVpaQdc7v281TaOtoBcpse
ZtMVZB8YUhjHr94aa/NBge89w9zlaeDeL9shOC/jdQOzSvKVXHvKy1PHlBlS+nC4
25MJW/tlB8C2pBB6CHNULCMF41EUyXAc1VRsySfQgL2/SwQYs4fUFkR7zUxcwmN+
LMbSUpy3+ITvxroBjydcDIFzyKjB+DdFN/A1wKCQLKCrrDzi7xFYM4hQsktTD7o6
H8Y1sNxKlQZUhTIoiRCEPDEquwUP3g2oa4DTnoI543XZolVLwaHRwQICT1T1cYy4
BiuXOcTUN/EwWuHzcy8YCFDGAS+gZL2XeF5ztQxqK0L53jgnsuTT91kaQKKq93Ps
ZxjWS1Ee24mY486Y0yDAGMGuZdhlKRLX2F1rTbbzveyc8LQucG/a66VpDTzr+Qpy
m+BFvPd10RmGevhrLaMDVG1O50KymH8fE4ESYSjwve2CzKx5bMm6ZzXLg5krzMwz
60yuZNxEpxvKJv02hQ0NE2ZXN2xXFsaw3mXDabzrZ0XUC9v8mWOvFwtFyQynT1Qs
RVH453K6lEBZ9iZxarZbcucEva+oGIHqZEtbb01VE1QXBix0XdkTQT8QUdiIxpMj
A67YgQ/EpyF4VBzlgxCgn7jhc8xOuamlC/jNs4CVv25mh0kOt1CQJIdMCGO6gFok
q3MAbXJE0eG0p2dM3qeAE7RiV44hODqzJ09sB4o+oC1DwqYpwELcBSmO3BuchZ4E
SrZMdwuS7z+sJ+mHSuIq7G0jsIfd7uMPDrjge0spXlsTl+8+J8xh89CqXj7Z390I
zzza56uWYaoBk6RIpemMEL9txys1VrgT4yfnBi3/P905yW7FyPZonoXWXSjDjAMn
nyJgsMjWVHZZTCIlU4Ql3jaQtgtGxtvakKBRUerNYy+xcuMD7LEe+FIPo6IPiVwu
YrCYoH8g+n2RCx+hxtURQhACsAWSB+R/CdXW4gzEkeYBY1TfDKO4dg3ebmhnWEgY
ryUVp2UAsb0MhSDGGPKjjyQKZVY+KmTmr3tzgcxmz5zVqaNOL6JoBL7JWHxXNNjK
QFakWI/RusmbTms5TZqq7kvdNUd4P6jhjDN36zPp+WHcM7pQre285MaIxJbPYHAk
7NmFawnuu9K1GTmv4114d1Jc8YGhNJJq2s2rQAaVK4q6GhPk0xV28sA3FFEsLmxS
XP59P1PSjGZg+WdL2wCFQOm+QOlfd1Xhzlzqbg8fhMZV9QFOPOEvWAhfKMwIyFh5
pLtPQ96pELczcana1bRNwSfz4ufdAGWgisU0Pa1BbCnXBpB+erf86Mhj5bnAhqA5
4SAQheDF1wpXqhuAkghPT+gQcYkdO1Atw4WCLNnNq81gVfipONumG1OQ4vauHkMC
Ohlav/uXuDOhW/UOLy5cQac/3qp0LAWSbcT+c4cmJUrfLqWY0UqhmaAd55OLMi8d
zoNtqkES6E+5dPdac/2XLk5KlAAE/BY+0rLQujYpMCtfFu34ulxuUSH4ufo0fLjH
1TQODbq07dOTI6905QoxXEFz0YC0CYJAnFVdRR9JuWm6Db+pWlZCKNL4TiNpW6Qx
DHM6F1VKvbE80c9nFB1gw8+9q9G0fNlfdMawS/h1ugjcbiYZD/71H1INEBqFyN9S
bUcnT/zeRphE5XSDVWNSOqu2xjtWV+adv5ovtnK5IQp8KaOtuY9QIvFQOKwuPz8I
mHqmtwrbWTGcorf9dCgxIcbHzj7zXEMLzL2+K59NVlnnVY5j4Qwz4u1lg0EShFwG
HQ3vLmrycC0BJmdAPLz0+T7+46Lp73+5sb1GZrK+/SFit0AHNLmrVuUzXHbkv3tQ
MbK2+ReIocTRn0uEvYVlJPonSg5aamvnxxljf7j2ZXoLTQha5BLwxkOJH+HmnlS8
deKu8Du2H7OLCATotZbxqy47H7nfj2LntGRl2z1m7KHji3pCFUqpI/koxcEf0Xbg
LebWGBFlgguV57avWd+5JLkHQpTZcWETaIuraczskvQzpxJjyL4TNTdTw+12V6gf
+8VQjlY7os7Gdq2x8DNGrzYJ3ltq9IdWRkDpSrRKfB+vNG+ZJNAkI7o6Bm2SNwS1
AJWEU23HrwsZS4yPeDqb8Tv68pOHjHXuRggk+kdxwcqe+n9geWYCENBQGAjuZLKN
p75Rhv6l9PpZLzBiuSC3LY/zQEW456are+Lj7KrQpdHQnfHK2HJaT+HqX6yYIrmv
DkSXRO7ZMjEjiH3TfQdeOQLwFbTgRR3ovc9TgmQ1BJCqAFemb74MjM0u2K8auXxV
eUCXR4Mvr7znbdMRAJfDNo/1aZYchBGM/4GDlOD58A11+2ELWJLOim4ajdpuHvn4
py3/oYhau0yl5R4H158XnSBXYDtCxaRr85JfdN2tg2c7QXoHI7gmBJ6I8I2gVN7p
AAhU3H3+qPLG62cM5wpL6j1f4MNZciuWrHN6x/twVuF0TNotW0rCmaNuLkGKkyt0
IVeYcOgN3GrGI3Mea0rw/tkoFnsgKvqXm9m4samrNjeVGbqm3Ood6U1luHjjdtWK
BlFrBmgWeJSmLKKta0p3oycnZv01fFbHFa3cRMMPcUr1aZ7iLem8MDCdmXWP178B
cqiK8/UEgPVhUH4r92Db3fCQedG4vAmWq6gmWi21ThDZUBKAP9bhIS5H5gY8EsDG
JpRUGHvqBegn4z8mLpNiIjthO2hgdjI+4IXcb7PjeJeLgl2Wm0o1/jGjJMSOxIEI
s36p0/R8oj3xpvZR0eKnlCt9eKqUhtKqIihHtP9VvcomfBuvwHTOYDSOV3pObKeC
gNy3yFyGz6NE2skwEytC1vKOcY8Lx++p2mxbwjT0hxb6mS3V25mtubexbFZsIyUd
ozxktCvZ7rvkHCZnKFy104PsytXNfYs62GaKLlK8ocHIAwnglQHgW107VoF7PYP4
FeG9ziYwwM9Jd6hDyGfOUG+9RhyylP96yMUaeTCRpHbUtrHXyvxNmn3QBODyOW9v
rVnllWzf+5asdGEUgehsoUGZUsnIl+6t7Cm1lM8p4SzoPOFipBZM1mVQ4OZGcBV8
5PWDaBLuDDy6w0rUD2NN4kriVrNGSt1WrV61aqv+3uV1++H9iQnhyz5w7Otrti4S
eq3boD5by1IbIpoQjivCMfJGkkQ8oEkKvyW7eTufYzL+ls+g1FJGysjaNu7WHQSR
Iw4Mnh5ymIg6Ks/2g5Ff9oGEEGdvxy1ZuMeXciCYk+Xfr0Rpx/swx9uNClCj2u6X
LKT9xGdK00arUomQWaH93JY7kTp5rvqbYtZNx9IkV9GvDe6ZqSGDL8VtT0t53m4y
hrrJYgnvBhMhm+6W6fY0uzELV4IFskIK9gyaO7l0EScx3ICPE1q5TvfthbLnLNRi
gYHwfCT1gD9NdZlNApnQ+7Cr7PF8ElF0LPe0Ow/58gmj8N3yLAUERlooxL+ugTQG
QPqtOl+CFb5m5I9AYORPna8DO4/NLtghU0vSRwvAaBlbF5ohiNTkU6Sp6eGFNoxI
MslJvZBWTw6dT5xkSdWOSdokmkfc/VgrUKkbkqod5XoIcEg4INWDAhXeVRnPhQWF
Wtuw4JY1oQ4OJbwkEjs1nvvFErEEVA+wJwaHUsAvucdh8QM7XOmcZ13g8Nqe+e3p
n946bGsIKDdMNlKDYv5NtbhEZQ3wrPA9rCeucnE94VDAfR9/kY4kEXHjJIsUg0Rm
ChcJ9z5x0X3tTS1QznpkKWPoaNSuIAgQ4lGQStX3kcIwwTGgkw4u/WAtpbZVm3Gs
IejEBH+mgTvIiAgKyjEXlSWCVPyvSgXJQKWbTKVfZkr+hKQ/yMG2QhOY9joegVPM
8uTpuCgd3nZufJ2EWnqdYr6ujg0MRfZrrkS2k9B0er7sEKqZJ7hJQ60jxIas56Aa
CTK4PkNGspadXmtvCjmI76F52yf9/iLedFs9rbAgKFpBXK+IA/mGEz00FpdAeiMn
O6vPa7SD61BTMTp886YznXXwvbyYLKyizB2HbbfZMz4HiZ06i5eEaaiD59e6AhKB
rlXtHxqHGePAXrwmyjRhMbL59yZgOVvZO84na4NJEFNPtVl9IJGrnp0OIkuuTPIv
2+LZXcjBTh0JwWDuKyShvm9GT9is8wHjuOU31IuCV0bPeHqsHDRfdZlnJac69H0J
QE+EH7Em6f0ZeLYRAUuvKLxsTvtlwjoS2KHRmraqMegIt7s7dVSjrRlxgEGvavAC
U0Z6+tlAD6j41rcBJ7MQE++9Mwi3iTy3EI+GLsJlFKwmdFa31PlQT19Md7YNnkc3
Tp/j+27rppUvekseabMc1t2IT+pO5+DVlAQGcGxUS5oCCu4RNHmrgLDob1dkDzvU
3v185ljPw7Gmot9M111JYd/xaAcCkXR5yvaAg/UcGl6wLqjxMy5kkV56gl0STfu2
oaMWs8gy7a4G6EwqqMiVp519t5i0iexfUS7L2N2BW1wET2EvwMeI46NQ8fDHvGdi
3NU6mkxQ2yCp6uylasjL/OHQAC/+srtXnrREMtiT9xpryc+VINwyhS/9ZPViQVei
GLeOT0y2l9GPfW6TRntH9P2dVYu1LjZajjnkkssvPPVcuOn+THdIuFyEwTsE9DJu
VnxJVlTFtt/i9WRny5J26TXh6+DjJIhvGkrO+2BzvLPXNjBYGI+XJ6fTz/l/r0DG
mHfpuMjkr+xPtEmFEVeBY6RPHwcWSU1RcK4Y5vT8M2cieltZ9M66m4FZhN+CNH0F
T/Q276rG+0ryrd/IAtQy5nF0dlIm/IMJwZwXr4Zrhp7HtynFvFPNNuYJaxvPDt6h
DzEtE5bs1PQ8fhYeqybbuMr9FkWOTXZjMOoKI4C2VtqHn8yHCU3yjVVpmkNy4mjZ
ffZLoj3893pHsHqzVQdSo6/tcmURgv8T9ddPILK6itaS3OjF4t1sQ+1cxWnjmln2
YmAtGj8/Id82xDQ17ov42X5r+MkxwFbhdFmtDtxmR7KS5Ntsq3wwXq+9o4iXwZDM
VMQpvkN9wo9qobXIuF9+hlPFzonL/itcjBTq4qIMMjTjCvyv/NB0XAhMMZssn6z8
AT6G/mhUKb/OwsL9p1SuHbsZT5DNe7bHuulCbSoNdf8qc2gdjz2uddPEO7vnj1tq
3wN4MpZRwBiX6q6CJ+lPzNr++eOKqcuVeoc9HGiH1/lo4EXU4/yTNOXd3K88aXVT
YkiaNiOaARD+Ktr3+j4jzAJAiQpVP8CgGuqjfjiRyJxfaVjLRzuP7+ToB/TTJlmt
o0QBBdLZ6lLW8/H7/gQ1ILNABEQKQYRLkVrnvKdBinghxNg4LK4VBH8H+RmyoVkL
RnVPcNevFUs8XI5T9BeT9NcHU74NvRCfV7aFYKc7O9QhRBQ918KhQKgq55MFxif9
1RPsS2uSrJQUbOF9K+h8SxnrppE2DrY4ehnAyVyAF+YJwcy1DJU0EhKfC2iApheQ
ItMZviOaMeXXKRxwPqaPwW4d2wg44ZlwuWFM4zUkMeBn5qIBn+ErSN/sCUjwXO5K
qjdwKHcbC9m7h/97bLO4umxcP8ScZD31a0f7DPb6ShgeEOaP7A9K7lHtR+e4926X
eTUJg1gfaBj+3yoWIf/TPlWsoP9rn/dNMRSN3c9+70oGXpoN9t72GLLlTymUiI5t
MPcgmuaFtfDOT8wwG3dX2u7YguATwSV2BsbmY7ihguD7p4aDtKhoR81CH4hDJE6E
/EaeOq+pvBeLTZ+E9m+K2q+TvELuXR6Uj3fdlYLABtAqc6qkzP5tfVVUAmcrVrTH
YuKsKxfINi1xBarHkPS8nAKLIw5ykvqKQd2WQ6G+2av+U7ksY0PfxFl3OyrIL+mR
lt9RQ4iM39evpyj4FzvRvLgw2H3bxdHRrYf+yVnkW5M8D9RwQK/3mlOHnl76O5X/
s0HOzb8S2Mjw/vewNUkTIAS5b5nDUbfQLB8V6kzIrAtvwlsKzdKY6mJTYywwnio+
44ZZF5cyWncC0uVQyj1Quc46EC3RsehX4sXXRLX/c7n3VdHycamaRNehOoeQpGoU
cBdaO4UNhWgetfUblsNAJLCIdchThZnjqCy9QNR7pRR6gZeFpljDap1VGaNbBn09
6Pc/4yysyaKTz8nOqoDMSEn0ooCDIuU6Wn/9M73mqr2FBsZJ5gu2v3lqYZwN/Lyw
KvG0KhEFpCugjq76jMqa55VYvlf4G2nYRBhno8C7dwFHKM+ry7zn2dJ2p13I/wVu
n8ywOlLolh9kylPLsL5Wk0AD/wuEE98d527dzaTWijWMbqGTvKDVvnCYVFwIHKDP
5tuhSR+jbvdpYw2/kEgUPe1g0z/kMbZtZaQKkXOlZQG5BXUf9lGVQvkO0H4uPcjI
569sylvR7ofuFSzWdA428v/OFDT/k9+lG3mtCLETjdxlUF7NuoswQh6v65nVn24F
NDIA3uGufKcvG1hv6Abt2P9mpSsvfd7thWoH9RX9Y3WYssJRPsrwEcVfAXyNKtb5
aUsPaV2pUiM4qaz6mHse+A8omNAgwrODWwiCCpumUSsqHJbTf9rDlOFxGny7IvY4
6nWhaufI06YWRWAQxgwsZfU/T33jZ79H9PNKLZzucooFkf+NJ26E9cIH0axgtb7W
kqXOGMaToA2tYrpX2F9qs9tih1WreopCFsGv8yQ9aTp0t8kqu6250RL/JXfKMVTp
WRnEFdWxcAfbeNb+QpqysT+/4h1vmzkl1CA2b1tXhLD3f0ILwWshQPSkSd1bcf/R
x4FLPKEtxaJUCeUv3Np/xQJ2XD+Me9YjqadnAvLpGWLO3/bTalv8UXoolPTOyGza
dRD6TnmzmBOxsTXmqp+HRnIWMMjnps5949MyuhV16ZlRJWW6VqB+rAQO7KbbN10p
4c7xlLH3ZBAPIM7v36SVse9EO8AozpOQvjKpJX6nvoPowAZPJOpoA7xQxtdIYwq0
Ps0niVPXqqNBx5xPVmuO3uj0pNsMHUwriS4LwqB0AtZzZt4VoRBevEGrVosrVSiW
efDoCm1IQ3wsFOkP3BtGiiHysirvWFLEFkmvbkzKX+cDkuYXtVISiQQqiq1H+ld4
REVLiND5dMfqXuD9WnAFiVfDUwNmOQ+nQaJqpNS1LVt2P8EEqNjcG8yT3LiDOQ7I
9EgGxe3tNSFolWx4dtuyaD5il8+pfhRI29qWwR5v99G5u2e95hMDihTGhYga+BZs
vAiJ9Dqr4AARRfGTV1QyZPW5i6ntecL+aqvd6ozv1pbYiNRBYLAya4Tp+dHIaWUf
MeIUBdYv1uG7BLGiBC7sEEV2iXHTt+6gEGUhSRMsLjzmkDEQqnFrrcVf+7+T/uR8
yLWC0WMqwfqZ24/iH8G5dVSYXjtlLtdHZURUoSy+lWfub4EV2nC6a7qLWwDuynWZ
jSNDYNiglGNM9cFJFTykJUilaA5CcEUdlThXRSSZp2M7ch0LJ4uSYGjB855IHgiF
5mvhtfW0FxDeL8ynhPl9ki4MXtHZGJ0V913Rc0NI6G2BtD6O3ZYzP8hrL+E99z33
qUMJYLPU0Ic3ziiHy5ymXvd9Tx7Sgr426cU49TLWoXR7isDSD17IX68Qr3cktLi1
6W6Q8BNixhAh+2bhClyLbvaWmWySqLB1ljk/BfriNvynIjioIc/Qyf8BBIdWd3lE
QLS4qX1dWqEV8aQ/BL9sUPCch8EYC+SC/ngvFJEF8tmvSC6btOgUPQtET0i3qGjW
nqI/I3vt+j6qkw2QpWCp5hHLUKmaUs6KwBMy3DlRWusmxNvnvjFH1GGBZyzva8P6
VoPpViENsLrbikNgJ6yakHpSvDWXWp1DZAg6m007ON4C0c8G0O5q0AVw3VXabyzR
rwGkrJi6vX62TNncxH5uMU//HoVAvMpOvThmHOUpXkC/GeSrek7jgpE2WP5ycKaW
nSAWdobMuQ3YgA4D8ky8mHSCyV9aZF+hrrI6xuaBTnu5KzYGFzCm8wqCaqVuFNk3
xLShw2KXbaSkhJL2cN2pDh/KF3I0KJnYiYezj/HxKt9GHLKjW96+jarZLWGtg6SP
GiQu63vpBd8Nur6+vAVWIllHVaiojmdyaGe01OkR5XCNkmNVwJMR20S8SnmN21qc
w1OhwgskXJRaMWb+yJV08kvkfafqYuUp1JJ0ULk8/Qr8bd9/HDMmrJFvtqOxLjUO
wRdGZEy3DiPCn7xtRkARBZul7xXpnkQZW/XvaEWaUhFY538eAVXdBJNfKTDLypZx
AHCU+KRVRbHkGAtvT+i5z6LSqLaHBk9O5DbnYfcEGCC0McD6FtLfY/h/7XxkRrWg
lAaqciRZUb1ys9T4gl4MGsSK+UV//6hxZMLJMcrbT3eLvjH1ny5qme3Ak4ReX6Xr
kfezvbENBAEriaW9HumxqgNV2MfTm8/AqJPTbAIZZXNmaOsRUOvzaejvLoe++7bH
+gKDOYzJtL6q9FX1UUBDNSrGcODpRwj+bqH/s6IqR3cc/DSG+pgy6rWiKxvNw6Vn
4eDnVbprKMEC5MUy6U09r6xfCEPvyAcVTnWebOFDYpuKkW58+1RqipnpLkxubv7c
NfZS4MxKbC59C0le3+2g9Il2+r1J9XpijK509zKfy7CgYwpY5nkRGwbTmAkfS/wx
rsLWlQd3YOQkbRUcN2GW+7mdMFT2KFKa18A3bmmbWaepmGTNgDG3ufgimgpCGdq7
oksAXCJaPNEIzwmBAU03oEwzeEn72Z6Ang9sJWydvk6bWedyLzDCCScZvL4E6W65
mPp6BJBwHrNir1uMl3cg57TPOYXDVNYHIcVBCNo+zto23N0kT1xr3UHA8Iw3tret
6KvAOU6cQBCyzFgNIoQxodrbM4+YcYeMr5iEtsEk94EvPrD9ow5zA0Jf/qlvy/P8
+/OeUhtLnrK/hVsKHchbNmwysLSDSD31WpJ5Ra9IbIiGo5Z18lBjZfuleBT1p7Rh
L5wdM/15SOc4YBmEcJk8NGHyhU2yHFrq6ZBzj0GUDGyiHq7v6kM6fFiL94oba2Zd
LxjmRETJal4gEtafihSLwQvpiTUh1tcy9M6CW09Y0h/fE3luQU7elfMJdXpQ+icd
cU08VYmiU6/t3F94e0ad6S1nPj/nQZwAHnFob7Pym63IaXUVzjS/CAhDjaQA8JBj
yX1xzbPjbBjy3VcTdYBMHTIgwCqaoQ+RWnMyrBUrfqUvqd7P49XvSh94DBMD/UoN
pTuh2WL0+FDOlkcixMW1j48agU7jnsMaOHoBKhl9OZ4+ma5H/qUvZP+fbpkacPbU
8gVzbj9dcNXH36zmlSwp3104sgw3pE7f7kk/hCksUMwGF6vf+oGLDS90ZapICQaC
8ZWrUSW2Aik9zhpIlcLAtlRkaKDEjp2jniREajO6e1143PIZkDldPMhdOlzfcZXs
u2rpZ7FCJdTw68GjLwGmelVaTVGAI26pqKOXtHbFc8aQ5eyAou8wpNfNo+PZbIFB
sSERTUekuE0MHcY+Xv52f41vYQ5DhDTRhAhlSxNQVKbYcTgWugWazNyjn9Tvn8Qz
I0k4o6to+zpT43KzQMc6uP/pDsOB3t/FsdX92/bTX3Ne8PQIVnpS5raDo/C0XegJ
f+ZdalsD6ZibElY7d/F6+e9AaWHsy7xKmRyHqolAkkb3gV4kUz3NvsciYL1p67Xb
4FkF2mtR08EiU/tLdoMMJo94qcpSNQx2RCxuQlVpPSCAU6mgG9XkdJx3Ky7ntVHI
kyK/6xc83pNL4xWCzPujUgWs2xFyMu6DGmJnlISajxhlYFCtf6kSGGfcsf6x1w/e
g0/IgVgcOtrt0mqlvG18dWysk+IF8D/jmy3jrG/yyXETV0yhq+YpaohkDSLrSBz8
k5IQhb3CIajwPZPOQbpRq39+v4nSSMn1E6UUSWP7RkBkLKY2sy9JGcFqzZMdVr+8
p8k5/W7648MBpnICvNzLCZGApQtEPE20uA3Baf4oDzFLgHeS2ETqWFUYtPMTGhSZ
B5yfNm+C1htKZPwhvPdhOPVp5PDvQRpEDMEI6zI66g8dTZZ5bVhYLi3ye5j6QQVb
QoxWxiM6ALwcW4t7HyhBNIgrthdIaG13Stydsns16WyeOBkzaVjqbxmgO51Bbzqo
yhqJmu5mNJslty5lMxlrWAhNrEUrHsCz8CWREDj6ycsyiBiR859r717W6WJfs3Ju
sN8sSKH9zskO9MxXjmdOCATXiX7P72uOuEwn6z46qNMv0yNovsCKb9Wtsq1SPY3y
GjjcUol/afhYEw1ZKGumlkOuL0S+uiVqUEHbGr0R/bPYB3P6Hf60A6zarEa6SfCw
hlogJ59Su2aHcYxX6vBEFeTK556v5CdCDeufcik7Hv8uhmghnDqDi2sXw4oQr1aP
dBN2bJkly1S/Z3Dv2f6OqE13sPKayumcZaitRMyM9a6Hxgj5tzG7gHa4XSQCZUi5
GGWOBg9rCZ2SBcn8qwYmWrNhwZfZDsRRtOZSHiVuAkAhcMSm2X/olH097eQTZNAr
2/1ujYZQwLYJuUEhUKdrb1auGSIAXZ2GLBgOLYtubCsxNpRLfqO9tlpq6YlxJNdP
e5vTzdzbzY1T+UTBQxWBd44kiO3qtWkr9TDMDvGJAgquAz1y485m+UcGR72yqXN5
tTtOHmJul030gspk2zV1GJ+H3/rablO8j1DquieCLOfzSFS+QEJeTnLuGdB1Bm2J
dAjMOfQsxlyXGMRSHb69XkZDeKn4D4qIa8ZY2wRYD2tcAK5TiFIuJX7OH8qsM4Uy
Xd+b1OBJzVwMa4UHWCyR9xFHNy2+4WdEru+VrC3FidLcIsON68gxJwNRA5MHCSrN
x6lPDqqD0V+bqBVsNbV9b9/G8zDleCcBJuydVKIE7ld2Yg/CF3wf8Wjm/hssxqbt
zS9h6+3e+MN319hKdgVwMIw5lnSWemI3Ccq9Ivjy/e7O/pp9vUx8d8xHsW1q6OUq
lEbu6trXi3TEqOoLlNrlz/Ug3eFt1TI+WTWfLuGjGI69IwV4W+PAbWFLqkV2zshH
wX53OeLGVKAzBt90TUfxAYSRIFbqZ275JvZNuk52dbWw5kMo4NRnq64/qBAihxI3
J7XMw5pWIxoWtfCV6Kza91d9Tq8j3CAIZmiMwRQSGDlvrGGn8rE9PJDmRTVD2kPd
T8rXSWdVatQeaFT8+h0AD2jx3IpmeMt2sgORqkPjWApb2MgkacT5MwXbLQSavLdt
34PuUOj5bfJ1nkCWGI3PLlSxkyLQ1dKVqrYijFoHLLk2VwDMvfxGW5BnRikWfyAu
8GBMPBvHIr5MrQri06dVVVVEyBsKi1amzLZ1tdjR7W2JX5JZXx6+WZPM+FLgl+5u
7z6L0uUhBxADACygM2EKZYfmm1kRuVvPmRwclVM4B7euo3LVBbzcoSv6zfA5t/dV
CyVldgpqIiFUI0NVMTi5AwkyHRuSrGNgczj06LpwCQlNOnBtc7QePTmyeNynmm+T
per8fiUM9EAR9DkoIeJdBztbawqw+iIXH3AttRuZflJd1H3PXSG33jP7QWcSrmsZ
CRWsIt/lwBtTtosW7hgJOqckZsa6UZPDoje+ZKNsVVT0lzttbzAlFPdfEcn77r9u
bIYT8Kibhd+ztj2mMC0AGOWOBGcDqDkERAhDTgXzv+1/+Kufj9vqBm0tsqgpwIp8
rcDUtQSh1y2L3+qjCjwujAx3v82uzhWISzVVQ2Lwnf6ALLy1DeAu7hrJKwCeB1YO
rDMBO/uBKlIEyZoIoMPNih3nTLoSP7rkYZe9earclX+3dzshx394WzZnKzUfhvvq
QdS6IiYzJJibYhWhONtjb2V2dtsE7+n1dw74g/tkCad08IRMe0tp2hQlHfvPl2Kk
Aq0EDX00FS0j69PVkFJ+FHSkVZ5S1UtaCNqWusI0qzxbOlQPrEifcqIFw+pFTgSS
aC0UGojbrWmt/37BZMq6KRi+i6c5HwW45/3+PtTRtyUj7WA4HyLVaWACPI5UPMwQ
vwrEcRBpKb+z8R7N4G37ruR2TE4vaRSb6UCve+GJLyapGAlGawpdRF5XLmIho5rc
VulBHZ7EiRGOoTCFzI3XHVtuFx6gPafboObbodrQ76LzoFS95LIDM/EE8TVXdFX4
A2nCVxZuDJMYg2GGHh6n77TQiNcMRoiiFCqGGbFKwFeu0VAv2A4dNP8auQpCnQP+
Kfj8r0JR1wQwkcqcO5Olm3mQm6nhlkgMERTiG85NQol/OfWVk+rHfFgNflBJHJZI
7zaErfTMxh8Ghw0NooZEKpkF1R/bEC5RVE9ay69DPuaWKxovf5bQXdYtQNiF5euT
gQDuUotTZ+8mcVkf/TIUennkLW4f9mIpk1QJo1lQQh5b1P4UFlUbUQj6PbqFuyK5
kVLQ/LxqmXVCDZginHXjXxh7P8cO0J8QOwa15WX+b2Hwpm6lhRmfFrs5IlHf/Plj
Ul/r3i8wx+eQUiAIITq95SYvn2rpQr7KWpzmBkVy0GSm5auGc/m6WrKDq+vfwJMk
6Bh9X/cFMwdYj4cJSdGtMWQ47iXSKW5PZEi4/hVp/z99OKY+qHqON7ZW+YneDLoB
0UtEUZWrxRc40D1rpyWaNxGoA33l0m5Ust0lMXtVqSmjqh5Jh6qDCL7clfTfaaab
Tbu0oA+iz1j9YsEm/vqWbjpruTfYFOt8LMdan5N6nyG2717GdFDFCVSou+E/pU1r
aiorkSMIqt3ScDjMKd3S4hRiyx4qPP+NqCbSsptIOxUr97vUBF6euF0kIODdTvsq
dREBiR33DqEme8YTVUlA5UON0gzczUx1h8MwgKu9PU1SGJmfR8N2hKhBcDyS58uY
pKTeOz+6nf7a4pgXx0ba8tHkgCu6fg4u3bFUCsoVkKedydMee4U7tPKTX4CaSDzP
qRgCvbp8no7Sk6HYLuMPdm5FeG4QwOQNgn+lzLmjsR6YBAhB0AdRIYfUkCB58uil
8q1fXcidzPSVsWUzHSQPQe8+usf747hL0QXg0z3Tey66lvzfb4E73qqHJbv4Cq03
z8THkY90Fei9eVVgEGMGBAVOqx90leOjt6KFy7vZdwzae5bxwJVSZIJ/ud3Km8SM
Y+S6w0R3UcKUKawQy2Z+bzU4UJBjnKVcmoAue8o4nKZcIoJsxIe0e5JtLih/tg1A
wgC8qsKMDVxmjMz+TvH1ppthuP2bGxxvYyoPuyPy+RqBxTBln4JbXStRwp4A7YWP
GDiq9BSX8TdDkNMtglROzZvkUsf1Um0S63DDA/vzJy91ydrmmwogAxiffk9scPjw
TqXkrCYUfCRY8rj/+27wcyz+uPWd2yAtBxc1LSlMx1dZdKsiDybmGtzYsuWjpWQ/
NN/Gru9eFW3SMrAQhxAi+KVFpu4XJZfzMjFt8QO7jDe3xRQhG5MV8NuYnECph7Yu
cEVGfFCkDxCajognSipVI/Et9pPHvQtT2tqbYQbpp4LkDlpiyE6g/tXJohPKQfQ6
uc/k9qrjMzCPvpbMYbV/WZDmI88VA9u5dYuNbHWY0UsJl1BSwJ8mNLAFD8vlz2oY
qThc8jrdeB7lot8StfxqumjNu9EOtElNfsuHDwnvkkumye553y5PY3ZxZGESV1Cs
MhidlPtly+toPrAshr/nYUkjLWOpwk4zvZmQEJgrWipWWv6X/YYAhjXczhvFng7M
dQ6ifQl0sczr8sJI8TPogzyvvO0+lnrwcSFDli/9vfvvtOLSuuc9WZoiQARVZYdb
t/+H48l97FuuAewG8in2bP/YMunhrzB2BleLkRTIAdxHRnhQNAWR5qzm0SRpU+c+
8y5wX5AEeUYmUp2JswktsG6h8mBc4G1uvVlRkPSksgjLbz+T9RY5wNGo0umGC9fy
ZV6NkNMpNzNFxh9q9ZFfR95g6jBLkuCrNNLXey4xxWhI2UQCp2HNbNREcHrzMJmt
1JEa1WlVOFv8pu8nQjzySOrfMILEo+PNBP3WfPN6dsikqYyATfx4vQUXGoCOdz4H
PqEehIEfQjnMuxVh0lYj+BUo5dDRxBzhlzDv13wwVQgqYQJgA+8ObCNgMHdBRIqZ
YvaVPpBORXufk7/2asqtvA4YF6vkJBIy4y4uKIt9e3dWaED8uArn/mjqcjjPUC3y
wVWqr+FQfwNXadoxp6R+0pjtkqZ6uRaXTwaFUTea+n4zwCE5e7Ai1CXFx+uioUbP
HpemtPwwbgU0i6xfxS2BvRYkitO+IZaQabOhBgo6XiejtveyyvWVU7oNSRPLp8ks
Q8YXsV0ynGDZi089G/0PPQ4kmIW87YxQAIG+9A2BqBEwGdvqzvH081Ko56BaitoC
BNtUMXison5uguEGYQZpfBohj+1otyE2ZCz94Z0NXAslZ/FJNBiysNvqozBo53l3
46+PTI6wtSNOf6dbm74qO+HRg0Opsafc3yHmbP+RQN3JTQwrkqLzWC/KDbKF/7i/
aZbhm7jGnGcAD7+y1+pmnh0p9PgFaOcQQT0ZSjzQV0D3DWLpO9X/LvRaSCalnpUP
NDs6mr9D4XOCbBj4dtrB/4mmz99oYr45lfnnxEeVAxjLvphRgxXgpcTKQVqzBC7H
cYhhFYJ5WhaQqyIrhusoFnWBOE1u3hLNrl0GVrNXTZkx5Ay24vM968i6g9oPIzCJ
Lnwrb7ycBOfWeih65sDnyp6XujyuX55Z65LOO6A1fckMKKmXPv7KtZwbv4Z5tvZW
gX369Ap6kmEuJdu6lkae4r33WfAju/FvnGg4U8k83HBb+xdUYHRELCY0w/fZISKr
nzbaDMpOJnGKTabnQ+jzQuJLmOEHi7WPo2khWYoXQ/P80+4iH48JN56uN079pOn3
xviROoZ3X4FeM2bqAUn3G0cznnCUwI07igBnoLC8BWDfSxH5roTIStlybK4CPKrv
p5gqaJe8jyc/orjH9pOohKZXBjbK3tzWuZpBiXBM9gKRFKQ35qqe1/LT1unLiVaZ
6jHkbjApEHvX6ChLgLLYLdzKjCoGvJiT7/ihKL+PWASZq/EFb+VjIo8NeoLrbogZ
MPw46bGogHC1rcy4sv/w5LRU8zLoiIzVr2XmnNGHssLpkYU2qG1aUOcJABSm9oLC
H5fvwL27IU6Wk+3Jjn0RUgm7Q3gZlOzTl6kjZg7a+4Bq0fLxSRFp0WLztN9tnOxM
rV1AbPX/irWmS4t7BIaA158+AX8mZabodYn9+OwEXyL292c8VcPhvDVRw7WpYTow
l+PTsCHDQtztebslrzASpe+qGv5LOvn0HxRKAYZMDZttKdtM4aAGn28WydWCbWi/
hBlIh6ePIsXAgaf8xf8fXjPp9RX3M6APB1E0PbUBzHGfW+ZrKq7MrmlA6rzAG7G+
/sqcawJHRgmMG4bhE+EuPCwuLIVbYV6SMGNh9CYoOxPpG0cCvz4irbQfkeNeq5Tb
ibQ8nX1hL6wkH5/Igo79ArbgEbgL6+/fy97x8vRoEmJH0gcjs5DJsmt/CdmWpls4
6MEoctMZlUI2LzEzg9B4bcRWMNiJtbaJS+8uF7Qi2AavFocxcpu1jYjc4v31biFW
GEmk0AIK5l7PuJ/0Wl7EOnC64qL3oh3vXt1iyUmbhBuKIgFveYGGx3F1+SXPLixP
YLaNMsREf4QMX9y503PpFFoPvVK9IE5JVCZ1gv9J7VBSKOu+FM9yYwRGMrGbEkH5
zkvNGt/eIkNP/P1Lfj+nWGP8GFtMeHuR1iLpg+MzMYTl9huidYaL/P7mS6p8/Xq+
6a1w75EILrQMAnqlgfCioJQVr+PXrUaoQWvztno2tuY+gJT0v8Gkc45ZRZc21D8m
+W9DiqWEGHQuCnVhDBNZuwlv8d9W7FUZuh/zDNCvHgY4yxaPJ1isTjgkwdHEeGwA
frsXVhMuzflMyIKwvBQdWyIOXWt03c6x3v1wrrRY2VX8RIfpXpGbrOFHrDfwCXDB
Mfnn9jr7oNWz7TAPweiDCPDko9yMUmIeJH/Hn534EXBhOJ9sGm/jYTfv6bNEW6/H
2npHWpwF1WwQVYFMBeCQdRVJEu13emJAYgsplqBsKMzvb8FOgCswmYya4E1slNKT
SJJVaFDho196JFWvE/g26ToKtPXfXcRyMcvrg4fL1lOVsEaqhWurJ/MBlBWDTb3L
TlDAsLvjW95dBxw/mAChmgbSHiQXhIF/CdbEFSafvul4SIJb+r/N4x0YCEX3qjmF
DgnTPwP0CCxez7qw/5nX2uqSzPskk0Jsn4Xd95hTOFpKjuvdXk7Hi/HbnrOFHZjH
V+UkOmObbVcRcIOKbp1b0TXlWbMrukA78D2rcGNs4jewaamBAGy1KuPNTxY1ZJux
AIkmmwgmKzpDHs+F/CfnqA+wQEqJvUZ3ZfvszSbEIguCcn3qVFHDbEerH86N7mNE
7VCznezZHW0+LvMCMOIFwq6kkw88XN5V6wTWnJ+NuUsSPZGo7LS59Aehh+81O8aw
psCkIc9hUY5QLuix4dNdvH7xbtXONIh+/wNXl5Ij66l3NOZYSwsnOXilI6rAYCWD
TVtZhlpGMzOoOiwwl0kULmhcdN2f7p8mJtnS6d0HDrLsi4VBngKOkL8w49+gPvO+
K2zYAUH076Y5veak/n1vt3x7KIQvEt0+e37vKjIAy4chkVE+h4z2Q0Th6lPQjASl
gUO1xrELV4TIyNsdwO1+T1Vxeq5e4M9f2Sfs1P7zym5ZJbvkpcpzOwcW8t6FPVpR
nzurnLWMU4ml6aAyRzeijwNCF+9OqYZVHh9rR2z34b1AAE87ltAfrsiZ1Qy7nQLa
8uH6RkRMHgRAYq80PnjLJgtLb3GHWmdb2VqtptWSG0RpIbbkM+xU+iE5Ck+xkHt3
NA9lkLlLrvoxWvfS4NI1st0uPRFY9tECMAGNEkQwRA/ngfeo0kGCOeL3gweEFumn
ETf9kH8d0vFud+ITxQspspU5nGdJPiN0oXZjUieqcnAQ3sOhINjHFtqQTCvkPBUY
gvJvo9ozpYudq9Qf/FDkzEMHCHgRnKYdxLmzN5aofLGEwXmNSin9RA609FdHNSDS
I7gEKt/0c9K/eMb3eYWurOBdqPiQ7ZhpbGHBacyDxRlG9ROfSERDYwg0ohsG8AcP
/TNJfNRwqg498VMKa5eaF/fgaraXRIsLf4Ua5VkUt4OZAdaaWD7TuQVZBNm1Hcvp
6x3eKzaJPMiq7LSu59ivRsEuBdksix/iFhP3k7kc7E+QjlIN36vE/ozB5frgUldJ
1JXRjIAPCJryeX9Tu+dWnj8WQkG9V9A3b9ohmu6wCIaYZ2T+EQxhv44vTB8LzG10
oxC2NbcawHfd5ABciNj+IP+naAnrEgfB7PrBkjVvws2GVC9mGZEy65BP2Yg2gSOk
H4rkWmGCCy9hM+dN5GclBdhsHax2HMRRzNe9Wb3pJV01YIChRtGUXvQ7lOJJW5ev
Uygi7vVd7BliHRlPyBZgcky13PwTicMn1U1Q2UBjY730JYVNyK6sOwsXVnKQaq5D
5VhUjggLL0UHtedl8R9Pcc3B1gNHNWjJTAbiTAxPr9+eT772ZVB7ZED0eFIqxAe4
wH9mP302i1P+bn10N0wjw00y+WVb5ORFb9L86A+SA1M3rI1hEWnOWPiO7OOOCdkm
cwuYU7M3D9/CQ/ccVSY43Dh5jZ6nDtZTbslaLiQLQlg0i4rqKuj1USsNAU6nJUuL
9xEtUuIQvDtxcltgToaN51/ZfmHpB/tekDRSUSZXT+x/CcEyut6RDeotpNsGVn0p
QPJt5nNflJIyiYw8M5W/cKBRb0eDuv39T7vhlt3CIHVFj1y8LU+orP/wWjX0Y1dT
9hAGXuWH8+7UcB8/auzyv3P2oo7XCLj3Mp644JuERfqWyBOEiM2MqlfsubjQgY2r
Lm08j/P5K+7yjNCSjCG40ttLW23Z68/HmGsFct+Q4zw5iPXvhQpFe7bToVLPE/yM
LJaGbokzNonCPgwKq9Dfj8Dx+3WEbzP2GQxbizRV3pahdlbWulfnTf7we9TpCWFd
IhcqdzmNUInuKePm8sGEp1zzdEuxo5tosAqqvzalfwn1ZPNmEhXrO9LxFmKomHea
QZs7nXEDLowLL+zV1rRVL5RgD0rjVsphtIKSpz9KI+8rWufqMNiB3FSlUH3tEkCC
PEkz4IIpQKgjnkRW0LXNCNIuSw+htFX/9ep0JZVOuqhbjwKimshXPUTU7Z7kJwB1
gRiaraMVken3s9aERxFEK/NIrxYWAFbZasNu3V45bMFNDCky5X/cAYt1FAhbT7LA
OTxQj2wjCKvtYOkAGHCDc6a4+ZYQVQHN4jiDnBdza3gIALaimjmm+BJUi40E/cj6
M7cFfvaOPLiDIAwFPS7fifoRZrUTooQEPryZvD8genyfvCknH+xc8mDbPreM8h8a
mF8jUZkyk35tImK5uiqMeqWLZuXp6HcIAMzAMB3M2Q2fmF/FjPVBhR44d4G4B2lH
bu8b//Mmq4E/0U/McgboxkpYYKOakARidjwBs/KyjzXq2DC0QqRcLeWyTVKjccPw
FVZ/bgsVXmGW5Fg6b4RFc5/Y8CHQ7kWAuhUCo7tkS1+7PvEKplRt/DlUqZUIh5If
6pYHXkAroKF7U6PMFM4NPwmW7YJB/LiSt9xCFskhAnMgGpt93j9KbUAIM+67BxsQ
+ay37bryj4GdrkJzAhhueWIdJlc6Nb2RJF/VcZyvM0v6C1vtJPn3oDfh9aUoAGfQ
wUSYjwHyts6+rCCxVFBCtJbK4W2YI1uk9PMIQRsSto3VwTmib/mHkXqmeLC4VB7B
sTwjYprmQBQImoZCY9ayaK8ycqLGW8z/tKeXx3vHtxcBdpwjEy1ptVVZBlTlG/sd
iBKLut+l3SMW9230yOD5r5gJWN32/PqK9awCVEjO/kPWZ3duFyBEaYw9AiZMjT20
zyALHb+G2sC+F8nTzoHqnelfLyEySRTyAPc7b1c+fS8/R+WaR8I9jfD+LbJqvlfe
wsj+K4yjc79ikElD3mgdxiLvsebxm4nlR7ffxy7niu9aBjqheelyuKt9WKdePr3J
uPS+TDdHV0YRFuVDBdKhbzLz8j2hFus3nCC8Q4zk7lm6L7mdnbTwXnajswiYWHzU
D+QEb3eK7iWD2qG5F96CK3MIKsxW5RG0nyrz0I2JXBv/hBHYPxrwQ5HhlE8liJOC
euGK3ntqG8vSJU4flzuxn1YRTqmeiEPVAcVTlewYvmSnp/yKMl3IQMOpRS2PdvB+
EZ3rbGbF/9eq+ecIMCY7RgGa6Emj3RkyVdb5w/3Inkp4t8A3rwLxJnpHjtEiWwbq
nP6ZdJBxhG4GzMTtJ8HBcbBUDPYndxHN7hiCNL5vWeEkaVvLa1JIW6Dc24GM/53F
s1+SVSpMTyV/rwDNCFaNltGa2bwUG8T6c4R+0AhgUCxc7t3HIReW6OmZXnBcumi1
x4DSPbZxs5XwGkmAMZjSUCspiFvyLnvncZp//mG++qAy+fcECGUxuElOjRChuKvR
Ag+v+ISM8vXTyzJtgdJyY4LDGRheDtdejL8we3cJEgtF06vquuI+WxFCoa8NYAHS
cep78lQsklFwVOrtNCcuiWVlooz+u5i7NqrmTlSOT2DZvzCGeh4tbEFeLQNY022v
EWfM3suhL69/9a4rNxIULqZajOPJQvg+eHcyFT0od9QFvDPVQ9cMqKysj5UFVXh7
51RK/V7rubxdc3yfUWL7wdbkLKEkc3I3Upl8sYRnY4jK1Pyf41QE0CDgOw+5gW7T
h6NUXAhrZ70Ln9kDd2Kf+ITbo6y//tnqQIZLtUIOEJO70Q8cEbhyVXQw1diMw+Kk
NZcElvKjPkjS5IPkqTHC9oNxHot7GvNIEJt7sxHi7fkV1AO6ERv2NHuNeLomWEoH
D7PlSONHi/bpdMJBsn6TmPCBtx2tx9HHZzS3X+XWxaithgD/v2fDZcooGlxcagIy
AMoozlP5R6WeQB5mBozyesJ9+rw70/vfZkUL62mAGS1vsKzkQVXb7GfULvyvDhoX
64BjTo+Pwlwx4gp7j9+Q96rAjVqaTptdeHMV5FUjeE0+E5lbHZoqNCTS2KHpfbtI
DyoFdHbb1o4YSC+ydk+BiMtd2ZP8P4OX9RorBMLRruZxaL31fQKNe6DXxg4d925y
IcYydgf3FoOgcD1aDvQ3cubvvTRRvAz2QcyFKcpDtz1OrOpwiCCggOmxkzmrkvZU
coXWx/aoEOT6pKEQshJzlyG+0W9NXvlMvDPJpylaaWYFfQRbE3++kYp2KVqNxI7z
6ASzvsCECyEuLn/b7kexsRb7RwMfep1OzGQNGpOdKXravZtOGBGME83WvgLXUqTf
kPt6wORqD1UDx30BWXbxCtSt6PKKGs1tWOXx9NP5KnYnsZhEVYvToH4aUjJ2qZ4t
9GdVhJovjanAwu1BuE3ihShjMbfvSL3463kJ+x1jPvw+Eo02Liracy1NbALXOQFt
hOuYWSQUSLlokpnoD7HtMJUzQQF9aVL6UJSxukFibg9x06wWlMCAl0eEfOM33EXR
Ga4In9YJYqSsT52gVCS+cVjsclMLGBc2bcJJq4YEaRcUjTvBW4ErGGvqdplHjCtE
PMRocJiyw24Hdx6OHTYs/5WHr/kZdzqirSId4pXUhB49pOthzT0hohXUCzRE850V
Y26jnPaX/8BhNEQ2OcsoYDkbgCoMUXKhrn/9BZ3K/4vDcN0R38gBcAT8MfHwiTCt
5geT6L9XZ0MvXM+wkuB7dTY2qO9OWozmsSXCImXugCS0tR9QbGPS2L20B61hRDVN
mBVlY12jYe3988aMsc0rwK1fm+46mwq4F4Zsj9PZSTJZKK1ukJrPfC1zldNhvvVC
g6yqhMwycOrRiSBMDGyAdDdJS0DtPd8c/RIk///WIZDWb/LDNWLyNrGS5S4aUVjT
8iU9+74xottguzhlocVv5mgKjR2uKn/qX2bObZaZU2DhuzmFuIEoqRc22PIzS59Y
JfedevNPTLNkE4StNeGfHT8h07NII8xOhYdMXQmCQYsM0+OyvIbJy79H1jcV13lw
+XPhrWmzgSIhkUfLQyLBJtHde8io0KGvVQGgHXLiUEfJ9qthzvEKMhKa0/433GuD
sfXIHvp5CzmtqION8IeGtbEV93mwSZagQ9SZkN+NmPV6DciJgDegiATBAvB/c3sU
wID4nXXRx0ZhGBKLhmUqmbKAU7zgoHDNsFLGB67XS/yV27bVnLywRnYsO8Ws7Ssa
KGoxCNnjKRjZev0HcCaJqvnwwIpaLB5w+7D65sngBNo640IiMvg7Jh+8jAIYoLKf
0NlWR7wSAUNbyFNws1R8wwWGwMp7Z3awTsgW2ilS5yHbUDHiFiArlP9a4v3pFVid
iLFmyH7j8lyPwnDpP3FpXeVaXWQHcjfn0NVSl/qdSMa74GT5c6vHD8oI7iJkrtFr
N4TgXo3SZI5d/+ExShwzqiGZOj57V33z2HGU0mGL9T1MtNujPRYU3yeM0JVeNIvk
vZ5aEFnCWmp+xfQS6z8g5wVRTxe/1uj37aPQi1H1J+6J4L+kUcBnw1nzbDreHhrH
5QaQShzSuV6YN3+Xm6C/tbwK3Rb6huJiTinyzykHMAXMXsuQGU8ZpCEwp5OFqDqE
RKgmY1fD4FpdDFDH7JzNJUgRyyI69jnv85kw3+sVepHDhNVW6KYBY7aS7A6Fz7ph
2ELUn4tDtbp3RjwDhANRlJnaFnPQ0KK7kEmJJO9oqZOnNoOkyK4Eeu8YbY38jeeh
yhAC6NzQU5Frn0zGp1tdIZKMCpS5uqQrkjJp/B+rBttykViZGFlT4BtC5eJbk50R
v5Dka7B7SusPYEogELjNPk1EAkvfWN3dh++IvzaFA011FvyUXPhoOFTeuXZPnnRE
FdPhv53y6BOJa+4VvZKdK9QtFfBit2DZ5w/qJfHALyZUSPYfdlQ1hxRMccjGe75u
JmV0cYr4mdNWDG8T+M897IdsNjXfSTVBzswMBAUNMBmzEEQhnTMFNSJjKL/o0c3p
xthcPdALYz4LRGX5r/axeliYdi9QxuONyasHPEKy/sp0m8FFRvjCjqcG6qBi4h50
69vBOk21mxfIeH9hNM/FpGTCyBTpu3QZeHi0v2XzR3lGNe0QZ+2d11UzHHf0pS/D
K1brtjOxlb0SxC0U+EEFt9bBhNIaKOHcPw2nddRKyp75EPyXam+Xeg/rfGM5APeV
I5w8UDW2kgxbVEIv1Puq24p2ZtJtrkvJ9k2OC5ZEzCv4TSVJnsbYn4VrKKMFnJox
tPZR5R5EU8whfO2P626h+oUQPffbBQDxwbcbPJ7U4Z8g+JmK4gQxCNYfE99HNThO
vom6sBUTWFTTSdgLxBemQR9tzZ/a1s2b94eKsAW7Ez81fTXImywBaDqJJJMWT2uT
/d0+MMbjZhAmtIR69M1wIf/8oguGuAKBmmByrwCR8Xrdj6cDZYrfmRcuHeco/tzn
k17Oq0r5FVMlNqReQFkjdsP+4P5FC8ylgXg/PnPGGlkGbE2BILFnLFcx9CIUguFd
ilhbX2Z93917i+Df4SZW+8w5F7zuu2SsedqcqpNqblkeN49PQmqkmJunGehEcTft
C2Od3gP709Zot8VHRtEOAcoHWRU1ghxvXeTtAX3x36vOyPDuBEEYcFGWv7rA6f9w
fQtzjVyirEHOulM7ndkorYQrXi19LsBiSQefBTWScueio6EM9zap0etwahvlJttF
w5b6MyXL/t56SNNhTtNKbEfTE4YPP4j3FqdpWW8+hRjIUBL06V2jHe1aGDoaHlbT
qcsS589QCtbNVlvL6oLnBPsneQWuvZ9x5TcamaRQkiKJw1zX+Y4gckNk/ANBcrL/
+IhgpD/glUiX2dUxvVOXne4fw5idoZUEhfxZeS9wrU7KsW3KasyRC3KPirgC7Ee4
cKo2npdlX9+TaiOxGe7k1upqhzyVpE6H/60ZItPcV+ykSQWPKpmDJ2P1L1o9sSLA
jIeS6/dQ8xR7rlW7tZ5xxjLdiF90JEoiajDqs6JbRuuXWCxsPRKOJKQJ+zr0xiCp
NVO/1TPwOIC1L6/GTh0EkquOQpBRzCh6MSxWWYvG8FqsMZFwizibOMPH5cly2VVZ
PyWjGv+CIiW/FfcUR4WhmCvwRb+lSdgU9Xq+EAiPW3uKXjpnudSjnpV3y794LS8k
96TW0H8PSFzCf+rsHHEWZRkAS/AcsyjL41s3pDQAXt2gC25hxqC2i2ZueZAk8sib
rikjaWZRTMCCVvzrG7GqqA+5QXOOO0l6W5Du5mCN2wXrstk95shHB+x7tpA3hYCc
8AdqOeVtkTcWvrI7ZYoXSIPGsPf0s4ebIudxtZG/x+sr+SGSgyX29sequQRXJI5Q
DCi+RS4LgXUGNEkY2YTzOCzM+EgPLtIgbWzWqoY1FsR2UE3oE64BLrVywSeaSzM1
dwjru9Pr8J1wHr8Fc0vl1a31QjMNhzGFJ4iTZHjJTJut+2KCY7ASuobp6Hs9/6p6
ZrxOljBaxTKAxqXYudecCOMzUyjclLtxYrc01dzAv6dAk7y2Ksbn70e1bhWcriUt
WLAKeXIWgrPsNHutkYE5+o1AOsAb+H3ZIXeDG3a5dJg38EtvDdM8qcPnPDmlPp1l
oU5JvJH9wOVZH+wBSHS3FCyoP8YveXjC8ekHu59cfAebtpi+3a1hVU2hUNCwqYu3
4+GIcBlDx40JyXStanr/mWjajVVEGJQr3kgSNaRpXmmra4BYZzhE5kqRmg6+S09q
tI8j8iy0irJsol1Eo7s0+RAH9zYqEw11lhECor7ah62DRR66PCSTTyo0vtVT1mh1
XcEr9aO06NNqDkYicnLbz49N5gLG4j+5PaWDmc9xsybCMbBRqn8RkU0tp7sAiVp3
x0IRWSpHYEv56NkOWE2RwTAXXguXzwi3pwL3hXu9DPYH/ih6zoLaxUQFwZpoeJE7
xXZlWvdOZIk3ca5Yya34b7kbs26w2O9IEItpf0ynB41Gz0RIKvztnD1rS9DsLOq+
YqgVxAIVVeNZS+BB1wEaF/om2PmMEsQ5FwEkmhtW+7SGFxgn+1fB1W9K2ayTswK1
SGyD7a8Ymqq4yWnvBEEAo/BZ9qe7m0PHCW1lU/V46aalgRpSFcUwWF3lx71NVhoa
4pVTYgmLpB6YsmSm62riLVsbb2VFo1tDl9SoJ3VINwKuovoO2wYBg5uNKtzHLRG+
LueScKTUKz8dEdK/LIxcFVT5UXbwO63+GnlQ+vYb3rjJzbYkmGXkLTSFfXdI9+no
CL11dcUk7CCQKD6nZX+AmBrbuh084tOttRZzANajcEZF2uCAD+X+wcaKvXlzCqn9
1q8rlAE44qwvH4e54X47o1h27fI50g3mPk+T4W9p05UKPA0FKLPTa3axyrA9t9cY
DCxIFjkE7+Qhfu5s5MEdfTbPwjks8gdEFYyKT5GPyskDgcSFxIIfcSq0ifYI+jVx
SOHoVOpjmIRlNT5wgklK+JBhKQgAtxAzL/d6GbCVZwRybec5TlaM4XVrhtirx+6g
IO581lwgLRcJrNSsTyepUacSVVtjPzlVgNB9P8Ra/LfnG1F05qvgA06biqZ/yEh7
sTwnKtniNkIUV7jlzKFvppvAfYEJ3j6OmeQUHXT4GpXuxVOG40aq/9Vn7X52S6G9
DTYN7Xzsopn+2fa8+NpUBtdb+oEdXyGoq/NHal7CsmYf+t2yjPohC0/KXSHK4uzd
FnjUv/S5E9VJIRVTMvg57kHmvJa1X39IHwYcIVumVCECRd0frJuAVZiYf4SXR5VI
gzMe2/47KwIEmUhrN23bORhDbutrrP2H/vniEnXwxoMJuCayNHSboT2xfodr/hAP
k2jJuH4if0H0i2APA1093irrB1zLA+S4x9cad8+WYzeuJNyntXkqltAQASsNlvYc
cyFJcSwZQIfXtg/vdts/FFfuM3y3T4ioE0UplIjorWZ1t/qgxXFIv4BT82rER3nq
khAcHCvT/Y9Prg3Mj+3Xfrrnq6bmhrTT6ojL+CqQi/DDJJIyEvfMjIknCZRCr2kx
/1kU1wHcIGe7+wBTjfoAV+8/gez1EtppVHEdwSXh0Amc35ZdGghBGs8+Iwf0HE35
qwRk6GGJPAizRdh6XbmbFRiX7oGZW4D52oUMx+DXe7rIaxWN2DSpWRxlIV3ldT1J
gySDf05vT9ytQHN2J19xcaMBu1oMvUSuKEE7HDAyTII1yrHjxJ5sKB3W/lgHlfIP
ceogf4PCcplFbUeyFF2SuYcogsBRPt6E0p5x2l/FqBLJWw+9ZTNCkia+GBb7+AE1
10Zl9chz4aARS0TUshsmtwhkKJOC7Z9AGErMXjmgX1UKTaEYCqkP6ZIcD0iZQNgT
FoTsyCc18tJIVga69NZwd4XnX3ECnRLJvOh+zl95SVjvsaU+g59PlfT0amUlQbdK
8nvjRo1iBme3ITIQcGmer9aq23rcJsWKZUka6/1P/FihuLV7zXPaCZAK3wXglUD6
dKlj5ubyNhn+WanYE6jvnxpyXGv4Ly01niISMXYDroh5zhOwNxbLgqmSNgxKg+dd
pAKtUWCcpLR+rcxcB8dbY5xO3YpqHzgitjrkoijAA6AvarBW6YwWnt3Rq6ijEEde
BPv6cXBtjv3677zPDINif1WywGUrL8YQi0eNaTdmwD8rBTnk8E/9gFMNgcVqO8Ci
r9IViELzc8o4pYxnwJ4VdeLnP0wlotdySgAKESDsgNmR+3m8ke4Kp8IP3yPO4gcP
0DEovKMq7ILO+dxm1zqzAu0hQeIX99CZe8BbKE13EMqRlxiPZgD4p7g74uk55MqY
lb729Pasuu9YksWNXth3l6JTwyk5Dmz1oC+udVN9lFEKvf2L5UTOJAWbgiZ+g7TC
Tfu8nzi6PNVmPlXYoUzYFHls2qpo1Dw4FQ7cii6wxvZARs6XOTrXmlxh391fPDfM
P0O/EkwLiX8o7MBSHNR/7iDVbpVb/ohFKuUmsE3j2qJijUriw8iV+WOtgOq0YWFr
HijXasiaP70Fxw6LiglvLp5wah+UXvqCY6uIfUMsdG7pMTiS7uKrKJFakx8SdMWQ
7Ao4WOdSxEXCsvl05HN7XYbco4L7Q+sBiAF8ER19Vf4U99zI9MAmB4E0ujqISwZs
4RgRRMdrULGCm03P4Cukf7gsxiHRSREocwhZLj5kVNe4LD78/SrqfUjYG0Mc/NFO
GMjl6kdkgAvx2vczPaNc4ohH3AUnGoNepLW3sAmFymXJwr+bHYTzS/nXXBphL01L
33uKj2lpKIXU2puEo8/Xvg2A6QnTTEQUlS2XZr+0EwFLmeCUjNjH2QdxwVhan2sO
9/d2H9S13fPmlOId9YE+eeUok5gBl3xfxJ26qFelDbQlg+d9Bg1R2ob5MTfo9FNF
EbufMe8/OCYZKy35ThuzGtC2oGycnkM7+A5h1dRvvwLoVOcdKMs0fXlkBQWadcXs
ySoQg7Dh+R/u2Dg4xNBJbWLMjwU2u1fCIdKpzemQjO9x3NCiGzItEDJKFfj5d6VD
y2t1BoQncaVSbfYXYc6IqI4jYpV9OypDToBfAiBV2PNQ6p6lLC6WmJWjJXtdfjyz
7QrR78Ud6HfyvE0Vn/+4F2DFiK5tINEZj5hfQTdr/o1lHuNbNigS0syiJeBEGzzc
Hld9GyApYOGZ00KdlCb63GJWoKpSzZBjU8fzEjDEF0V0JPzXERyCVzAAbJpZBV5E
iGIdzkNKPdD4SdD14m13FtN65LqNoynrgsJMTW8m2mxN0LxWFntf5K7RJ5c5GGz3
4fKO/PTS0K6FGcidHQuIILBZMrt3RJnPzorJgUXbvZqBrjIq8nf8hMftuiU17Smu
YfWJ8iWaWnXz9gPAp8KUYDhdCjycpVPEs4xBOTOAZMB/rFGmvjBug0CHX6ZGjk57
7uJ2qhpUSvN9j/X0W/ym46xjS4Mf0jEBdP1b3bkSf4Umrkzp9KeU2HmTirRk6VlC
z4HhWSwf0h/036aHTqHeACTOUy4GI9xn40nyDil2StFeUeHxHAiBoh2USEPL5XB7
WmhrTTzOr2MdY9QSmi6Ch+7HeZ6lRH6dRXKeVfsVioiD6sDWgczpRvxrw9X8XMzq
eKRSM7oVkAFjqTaTWwWNW5v6V+L2XHf+mQSjKcGIqV4jrAhQFHvzBqjvqB7pu5FZ
tOKjYdiE8cTw3m7rqq66hnZ0s1QRkCl6m2bYP/FWLmutWKf4EiCMlgI8FLNMF25G
WmOSPrmrAw/SJv82rxBL5r1rXvIegkGLfY6Fo02HKxq5RsV2XTyCAq2YJFZV1EOX
tczHOWhBDsln/6OOcKvccN7KWGwqLPvJGY3s2ap/gpEE4l0OEQHNIKiQNh7eEgIr
rjtKmHhXk3+mUCT6lId7zqVkJnGu4TP6iTyPkcRFWHwI8j3i12d4n3KlCT+of2dd
gVRO1xCbGHue0kRRH2y3yt2PGBnjvlnq9+wyIljBuy9GqmvF+GmuR/QTKuPF8pzD
+X+jChbvFajSHwBN1lXHYeUQk1qCd6ShAgNfZHz0HCoqRZGtWcNWbbqvxXWJVTuE
BQ5/0AjEzCj13ZtBOb5834wBl3BOgOF/Fpxmc9ewU05uep2xbjgjxin0zbMN7A4A
a+j5g5XkU6oUWBNMbSB/BLsqCjZvSKqpRDRmLOdfKXjkdgdINN7Hqq4JdNjQRODy
cFbtXhyj5Dk+hZQ+FStJ+EwNd0UV3wr7tkLLSuLg+9rrjJuXKg21COjaLzwNprG9
GqXOFYUcSAsmaC/kQrrA921p0Cfmx5zISRhcIyl3jmta5uMkuS1e/hu+i9kSv1cK
K+H1/r4boecRtDBmGTQjF5xr49H1Y+j6FHepLnzoSME9dWUUl5WP0RLVGZzHmLKj
w1JRvMoMVOGgkOYut81LXxP+8ph1jXbZW2cBDLyjhtbGgvPy6pUIEv4SFONKhij+
4sl576cl/mWH2RHfOxwxDVQ3a4jHi0uuSkfz2IauvJtytlPa1bLTRv0cfqGe++Vt
rT2MiRXpMJIS8lLZLQ0Z3Zj6TIuBbj6g3T+jF/GIKziCRLn8mhhewH8tOYoy1Ijp
ijx64qN6jyWmCurf3c8zRDCVEHpoujs/UKI0RdtCyjbPtdPhqQ+9z4pvap9VYLmp
qV8w/8FddF/jqD6AZQH04vPrrLJYvMuzwrJ13/FpxMV2SDoTojtD9Gp5R6mjxGtl
UXtkR4n25PghyRepsMDnTNhh+GJQbbrgsUA1ApLfSrGx03GMzYqUO6izUBGf/tp7
5MogsUsd9FbRtq1jPuONkkjQ32DRd8KjQBKbYlQepu3akH+W7v9IwJRXmVaL9XO0
FTpVmyKxzdTYLXUiFjExr2UOojpq7klZdbKPKWZ9r53emiqv3fn5hkCc11SaCXbB
sCRHXOcQTZql0ltNYI0B2vr+GIsvE00Ns6K0ICbes+/5s0UHZ5r7oYk2RYsfu4QA
dPdZ699svxvfGR2GZwyqdqVW9uZWt0Ipj07MXtyvDNZXn4QSgc3wSTe3qR05WemF
9DHU7iQt03GJL8xCTDNUgeKa8BOYsOBKpj2TXqOpDJ0KLaOnAkppdnnl85IGPgHp
nAG0wB4zVIpTiyjdy+z75Py8CFAKBLGDNu7SvKGY13bSKEv6tUaHifOvjo+F4rRq
1FbbkYNsfKkYntCGgVX2muUdAjPttVbGuctsgIql+KJe42cEWCywVbz10LAFgZAl
KE1ma6JEy0KpZPC63jrr1xDCy/yhhpgqK+kjW4alKz9gKqRcGys82vtqW5UboYbQ
0bggcyCQ3BtFNA7pmDKHOxecfmtn+fbT+NvIDN6e4YyASVOPL4RSI4zMZPtuIitX
eTZk/aKlXG5ZAoYYljK65dir/eBNgbPTHJbvKoCp/oQ98bmhoFVA2M9S/pjEI/tx
uYAtdnu2Qmr9+C4ZMip+BvGRRsa0pYGmeGZ94FVCcFWdOBfMEVxq6tQaUBSAfZRj
6wcAAEXFPTgpYI3cTqu/7cmW03S+OJhBvUF/Spk8w/E/XdqiRZycm3/zrg2kUjg3
HBOkaBcZU1AUpV/dJ3vwAXYtVh73UEdm3HYC6QlZ6YKKH9Cw/I9JGbQnXbLvvaI8
rKj1dVrwdhTdHPPY26YIqyQWEi/Dt0ZTaM94/3xsJvcxgBsgTakiXLakJitb2L0W
xCYRBMMPsskx/jo0bvDaIv5RtkE+cyXnwHD3qgyX5y7AQeArH3LidG9QaNd8PUth
Woc82p6sndYfjxGJ16nnG7781NwwddZv4H8025xpS+i4QLadL7ShWmyU+UVjXfM2
/uWEMWmAwhGU37/dw4Yn+tahxKDTnacSS6J6SCHDZe5+kDHM+fTjuTg8QkwUNklo
9E3UPLCqG+mscSSrdaVNv4dbN+m6WYJlteExfEjRTaJqeC7tswLT/Tb8uZ1mqJ0W
JcMxLXBg2Ni6MivcAGTyGgYrm+bWdcal6TKvaoN4brtH1wfqOxVyx8w8bCOZ7WTV
LjTBdJLzUELH8WI08l6PxJbtB/LAOuc/K82VQEh8nSHRqYhR66NvdMM7lBFhq0wT
Up0pF86QdXE/WG5q73gpKIR5Nf1hO1GZQmLqIM+Zf20fxmYjsjFHKGAIXEcVfoRl
4uktiuFxkpyGNxVcML8YmlOC1dcIOvb8i2ixpu4WLLJbY3FBJuzqLMpCQrxWSlRI
fXmuYke6LejS1xy/BkH5y4iJtuBIsYdhvIi39l8XKDiJTj0TRiLDAJY9ZjyZu2AA
rSuURfiHoj7WU0nkPeQrhkFd2O3p2jP389xeTHIogFQTOhp998t/7sU/YrwUWqct
L+NhZuGKPNqrfuCb1zo+QgUvozhnML8+uOeyndaoMB5bNvKqoI+hjE3lioMo081+
h95+iLA3vA0Qp+BrHobou9e1DoZl734d9zKRSTT/yFV4gU+d4srVUh5MliJBRKM7
ppKNZ3krGqE7ET8OwhLfY/Qo8OQJLEr4gqRVSOMCJrF44lCGx75iXUNGgUZOyoR1
wcTY3nm3f7FSgbXg1AKm3ibP0oN8HM1y0iKHrmYvY1pr9KJ5mrbxVOTs4sbrWTu1
Lh5eKdXUeIkHsDCniTibJ4fh+6w2vsXr/k/jjntcsUWmertPBVRQNNbVLtD9z1uJ
rqp6nMaXZqMxuO8OnxCwcBch7N9eBbVEJ8koDYajwef1sesAcn7+0R2RMfCvSJEl
LdcHPdoOwV3y6fFNNKc/mxPyL06Y4dovDyLqSv5oLL3RmfwhgOFFX0M6m5donLQ6
I4KDoPTVz7+w3L71zgzuaVTJRKocE9bbOrmZNn7g3kPXxrZbNy9Y7oF0gGM6LgGM
RwK4OBlgHf5+EtsBfeQp3nln3hvXLATMH27yYV+lakrwSzOfQUO3X2qy33bQ129t
MY66KhfxlgKVTZNI/CRAFpKG/KjUnEc1C4c1DyaBnFicWp5sZj++/ifdYLxGVvHl
0brHu9Egh+5x5wGC48YiJXJvL9WFd7eBmvyaB6MShF9pqXuWJMBdsqojf1N2r//n
r91NswVTebzDu1wa3WvLDzsd6xha9S6OKLHDGTKwUoe3pUSL2ppMuqlJ3yHMYHOX
VNIBEsclyBUGcT6LjqDRFTtOIO7vr9813t+nZQhl0Nx7t1Py/wA9pH6cIZ6aKm0X
XlE4Xn3HzOWmTTxSlpL3bhaD3j3au673fzBMtz5hgBujf9u3IxMM7dFJ/3skufcN
aIRCPUav/vdtltlw7gLFKU+IRNlwwD2w03253a1SCZFsrjgJzlz4+pQ7R8/wOoYT
V18HuUCWAXoG9VcFYgTPNlUBgoR5qLt4wKRBHSzctfAG3XjcapUMX9h+tdqHRQj0
/ZBEpMVrRQizgQoFZW3CndPlCz7NcaGsVzs3Ds3e4QIJcDnKlhzEc/WrikMZFIWL
Ol2Re06stBEmSvVduuiTkWrPo014aTNpjT6TMyY1nJ99tGh1AAlf24UKl1Bzgj1q
Qf5w4ddCii062EA0XiAaPOUg3DRYuKYjsn5EPneowZjqsIkLxj4f1DrMXBieN20D
vY/0SpCAQxcZNYnQ4BhifA01zinFP8ZiCUqNt89MCJ9HPXsde7dK32azDDdYHeqq
ESCd0/JyJO9QszXvS68sAjaJxP0c2ZYr7g8YAuK+wgoy1LE4jIbAGCpXQGapZRE9
wZBFr3NhTBJyb0PMNSbcUzwrMt2dWOqB3S65+6xg7TYI8c57hoRtFw2cQM3Z1NoH
Xy2+mdLKE2IgJplnJ4QnV5d14g0QYs1elJoaAoK9EhNuSepwuWG1bHDU83H2bjfU
42nzm4wrF726t7YFKpZQ2ryIlteGPyd01NtFlIW9woA3YgHI6Xo9URZe1NRgpEny
1qUP/c1DMtJ4DsNG6/kOPTN0I6RWJHBgF4KR5XH4MCUSOxto/ObvC92uCRRTHMG0
bN8hkrXcQPMk1eR1emdHADUtmBVebNH5n6SQrm18a9mZJCYOvOikUR2xy3Vkuxhe
pxQZWFZBvTkNahLrp+aoIsm5+xWBj78/DC3a6WPX6/axid+K/i22/RDKk7JI052b
VRBdRTYQbpHyQEUiP3fBzUO3i76vcllq2WPnmczHO+mM51vxnntHPo+d5zDskird
jOxnKc0fylb9sBgIbfo63Vh54SsBomcUS7A1EnIFQnZbIgNh5UJ9TzYaYuqWyIcD
uIffayJL+Q07KWi8WvQj2Lw7TgyQ/qgpbFW3lkt3piHHusdSf7+5ucD4a3EGl8Ib
rqK5dYpWF6stRortRaFYCBjmvO1xUVRgYC+qTVgBvxu0VIH+QynSUZ77hwZnfw9e
c8H16IJqkQGOh7I6K6ExYXA+0v7DBe6i3w18+ABlQeJxfjT0Dp0CbYGAA1koTxAb
QkfgXDmEaLUgokXpP8+anTlJJ7T5iemwmv+gai7BgEpEBhvxQcK60U7cIHvxjYoH
xDafrmvsSNY+xTQwRnzKkaWhM1CdDqJDhRN8Nuz6EtT2dFuBXqpuSFIOnF41Kb2n
pQyMY5cdnVPk0EzTygRyXabajSW1MB432WM8ZxADZXbYNY9e4JjTtI3K6AyDkEIk
IfJRfSJchO9KwkJh/XRhO6Fei5/dKkHT8NwXwFDG7YGlWKMno8Tu8tesbzrl3FYy
CH08U8mU0cWg6pcMvaX8WiysyV3WwEZGGVMfXeGoOuXLEX1awN2f7Gmt7vJvdy3L
/IMNuCj/DtIfHtCSG0R85HZDn16MILOq5JSOgUAAuyfxFD1wz6Dkah4OqB6n+Kzc
GB0xIjL4Z31UkdSwb6W7TluQENF3shuIzyTqdK1mmnt2Gy3amietdwi3Ja4ZzaQe
9Vmk/WyDfkZ0wHBejyhCX9ZT95FVhkuPsBYKkKsgLwEHFfJTYTUOlyIz9+vkQCNE
Gz2E6OQd45SpyGh6sE2o4Cv5K09sH8SGYaufllrI1Yx1T298L9uZ/2IKDOW3B4D3
DUvY1NaFUNE3Br/d3NsP0m2OvlLqgynIMotSHburqNty3bmf6Wa6smRCZVwP1616
EjFOVK27N62px+Ynqpo9WsX6WutGbk2fHw/wkYIFxn2OalljH7rRNCvlOd4+9kEc
Qj7xStz9grsPGo77jNgrMWR0wDQBod3XYboXVIwrNm9wnAX5MPkqlNOF3cBuoa2u
qs+8DUVNyXbzVxdphdkxh+nxuHNCpf8ggvxVcWsHCLSluSVhZQ/bAZjJC5s+YfW/
YXcDDAJ1jMsjZg3wVi9hIuBS0cZnraNk3GVwVGVEoviQeW98a/Fhgvd2CPd3matS
f1m5SAuDbFgaYUX3sOAun0sPcgoMRzsRObUoZzRjMB6o+Zd03K5I1RsUcWy+NeuY
OATZ/qQmxiyE94xbr+dqCKlsI9m5EGecOY1bYWSddggfZasrdGWXHIXfseqJ18Jh
rQU8CDUf+UuPp3M3JpBGqzhmGm/8EvvMDm0QlYdBqug+jd0zIEPvUVHRdaBHOi2o
eLCREou04Fd3x/XUGtga+zZYyG9GFz82u7yDNRc+3RLUMx7/7hMKM0lU1ualm9pa
Xmm9RfHhPBMxMz/00C1Xbj7ZC/Ua5lbRDDaCch8NLYHiFjxz4f0nzxGtHu7jZ9Q8
BQhLXxQ+3Ahw+p/e3bCsXCKidP1yek82cIh9QD6rfm4g5+Hyk6wWfDKWtGXzq74D
Z2wLfWIAJi6vttUo9ybHs+rRpI8BPoRDCF4sKHlxBALPQdk2in+aREyBRtxYBFkF
L92qBIBePDqzI9JHyi32UrYIqiZYPQNJDhD+DDmgzeC9BRhGDwqtUFHGwesFXxYo
Jm/7g6MkcSrUDhn5RUdzf8rxImn7+fKIH4QWB5+tagtgWmMPaUnAyzoR60K09Kec
w9cu9s9sP+MYuUY5U+tRLt8UzZR4ZndOMK2fMYP2Ga05xF44fV5LocwXQ2a9Dn8C
Bo31h9BlBGjfYGWgSlUUuvNZLbuV/48BJt9208FsGPWtVpx7/41SRfgUbDLzv9SF
589VJMDqh0Wa+eLi2JQQeWWJjVE86+JJQ6eb+hF+GtOyr4VR7BoDter9oRZ4ejg8
JMuzTaZjdx1Obxi0Bf7C8GIGYNeCVfFsZzFlPlZzo5/C1IxX6eOljQp/5QCiEPLp
XUz5nfDpVOKfa1yamwEbBxfMeOct+nNOpjKiW+nye02eAf+U1nZzS4hdIqLv9vyS
UlZjeTJWbiRT0EPX1iselmx0yTe3jnifq1IRsBwJBg96N+wIqL0JgVQFn9zWlUFT
OthG8s0WGgPzY+UlcJSmTxsojArF8vu/Pv652G3KXWPqK5CfcL3IRpsiTRO1/U3a
9OjFyksEx9XuKdtjPFOODz8vaLBI+Pfjh2WQWWKi8A+b/q2BEdMuyK7ql/v1OMEc
gMANp0pBzF/FZOwTxhrnIjdkDuLLeIk7plw2zs6DEtzz83lmgo2F+QFO3Cr1a6ac
TNxp5Ge+J/UvB3fNp2D4bsZvj1ayJP/uAnX637p1sgUxeCuPVgFS+qtkCDItitfu
vl+o1qd/6uIIkNDKExutgPdlei3qScmTVShQx8KKQ1H7RM4bQ7wIWhgAS7ejg7Xp
+Ic++X8/7CySF9uLVIpbRcUGp65Hr66PU2/QHf7bekKnXXNtf0GWQbaAGaw09Ncp
YczT5SawfoaIfV1c3PnFAICGUC3fIypkpwGChXtBMqIgHxLtkkMxuvFdkEmOEbqt
dcsnEUXk309s8dDOPYlhtby08zi2r06u1G9CNirlHKqVmXkWV4oZjq2BINdnmUB+
QE9h4PERVR41mhj3RC/XvPMiRI0WUnZYndxWp/zqzymsPFtR4o46gWtIiNkXgz4L
9YMhX3DTfQfv5WHjw+tLVi3sdR+aVXz8+/BYELyTfp+NZLXSb4hy8BcyhWuMe8TQ
vO9mc4Ha0W/R9aUB8nxyEBX0LujAlBqVqK9Dmzk+uSxzrAHNREMhMKsJCsTY61zD
BJHtLXczsNF3ULLlHsx8MHre10Mxcs/ZKrQycX9aETPM9T1C1cO9qriS5CpsPPHU
3ImAF/EmSpNQt3NI4DHzBqj5oL2y6oBFOT0hZeeBY5DCQenE9zMAPn3dNdVmKzKQ
20vIeyRDfl9Ttv92xGp5SXARaQd+UkmHjUtQhsfzgWbSfsR0xY7wYmDjus4km77o
dSs1zcV204A+yACj9GgydnVxOFDg7Fl+F9zsa+s2wY4urKISTG71CriSbK6JIhHQ
0EpgOFkH3jLDwQ/zuBKeTvU0aFj2qhBvvPSQRbewtiWNaG/GBHOrnRO1o8Ip6w8D
oayN3Ll1AaFwXxzsymwAvFgc7EFrY4gAqo+VqFN5QvRIZ7SmiWxUZkqq5WElehJh
evGECSSW29DcOluzmqNopHgePlHlku8HY9P/INSPk8vOMrF0fLN0A28lHOsvtZov
iSzJZZaNJrf6KrNgPMzY1R4aeNDh8q+JOp98fnrHsCdEIcpcu87rU/orXIRTSww9
FE3e1UpeMzgCbJeW4YkeiFY36VQ06RR7rYwyJVuPvZqfU+17qNfZ4qSyy/F3CkW9
P+IlmfF1p50lzSNbfyNHVERaQk9VorR/JgLolI1xq6OoLv2loc6/85XaOKfmHPTl
ypCANmkIrqS+OrUdaaO/r7r51KNNd4osLp+EIoQE9qBxZOgv5gepMEu4mXmyxluu
qa0bJqqR8VZFyDr/kxoQogp/gIKRihVzicT4m7UBGeLApXOhp9n7uUN4rPdVSlob
rjl5gzQystnden4hyGt+RD584NCoPQfEw1bQbYohcYpBnEffOzfTuTGAWaD9jnk9
MXwH+FX5Wnx9jNFCLjVLiuzE0uAidPyuM1N9TV1XSaSclZxxy9Jy0ph14yWtwDBG
aIyHZKtNtqp/wSqkRVft+CVF7Diz8qn475vv2X6PVUtACUHjnizuaQTQ+r/tWSIy
b3zlJ2WXRLrXppphWU+o367V/cHJNE62m5nXwC2Q6hcfR4WiLSGa3uXFj0TCk91T
QLcpzGbDjZXSRN3v8gw0XGamXAB+yWMDpfQrpBgPAh5wHppxSiNGNlUH2sPtb/2g
rmKcrtWZrXWCTwPty+4uo+ZVG56tLkhtCz4LUBfVGtgeYXNgVdcCGMOOxtPgSK/S
5Wgv1IH1PbOxT2S0uWNTIzrLyX6X0Kp91/jdgdzGnZVDVy0Fa2+s9Za8HGrrUAUJ
HQ0TMAaDcotJxmxbkE2uF4JGgaIxeCwT/wdrYeZMt4/8HZH6M7oQx2wXAjTHUQzS
nwWY1xewr31dQi81NcwjYkiSJMhCiQlEMXBcFCYUhUf0bz/XTMaOnPS6fYd2dXD8
ri1tzGGhzCz5LVQP1MK/5syePMopGEueJHAiJENmgK/XyBPR0D6Afbe82y4u0ywj
rIo31WzJWsMOi/P+dco8o/Ep+gBljU4FiyBPkS6h+7YVTz3hukM/rMFH4ndCGW1E
wzQSjRaH1b48IReaTaE4J/1uwKsTfYOm+/VEraojB8f4cj4qf9s2603KaAbjabQP
9hoz9CFrXlkqXP4mkwdMrMRdojgJ5/3wD5ynLoxQAAtVxIFKndvffNc30OzYzRHD
+q5EPhXofrN8ayIyo9h3BUsgsB1wkJXt6oSwtIj725nV+yiyl6HPGKbzNwGn0CGM
DSVA4sidX1vdSNfrHbzo1AVwqcswdt3sxjjvBtYtEFDrfULvJ1+JsVOJq7Na74fk
Ytl8jCxqZQs/97/57hl087CSf1BT7RzQCU0iW3aCmozlpD/C4wZj1hIaXtBQPkoC
gWoyRnTgzobdRcro0y1edq/HmZMAB/4iR6GPbiNj14Bi5AvqzBGORSiefT/l9hyI
rRNijEwvS3QpV9b61sfiWMXzZVYBizkfcZYy4HgvpD9TSGjLyR8nV/XRJD+s0ZcH
eWHJ617la2pXFFoU4GClzrR3OoP2PkoZFHpwrO1dgfUZpNySsT/qYQ95luxwgQ0x
hDov5EJFK4ROHceEPeHhsRVc3QjO+Bvxmbe6kXpQYUYIHGWY4yVRvQPWV6JzYYWl
/PDXrn4iTyRhmV9d9L/WsBJu4grz6YKD4avDtHf76E8/+yt3MA0zyHh2KnA566J2
e9YCKj3l7SIzBtCbcSdgwJhvrhb0zb//MBuGzNwqNlocPUFylADBitx5VLXdFcpr
ZuekTZkjHWeG7WItjGR8X1Joha+i2OvJt5SztC4D9EEq1AtuXNeVdi8fZlQ3FxtA
XsER1cN0tyoc0j5c0alJFVEd5ZkiSIhqiyc4TG/ZDNkq+YamWzUP8+i+QVMtBt1m
xiNAnFd9jJHAyUZzk6xlrVs66RWL0wkhEWUysOj9ZMbQkh7YoXT66/yj8qfswnSo
wM1TUSHa/hXXa2dF943mItpA6svb9Impq3JffxYKK5u4pLk94M/jzAUjC31mqe37
P86qnIdyQh6DMHwdmQSLpZSLLRahtMLzD/JJndnht1ngXnJ5kqyHHiEhiEphuBOQ
H6PrV9CshMlXyacNZhaFrrEIAqPgO2rjdwko9Q4Gs/sMb1zMz5wM/JwyejZz2l5k
a2L+2yMVFJZPHesys4fRKxarOmfpEoI2GR6Qytk2kUu28iVqeNYIjxzxyAovhd97
awADZ7V4H3y7JW9Z3NA+jVvLoBrXr+zaWjY6VC7gimd/cnf06FOGQSf97/pK6z71
2BiaB/VnWgWjR7izK7KGIb6ehT9no+jWfylcg1XwPh6MU8KK0WqWMs4RrLwovtyf
c1ctHLtTjfNsOoN5uODUEGI8O8rJH7Ot5ApJFBG1n/RsjrvoEMqEfy4df0AadCIk
9O5UxSJozZlVhr52hQSQ8F1t0LfIUR8+kkbo7de4oCjAN2CCCNx2SzMuwKwOLcDb
CMF53iVvShqEXOip+MRlW/fbT5Zca1A2k7Kh6HhlSClvDmgP0aj/vjQBRuqHOZtN
oZsDO5HMum5nhs9dqKk7hEUEcbJB5YKgQp7NFHKAbPqw3wXUcZ+r3uiAbhhuYYlz
0hT3X/A1FL4wpaqtY5+1D7l8X+hZCG50CIh4LjbM7stos1PDyVRBgPABCEKnlHZd
br1iZb4pJNmaQMAgBd5Bq1DKz2DHDLZXpPXhLh7Oc2WztabGtHy6Ql5DHVW+8OXa
ifj5pD/cghP3ax+0vbkPyMcD584mJ4NhqhDitJ6x3Y2wCVox1AAAN+xAgPVkzVdx
MWjGoX0hm9BSTHhGjSWd8bq7oC5raWO8kMYPvhyzJD9ZZzrh/y1P2V5ppADEzoFJ
Z39ouFvVXtRke+F7A7mQWHaAg6znWVWLY2lb0+CSUU4Zh8MOMOqnonAX9Im6XoBt
StqfxcHbPBGXDdUTITWrpZL8ezAycnAo0EGxxV4AKEc+h7iMFbgTYRdauVLDiZ52
4ib21Y6xh4k8b9E31CXObsAPFs7KmH3l/LQ1m/7FNb1DnTGKFxv3zeLSXXdaRNjO
Re/7Oi1rBTTEZp9idpCv1JXVDzyUsJ5l0ZGgWUgjHRXlgiv7IwEhpjoGWxDIvI6l
JM2ujJcp5V8GIsfXZzlmklnPHu6+5zESIfEqLK0wrZJDt2Js+Bb7wM0TgSeNTMCo
rzH4ZRQ23sDowVmcW664+Fxq11lhuFTAo28j8ucCRn/hTj0H0benLyUeqqdKiaWd
SR+5WljxiygA1jMhLxhR8O4PTRYU7RvJXH7qmhhAavaQY0If8Yxs92frDZ0svEvF
dstFq3eChD9gnlyCgSny/xPX65GEh8wQ5K62gINOvf2I0clsHyC3cv29EKOWOohx
pjw0QifDVS3Y5Etv18r44KfjkGJchDzuVfgpNnMG3sxmYhuOcz6Sl/trNLMT6umg
Yv9stBbmXT+S38j+tp6oxAkq7GemxekToTM+3KRdGGmo2Wf5amu3C6LSoxjm0mak
UplOmKWHMnpjJV248uOvj5FbqxzpzfXyTt5sc0mNscenacI4r0A1mr10vdY5lrxS
VWJfMVTGGmDhguOLS20RUxk9se9aNQWNclGIPh1IZT4+oh6oHKy8SUmMDR6C+HwQ
e8seSkRQ2E5M9O3JEw55ab18qSa0KHkWC41HykmLBdv4Mmi0BxXUNXPH4YE07yuh
CbywYcG9BKZ9LqAXGCXNpIBI/YbVk12IzuOwdMb802QgLwrq124eljUbvTK7Mdpf
3yaynVO7j4I60QG+KMgo1ybsZz2BpYzVPNG+IIttVKejtEibq5K9H3ELZfJsmWoc
icIAiF988qrlQY+qsWgcnzNDY32Cr5Fl4VtKNTQhI9UjrL+ZWo5YqUkbSdgfN+p3
w/P4iSvVcDyHh+OVMGUxecIk5bpG5tTQoSwPyGX0PIxF+89+v9F+udMpFdaK1rYO
UX985jktNnlbyywzm7klMPjQ8YSUyUqG4Abfg9rYSBhbYdeMIAZGfDlIFokPb/3A
HXNGcfvEucOncWR08ej9yUoHwf5W4cGXt9jxF/jjsy/s2huvSGRavsuHueruHgkk
e4YNL+LW5fIxtAJvUcf/31NkXgyd9EomlYfZrx8jBun1R8X7Bc/J6KM840efh7FU
RuYGMrv75zzCfv1374PoeZY1yIVFOfDgBo7yikOcd2Sz8gHvxOiCbbixT4fL8E5O
LNXa/f0EAQF5gyey5Lc+p6jlCbsoETWTSVyI6IMk6Kvi15MGNiWG7HoKoQGD6+LP
wuXGYreiE8aKYDEwXIH3uAJk69/6NRrv6f/t3iAaI09zDa3s172eWbFhokPv29Ig
ej3cvt0SJAHkZ1x7f2MzUgj/e0X+zlFA5wsgP8v6cgvJlqp9zgkyYobmEGgyU1zR
/HCns28RDHigxkUGrwbTLDdmwL/3sJKdNBuIt3y9n6lqj4K2Oi8jHj21d9FISs6F
FKZZ1caBqEKyAxro0egl4GrFPNK+iriK354CY7iUttFqdnOHXjl77Vq0igt8zXBi
nmvgeVBwiutxCzpeDzLX8BfrAnOOhsrJR7csRIe/AWaWQVuHz5cMnTD7OAj4J6+D
ES4KDF2rTtXYAk2pgbbtZGOxef0R6kfuFupV1YRzuTrTfrj9DtL/bOAbirIqLudP
ltteYkxKj7ZQX/yBygdKfxlVsS7zLbPXn5AHpPr34Nr0exVTwx5qY/SSZQhbIt/T
/un6/3B70SqO91/KRtCw+kAJkodBhpPPWP1Rp9kzs1XMxZE6tC4+BbFmFZptyFDG
TI2Ubuo7J/MAbVby9RfPoCMkldCjo22m4FU2tbB36U+oMzTnufbs5U9UtTOF1lHv
sD3R/oQTNNvFgHAJIe80gwCEUuchxa3MS+7nFjg2A4qeETlD2Ju0HhpipGStFlfr
y3A+KuMLq9tKSAA3Agg3Z1nsaGzdv4mW7+i7cR/bF9f+zEeoBpZ8ILNodLKhPQdJ
/pLAzfcZc1sDnQE47YkW8KxutPheVYm9dh4/JcmVaK0StpqqNq0v99ZwNLi1ATwB
TUZxe1YM9SNx82cRqvsued0Ri01O66D7HhnUXYIa/NGqiAfWXvHUNzf29V3CGdcE
Q8i9rDdAUmQmfv7RmVnygdpNSi7xXd0+eX4W1xTI7J1VPw+GIMOiOm9mGGDI2bEZ
z/O7hhqeL3f8TAa4PsbCVA/I+D8f84haSB1JOhXNpVVE4EVa1kqMfNDkH/KN+WOE
fjYIo3lV7ZcrcbA9qm+Q/CdksNwlkyDmuNR6CjBxR8I8p6y3eNez1BL72R74bz4z
XXmsvReLBCebZi1Q3gEa1FTLqV95JR75kabar0zfZlDE3CGpXZjEGG7gEna4B2uP
lIiU36OthTpGKExuTTzgZTlnBY0Wq9PUGy5nqIwgEMxAHSjJZ/yZDviSzGeNOVUM
8D+7wgjnuS8cypA91MEYhM0hzNBapclXc47Qdj0XLE04adPrgklb/nsibR2KLWYx
rDZpB9y4i3319H6sBS0ghZ3lzfzr4d6w0avgtaBbfHBZnxbcr1DeR5PEBPfNUAcC
NoKojwkCLaT7RtYYf6sNom5lyseio+tSJq+6R+j+auuCGit1ysKx0RxHsjQQ+PDN
aQMRQoq4N9mMihqQF+CxKi87goO9nwNbcCgzXGdvANTEVXW4/sfjVEkGwguc+swd
ri5V5Ng1IyZ4cyF2Z0aJ72G6zmOsTLNbJgwFQVSDjItYsJdJLe3phqyJtpAzG4AS
hcBapu1MhjU12RWO3lav5nzqCYe9o6EulYfTQynzAoU1AcoN0yh2X4WCghs3AJPY
S+zJEtXVG0wrjAp+ErgRFEXJJyx0uATXIyA+PX1Z6wy9T54zYJ0Zc0HsIXFLrPiS
u95qjdmpuxX9Vx3bVpLQ09vnjbnjovRoQGTKgqPvtl8QUjK0jM2jyzhDEzyrbrMo
f6axc06SAlTC2x0YjFpJaPs06O83ZoVy3O3fEckITHspTvpxUwbZCrHSmm3OOWxF
ZBZO55zjMEjSrop+cOBoYphTkoHfa25/8UIZO3mE2w8YyHA4tTJ8XBuJdu5IfuGF
dePuN7Q+SdEztlbrn/etWfcxTX7ppqr++nb8CRRtykl//6vMJjR/xnUPf+6J/gGM
5oWi2cHcnlYVMVmdC4aLrOj3+EMEXYpAYgs064IfWjRjju1zzPF7lw8/5WQVIgY3
FkWr7TYiCHaVKse634MWYQERgpSMC8JEZPp5IM6TBQcLACzEwg1FgnOkH+rhBRUy
pQ2huh8POhpf/Zv+mpnRmDGiqtsuuoZTkOCGWb2Ss/vqW5bdtf8GSshJAhjEnkvO
cE966qG+DAyXWeFHtRXBhdfcaiAjOksXL3X3wY0aVE9HvIKuovTm2YlkYaRP+h4z
TuNE4AVotfLZJE/izg4cQV6esyElBrNuuXeBfgZiLr71BeE/Vf7HoqBHypFo/CIt
aQXAtHE1TKnkqKDs19/Yq+apXUnWF7Cv81G1uN8dgYLVDoaOJwZh6+l/hLvUfNWJ
ZFBbc92PoacY7ULQi7Qkd4cXJa9FizTbNaIwDHn2TrBQb9JGQY5k1/t+z0mTVYYa
5W8hC/Pxv7IHXdSkwFUuWd4AkEw9dy/3AL86jTLNzTz4gzww6Pjz8n4v4LJD6XAW
98Msskx/DrJReen16oxoq+V1B+/yHyDFntQc7B8lcizDuVVCzQma67anyOR2fMeW
S0RFyWbcX+KEoxIwe1oWAy71tQHANC9rYqSJVNNP3RnkXf6lMbdXAJ2c4IkBRQht
5LxOYScv2hPfXkREoJWuwOsZdFiQZ3sMhJwL/Hs1tk1jkZjvu4cIsGBcO9MqLwXz
dAiuBS2SheQaci0gX8IhqfAPUKN+Lbt5NIiTCof6GoMhYXJjd6dxLCk71zy4Hd5U
4+ZEr0QPIB9KUiYRDjcCXyQ4UbIwtWfzEDSGEmqavjY9hyA2e3xBknkFSiL6dtSG
8buDo+4pwmiwrzb7Y97wo8b+aoglyNW7BH/qjmigiGxyxFbwrTtjaejBHfXbVccs
OtMBzpJRKgLuSJgSJZ2XMWROMPQyTqh4e1JAQJAbzvPQ3vD3T0V42QNxFblsVosv
ExOtWXPcPbphUjwBi25g4mjLsqOpgW7GyE9AUSnwe1nnoRNfGopVsB+OCrHYY+6w
CFVrtlGNIjq179aYl4bHqwDLkPVnNQvOCBmlZmiI7vq6QLcHmLRK3Yciz3jFOkwX
+Jy/99dWG4fwhsqNeoHE6UYq0G+zu6kR1OmfmkbueplxXNfobp1QULfK46Es3/OW
k/X6PrbBtKXcexAWCVw9qqQtZRCKjA5KQocS4udefdLDXbt2qYU/DA3+8giPiLog
nOFfk/4fqo4pdWZpM2FapQOqOmZOXADDUuzoU3Pba6pDCCzAiy38AMWEBc16xR19
MARR3ujXtDzL1gqtui8qrSclGoAPsokK8ABwnWGItQUhXZ9xAzeKgatCda9piY4a
6DzQHAceLjKCNqqVe1r9g0qy6eWdhQdQTs47iSfD48bLvGdshoH0jKR2MaJqkoLY
rkSISk/sxoLCQcfK0+z4nq13+7+/klDrpy1Uzpc8nG29EvjFt2a6j+ebeS9BRIRU
YP5wxkOsHyL6I4n34jKBQ+cUsiNo+t86m1Nt52M37RdgH0pQ1/utnbPhuLhi4TVx
FfFrbhfWCkNWYIM6Qsi0a1d6GobClaQVdq18p7qzWzEYA1xUmO3SBcbWujhEfIaS
vnzEIO2x4hvKUJaexJTfknMNjaiPG9b1+GbyjWST/NgaGAr8/BJBiXtDnpTFs7Mh
7e8DJRezlIi0GDmTFKSuGLrvbzT8aZSm1Hn5dU4KK7f0s0p8Z4RmwrnvlsqprCEc
1+76r2etpaIi76D2BteLHTsve0Xhe+zTpz3TaWct74z/VzmPYFtieRCUo2Zhwj3y
Rl9OV8hizw5sPNgCiT4RdYqFQtgPC7WGWnrkKkt+xbghBwUaLGN/AchiKtDbF7eW
c7irekYP9vSKrZXFX0pzI0ae0TQJyc6wv6Hw4J8fW7fPfiBuFxUgDOqRyeTKn8KT
8AHl3SVK1jJdKKxMUj5RFkwS7Lt6qM5OtGF+yOZopi4+NRlPa3FOJW29NcZxgGIA
JQPifdLpvKVfP5qRRCgLTLaga1bB2Ho0t+W2N16LvKwKV/j2aHaIfo62Oy1k88QO
vGFVPk1eexm7MwKA1h0eKY/uDHxH47aTORByHXUhdOk81yQuwkCCSSJ5W53AYhnD
yCrxiwUNd35YTbKtoMXDqGWdIujtEbZLYLucG8k5GcvG2HDfzZshknjCl4mirm5Z
8fRkVjeoUN0/3N8YarA4S/fSCcE0hP6LuRA0opsG/ZW7Trrbg6PAV7+6u9caitPP
+CADu4Ly7aYZ6MXwsxZmJ4Q3fJWqzqAzluJsYo89bUo6RxvK0yiy1l1Zq2IBp2ux
efjngrfUJV+QjpVAFEZQtitHhsQf4kRYSS1hPo+gMYNufqvcIv1lkFP0x7JIk2aM
Jzbx3UrR9rVsnNrMXUaLof610yEC2VF8dMRgCQKIakXX5PqIcYmOaGTsM3iH4mc2
IPrVIVWKWPTy9pC/7+85sH6tf3JTzhDWwy+Hd+prH1fCPM6dZTWcMCkUfBq0CPCb
Chh0sY62ckHCHRiyQ8uZY/gINKaxmtTU3wyuZlo7ZaImNJEyJB6akzOmQVhOSH8U
zkmcsBeP053k5rLF6B4om+agj0/o8+AkkTLxXx6qKW/l7vahM6wawgkW9/jV29sT
KG3+3vEUGDr+pc0iLTWw30JeksWizPMU+3g6llC5zJyl7k5PIQmpevr7fCX4SKey
R6rGUtvZN4T2I+6D/nqQ9xm+PzW+AVXaXWZLCjD0HnfTaqCF17oXwfrrfsOM5NDz
lhg6PtXu09GDm74N61WZNGmgBaZxzxAoZCp9oOoAVbHRlgQHmzZibn6Vy3bIN8Z6
z3f6LioZS5E3KcpyoHf4lrf5NBcgTOkS48dWplTKwWf89MHqWmwj5zhZgUgiV3T6
hOdnkw0ontDczTF8ud8OoBw3fMQXiGKnlwhGhlJ3ISv3RUUBbmkWB+JBGXSbA5UL
KC0PUmnEqnDi+ySUFzEfecF+kDF2EacVkTxJtqF0G91zWYgq2UMh/S3hIETk2OjS
Jpz8PoTlL7y/TGXfJEk8xAgEGdrcAbA2YicVh5yckxZgWxt+MgbA9Brs2zB2qDbQ
z0wfyYsclyCO9RdG5Rp+SkAidnKwxpImxM03ceXmI8ovRC//gG0sAOHjtrWJ4bN3
9K+1cLZKbwE8jZrvvug7V7+Q8D1ws+J0Ys/9KtrGlxSBGDkeP/nO/7139j9Hp+bj
Iyf7DKpgJRE9cVqcru+PdXdAevXQchIbaYDVxiNsDV2s0eKjOp5v3V8UGSC/rE6y
qIU5fv5vP5tdoTImWPWkWJJbq/Ptvy++eRe+0WUiy2cdt6JjVj39w2RladCBW9z5
x5Hfou8RoZDnEn7rbVqCkAk70NfktCYWAw/woSosBI+QQsLMbtc2wFghW76GFuAS
MfVxUxMgdbp11a+8v/xMEQyycSL3F3w4B9jHg68T/CMKwktg6ynWeg85eDdZb8yy
IxyUiE68BIXTUlnZQj+KK6E4o2OF7X5+g0v2doUXnK5NEXaUQqcQ4cRVM58/TriO
S4Ingz0fcT/g+m/XR6WY4Fu/XfMhIYAcrX7GyMXhlLbtdGY4fAuzG5YMrwXmZQZ9
/xFCMm48lgncP1oK5o3vij0fbBG3xWeWBByh0j1TgWKLoQVBTWwGfyPCqiP+02YE
OA4D89wUJTze9iaaZCxjfdRNohgvcUTVrMaPvB6MAZc6qW6XZV+jNCFB+gYlkcc0
2NBkYb9QMVm3GfpA8Ly6CzygHw1e+kKXmyLpzS1EtyrRWeysmFHXNDEtj0tlEETO
EMM94GtAhnF9NQT1s7iuQzw/RcvIAaBv15LRNlbEgx/ts7NCdjZeStZGhC4ATWNE
ChI0W86Y0ZILeLvGDRMB58+7Itz8S5r2H1DKVC5Sw2O0bc8WgkgTviFJPNyTehrx
3JyBl72s8JV70zCX8wWAjaqo6E+AONwKFMx79VlCA8dJoYMz19dnpZ7CvZaY2jEo
yqtTYBm2IB1y7sD76NvXzQc4zr2sSjagEssiE1tI/p4L1h0obpBUb5HHht2If34B
GBw+hUbCOC40Tp0gzhuhJTyX0L4TyxLTz3gpa4w3mkEenZXfIs6iWe0mZCZOF626
RJFimbxa/seTpkFvANrga5H3AlXwN5iotRYRMynQp/JIdEBvWX8DuI4dIxYcu+jt
6M/nXlE8LeRkqOSaY2V+AM42jfsT1u9t7+77lbHk7uS8e8/5eT5ccK8bPXBjowy6
kP1ByI2KemLGIcF2N8HhV3p7XuQMajJXD/UdMffCxiktC7R27hFrSfyvLrziS9D7
Yczm660gaS+oWIDAD/TEfnS/srXltR0+xtM8YC47hDUFi9psnaxYqNPv1ZS2H079
zDB6BpKf8mMZkxYYJ5YFKp8wtoKILjDmum2KdH6sq520qN0Z+mTkH3BrX8yRmuRW
FbEMj3UDQ1Y5IU8ClbdUhzGcd8enzM9K/V5gpjNitNXPdQaqsfj5HFJpFDWo4IDk
TGD7XLm3hSreOQe7LG6XvR7mecLzBksxvfO2P3PQY8Zg15ED2tZRiuY7OQSrtR+I
vAuP8mu32MAmPydl2sDR+hwd/gkUS+DaDiFoHRfhHiSiagU08Xpdo17CiCgZKUV6
ZIyOdNgIyspXth6wXHgMxIwRrFnDr0KNa/8Wuv0OhzWI70EDW//ZPY6XwayaBsz7
KBaIgmB8w7ubK8UIKlkgG3dN6jsCcN5Ll5qgA/N7CopZk/EyZF0dkq8JJorSlyiL
zB1fnbTual4VWCmmJodlwb1E6zt+fjgTCeaKnMORhftn1FkiTsixCM0XMH+KrTIo
j/VE3cabzyQ6XjSRhUyn8nli3PohcbtFhRVSfKPzb9L7Lhq+lVQx8ms83ph/HlPM
HFCirgnV/utdWFao8I8RQWHL53lKX163paJUIcivgAs2dWUIt4IAhLkOo0GTKV04
15+xVbqfDBlKbM+GYKNzHjzFuMekbmcXDhd6OBw/BTAG+015BakCtY8NVPyT9s0P
B9w7zlubysgnSzg26uA1geRWJHRMecsN56rjTnuuMYyqyjKNaETxk02FbGRYIL7K
RZEbQKU2DgLs9/CLvAjNUrGzTTUaHmPuMEkow34NppyIf3yEvQNDa8Pbx9zdDP7e
Q9NlWnJIpgfd7AugjJWGDVSZeXlq3nlPK7NendXjVewg3rMmwhMlHGiD82RjJmrU
M387BDDAQODLhGvkNls+XlK+LwXv2izSmA9rdHk50yhDGzsVdAlwWsbVvSL5RPdc
/GWXPFsATgUK9HdMEBIqiwVQuUxsGOuQ5E4WBicSBhhbPiidZJ5BzToweqoZ4Lib
FsXl6shLGI/b1WWnmllh4A+FhG+6r74BuR4AqSUXarAxKtrPHDjfXUB02+MlG3Bs
fZbe57OzSySbSbICkzrL+NxC5KqCaMV/lLdD/prPjtCJ3YyUJstZw3vfqkHoJez/
e+DnUjnkhv3BDLb4zYs+OaPxwrGts17H53jR+DyqTcptpzazH90m658B081WIYzM
mtNV74y+C1u5JAsmMml4WKGxFpYLCnCSbBu0rFSEBKrPsJjwhSKhnvxkQOVJwqEp
ej9VXiU2mWItjUCq/ZNgcbXczYliizV8kgILIPwGskHyJpunY6MWwoqQojPbWwzR
n3Aq2ElpQCr7zKfDN92UDINaO3BXevUck/RWWaozytFYw/B82fKOUhP+x7IokpiX
xAIJmJFf8gEszM9bQLfi1kGqo9nypH3KA4Usa3oAtDLucm29LtGSrIXzxucwJpUA
3vQaS+fFmYGPRKaiCsXEBa93rI9zkoS4WwSyjgp6iZkEJnkakRvZ8fSXN21eH8+f
IuCn1ubicu4kBBCjTH6W6xxjs8lYIHqcCp9AhDG1hfIlEjZuHmZUIwErnMmOBXkL
m3srOwbt8skgM/DJa7hWXE+u/O62RNhVqCKShY6wYwyTisYm9pLj7oEACSF4BpDa
SlH3Xd2cPWCZiLGVPGKmdS9agPrnkuWkakd9s/ReijkkF/6+iGK29yyBcgGzU7tN
ZAqbd2YknJGb2Y4fxoySvXRdLmJ/r0XvtZ7xa6/7D8sIfiUOPeA33+L5nA9Toacn
MqvVeY5zjkPBI/Iqy1Rtxb8RClsym4rhRUAJ540Rwd6AMCN/4AChiiudwaHNQUOQ
88sbDnEe7AmtHDAVF4tegpdoX+nLnyf5Q20KzN8pHcffqr2sKORiCDSiTkLVkJYn
UHemXqr2Hdfux2jLgwqMGOxbLivPhfmpdGxFi8O8KVFemokPdBaB+PwK3YGdYGRn
nQ32fmG1hGtNiDxSWWxFK5dIwbBoAlQdrNkiHKV7vhs8lwv/WE/Jubc+vowB6vhX
B2tNJFVt5+4i7vkCOfgQ5a/TbmdhxEHoQBOKdLqRDGpDcMCJ3WkjMU75Adb8Y89/
vUI6WFn5Yo5PzvteFndqTkuDWvvXMavaJKe5AbGbjzzEGCkJDGFx6eRzvDLJ3Xlp
fFNPCViCJRtp1rlnpaOGmarPnNz6miCiPf80Bprl2vlQQMCNeMKPIX2RXr2x4DOm
q0Ombx42q7NjBt8AgJ+soTgcbzEhYYaRBd8lsgB86JmJbpULTWrW+JkMwTq30pVs
28WlKzm5pPc3lNnnHte2s9FFP539qzIUPCalZd8E+eLPC6b9WUcpc7wtGCSRUblM
7cbv5AQn03q/DJkuHo6S6K/E29FbKRhtjzMMoWwZO9+f6UurvN6vUqvtoxaJ6JW8
j1aCRrmAs5h+NDfnC+rTSQ8kDuvC/c9SQ36KbtKA/H2+64TZoderHOyqEsVm/SyP
McaMIh6G6SUoXdillc2erUmr9xv2N+uFkC9msHx7mSIRyxDR8z8ov39q6Jw/ayff
+IU5PPCryDVV4WgFl4bSA6eIds2/cOR5L9qNTW6EQGhK64Cm6r4iU/TqAB05lHnO
ASpXLO6bdvz06p+2UIv0Eft2/S1a71GJlXCxcdyVc4RWkwiZ/MG9qBVeN0ivk1iS
xDA4ZEvzA4AJFDQhdWfYs3AzJx0AzRDLjaALA/LTHfKQ7X18oHoLU9tt/AJdWFuX
RIa7vCOp2y2udM14JDcV+mm22cTU1+pJqWPHdY50ANnt55EUAZ0chGfMmbpiC5BP
2WShqlpu4sahKFbhFjYUoNQ6SArUIuB6xjqX4+yea4BN+X0BCMMrTIL1Ung8aOTI
BcUvrZRzPlunFrfSw45v67EgJ2shBju6wmS2m3NN5e5smLtFAzl3QCOcNCV+3ZHp
WqPJmNIfjbVUtJeZwccoAfY0IlN9ONm5hVfJfvdFswoYI9GXHVOzw8b8D/7sS7my
TQCHiQQXK0YOFZ/iws9sLElS5tmRgFfMvFjayjPTyUdOa40tKMrWKp8Wdc2GwD9v
TKimZJnq9VHGuXgbKgtA96LHIGrgGrd8RWuDiqpc5h1wgtXcQnMgH2ant7Na5Rhe
I1Iq7y80oRNRY45NPuKKP4cWP+7JFMsYVgdqD143+6zuLuLOxswyjd9y6P9NtXto
GWaPB5/wephsAYYqXaUvLYFjDGIX4VidLnAGEstM1QpPi2xQTFBb1GggVbNSTsMC
wkvJ0n7XVybU6eumzH9wgk7FYVM3NV+/qoeE6QoN3lr7GqAnPqwuqDVqOajLyOnt
8GAGIWSTwgdEAvm6F/6FiauvCCavGU1xFTnJRhle1N2Uq6nr98H3v9dF17h0SnIl
T3uCEUiosbC3yzWF3aodgrPRPYX5HNQHFbbSztiJSla5oAV28bn4YRVK0am4Y7x4
/JsfyMKIM2MnsR+yr7nW95bi4pVxwR5ZKc0uCnSEeS1Rf63dIDiHbAdbp1UGoT3z
GuS98zQTd34h+JOZCjs207UYxCSse9wSgHQ+H143OKqQ18MpUwlUrPnDIJ57XSWP
McssvlPHojelvJ73XLHD3+tKGa2wFh3SKqz4wGsMZk9dYyafDa3TBXKFdPG3Wlba
y4jcCkMjPiP7WCaxghBLgkL0g9RtT+Kj8P9FlHQqN4g+Wz/evZ5bOMKn0fZE+DBr
Z5MoASBQoQohfXdfW7Oca5Su76bK/ATJS9koLl1MFakIsQn6jCj+CH35KxVfM+7e
9iksn20rIZqaK4Q9XbouKB7gefT4t8BZWezg3fBWxRJJY7o3vJgaPoAdibLXTVDq
Y9fR5HfiH0Tt67yzcJy7i4WRKSLz2jw+pW4djtQist5lwUd6uhIqlnegJ2OnQmFX
ubO1b4ocwr8idodfrifvQxFt8Wnn9Rc3bxD6tdQ+nQwU4NvMMBtLhdrITEp2M0J0
KIpYySbOkQmUiAK0twK47dlej+cHY59E3diWmj72d5QUo1Q/6YlC1f6ZNDrkWbDA
wnem+Dw6vW+nIc3ElZ6ibj9VREIxzShACG7MZHz/UpsW3u4b8sf8FY/cOv44k0el
l89w5Emvwer5Cfq5qPcXhaf+dULDSmHxrJwFdY4AOhZQ+MQUHPCMjLATbfTsr3QD
P6PmGmziXW5Do9Cm9kWRqdiD9pp6YPVgOZ78vgU+4XQ87ADRzFKbWiw/iM332X/b
lru0bo8iXydfG4FaooaD8Ytlc3b5jLdu/HLULuIw65khopNscRMeOnEFLnXeCx1l
8PZNfh5vidy+x5bwl0KZMaQprO/CkxQH8Qdd15gK6mTw/6Ujn/NcEulp7I99i2Nq
If8dnVY9yHizyvujkIypQVyOBw+GcuxOXTDwYqL+qNyedF7Rfhgdkh9tIlAdkWmv
4tD738JAVhlK+xz1HRSTWVAmnItriVg9CDjydpHWfluEi2zzOsgI1rkWAS7HpsMd
f2ebyEH5e8HiQ/4viu2UKcPW8ps5sUFBqwUZzKngr9nWSYWbU4hLcaR8tCS64ljG
nRsRT5shhOWndNLecUh4Pe9coSA6sGvIfZfPAOm+2tzr/VZLP05azAGz/Pi6mnnx
psG738qfTAwiy5kyQ/O7MVsXRRZWpksuNBiaOtsxrF4RloNS1z4VLsmFVMn+D1d2
Sk5sjb5BsvmhkVnnpGcq48XXxMRQ+Px76D0CLMAmm0pdabT8K95cIsRWioa34L1o
kaJJgTFjvweAFt3HhbmMYlLrvCPknc7V1Kb1xRKIQZ30HcxD5RSLWU3vMv+jvv+F
dPdVnZdbBwLHx6ddHEAH4nOvFZmYYCjCBG90rt0P3Kq5LpPt+M5j4+/uxAUb+5hN
5USjLP98J8K+6Gg5BorTWT+Z5SaMGHxn3GQTOBPFSv8MIHC42v/+l/vJ+JsQdYgV
LPxunlnS/TUdIdp05OB+9rd+G7XxsQKHPrOrJd2/uhsnxO1l8nR5Bg0+3Z7ZFvLD
AemXhxsq9bJhd6rpzo3lQNVCijmG52/2YPsKBQcngC1mxEZQKjTyfgoxMCU44Ycg
eRNzJp31XcsPrRzG++jgaJZjQCOQ6v7yS0jKj4ZLdZ7kkT6e/76wCBBVgx3U/QEz
JT9GTcPXUl6MIdFIs7pjCNpolAUf/TS9QbiYEW0M/YSdeW0+zoUy2G270kcjNnZJ
xoO7zAFRFfemHeJNUzl+eVjxre3WV/7WgvrXsel442VG/7Wuo+fLlFhuRFak7Z7V
ICgupQ04249IDTK2S5hd+v0Pl457TAEs+5ceuv8XaJqye3x21uYUAK51a1Ce4e1R
eMO+6pLhwm/qI+qzQpTuO2aqWB2OSBtLrlnEh5MANEPELNZVwJ8HaVvQ/a4ngc14
4WdKu34OyK0zIU3SMOPKNZBsgJtdmCGVUOO0cNoGNBpHYXABdVH88Q220PN7ao4G
mg8AzF8+4Jq8g59a63Tc7+93meBMNqWDK9DKaVqoCpWqjqb+ntzwxsGFIWG+BBnY
/y2+4+BFT1JJP8lERmGGvSdwSdEQ8cCgRlYQnSfJ1OzDBUGezqauvmoccv4uU9tG
w1FkM8BDm4QKX0k9CQXbdQtKv1PsBMdMbEsL6Chjk7Ewpo8iNt8MLJv0C5MMvHtG
Spcx/UHX4NAxO3Bg55VGyPSDYVsNAN6jCRAdMLf552PjATK8lUAiYLSNoXl0ck7V
zkxPLRFHyOTcZotu/vlhPtMFo0h7xj1RQk2U1TcsBtg/pIB7TKONkrKrmb8R9lPh
17VjkIm8/f3ROn10VpAK//1eyjSy0SRi5wpX1DXWVktDgJvwPedyh7X7UbT0osuh
hRHPp94fS4zRTQxr+aSkzizhTnYOKvdRFVrjh18urDRkP5BYhUlojkvTX9il5k/s
oi3o3GBYtfVvAfaSvlYXSXPW+0z7F/fPXU7qHzaICe8oBDbinBO+hGEjYSAJ3D4K
ar895sieuf9gaWm2nGDgrDEKpUrmxjDas5TSxETFu/QdbS1omko1kqQCk7firtaV
L7Zcg165J1FPxdjJ9hzot4O4MCFkCqez8bEVTe6+mlptvqmSvw8S5uB30nebPtlt
eyaDM3NvWlErH49lbX+v4TMJcFHb0rivueQlXr/cIHeJhGAMqihL9rhl1OE0Ymeb
1t+q6J4YhU+soTkKI5a+I+KqKbltS2rObIvTGEgQvIYQ7sqszRUTQRYX38MLABAw
UjMTSbUJWGmQjmSUgcpW5E4nfgtNFCr7W8XbevecFbtF0JQ2IrKhgyYC/yiU2a5/
LYhKHvhNHoOSJkcro2Zylim06gMs5gedcOfv2g+D2FeoPeW3fWe4Rb7fTC9splu6
GDda0DoGC0KLjrSQYGVg9lHIoQm8QyNoml80v405vIOcOMlM6CGbNtkQDr0zfqBl
M5Fux60Hlkvn83+2WtGOlL7CeswZ4p69P4LdjInJujlrgCTiyAFLKzYL+QDM9DMU
vJLDTAq/6L5FIOZA/AoCdXCYtaKwNnzsnoNLhcF18lt0wD+2qG/D0xRZCtWcHsG1
dCy+NI64fvzFIloD9tHuauKi3GI985cM3OmexZ2Kak7YLLsmrmXAV3l51+aFvThk
C/dTEMZlAWhR8xtqoAgNdY+Y/UJBTHRapR8DNhowSYyqvSaJmUyk/GpE3Qx0xzxF
B8ISAdTgFUONK3iaGOL5R5WtNJolWY4KhTRm7c9ga4/K2iLlNRSLpE50dTbq+SKg
0NNjtwf2vujkWuifLAGl6A8lGXKLNR4q7J7vpc4mjVM1nL/U7cDlHXPQs5P98qcG
PHMnYfRNwcaQ8UVy0SSz4Sz+/LgSxxD3CxtygUiM+dLlF0d/J0h6CifQblnf36wm
v46gqPhHCVKKjlgs0E7mJa+4shF0Pay42kw8adDqjpUl724omJehE4M1TUYSzyOD
scBwO8x/94DYdNZyJhYLSqC2wrdMynfySoeLv9c/kdsY0EfwP6JZkc/BvOHAQgpv
pSxr7cwU+aypcFSP8fKNb+uwSsVDoPvSkoO1I/GJSb7R4CbTVfQzmf6Gi07xESQU
qqIAfG/ODqZbpTQgTp/Tep/zSTKfGH1j7bj3+VEP6eBMoVVu08w41MaXwQe6vmSF
6d4FV9l2gbEPigLpLesmBQ/cBAcFJVOt7ofqmnC8m4DhTApcFlkQHePOwXXztQRk
1P/H96mLDKr0k5w9mG6757YFuUCIZ+4ocC2eDmHjN0LGDVG7akpVqc4yOOSRSg3k
qnR9QMne7MHIGz/Aq046tLxUXUmz7JRdrD1womyFS1KWtyIs4ZGEXisuSHAz7Ip/
GnrYTL9INZ4TeFitHWAkve+dpf76uAai+K3h5zxlh5u9MFKW6AHsrbN42TZxbfRC
xUldaFqu4A9yBk/KT8LT144rjrhTtIAMFgdYsuUaKVRF1zarS5bjsVtR5re1hefh
HZlwyrowjSXU+pslOapFHW66ZlZjYezhkwriApggzAkJdkFJj+4zG1fPfP+bA8T6
/QcIxt9LOq1L/9+aobsNkVyawxwl5PcpVHEH5wg8stlzWs+o5jo2c2wbohwWd6hO
z1o92o1PWggO9a/D0ui1K73sXZ9aSe33zHibnmMiy0/9DdJHxKogpWrH2Qd4gnwq
/uDPMMcTXj6gJAFptVbl4CRh0NjNYcdph6veHhZWtkYHzx+AqjG7WKasXcaXfjJm
dxEYp/99hR3+aX36oRKQmpJpVNMu1xXYNS+VD1bkRTNPtFQM1dO49GUIw8WUm4bf
k9CiigJnTy8cPQr6IvyuaYXlX4neUD9ARuGt/4Ay+92qIc8iVSBvQ0IsThy8uZLI
VCTL7RWN9Ts4xq7fVj/jZ8bH0sIle6/lcZjExJrFZfB0RwgAOjc6Ih8vptPfBpHj
Tbh+Cm0FPPQQr9hE9R/pA4A0ptajF8X0ufOj+EUZfNDJZ0sIaQOsKh7oSoBWhhJ9
fWkC/BWDOQTaFDwz1IHgnCvTx4QbPpA3XsqVwhuTYTsIN1sTSchMS1FjaNM9TaOS
vPwOxRvL6Sd9pH8R+urUeHuZeNQmRzZYFUWfHdQ2Keh/vQuMAXDLw5XFYRlsGbmW
0Pi8SqE+KlvhD3VWLBScbNlius+zWSdzP6MIPceuG0OzXorn3kw/bwOZ6LdaGeyO
4dGuS342grpCX5H0pGCxdmp8BwfG+3GX2EtGRSsBn7zi4011NKk2UY9VIfYzjQsK
AOuDKoqMdrus6Ye3CYmvRXaHYiZUoWOiMnYEZBvdxXBNB2zRGYkxc9NFoCDlgrIp
fNlakstzcmtSdBu2enqNx3Pq+3eJBmqjg5yxqKXyl8GWkNMQtKjV/r72LnD84T9w
60WkPWoZkXbeJhLioEeO4sMDMR3yykzsTaFt0BU2DfukYmRXzwTkMsBNNdx+5hvq
ntpzXjX18MGON85MDUUegfV7kf672I6rmTYnj+XdeHXBLXcJ2KYig52w4a6Nwn4X
d+l0KMeg5Sl0zNIr5et8fcy5Qmpy0w3KfcndWyxqQoRBqB5e5RJ51a47vpWcBw75
k6F+ZQ0f2xXoEgHCXgYVYaR6Gt73LUW+bX9g+a1xOjuvi7AhpMfkBhyQL7LYKrmH
uAY/3Ubv18knF7budJYrw0zmZe5dVemFWN6s9awoppX/1ljJ7OtZoBKdEkhX2l4f
f0q32r/TAn+peSUy+SBmX9fmwwURSiU94WNHQfPldwOuor4qpM7fo1h5z8eejBPi
bvZ5JFilE8N6QAP0HBaqfbNGzrfMmyyZT2XCpiVhGATqPhj143CBhRyw66lik/Uw
ZPD+lHHbfCJzQdKMMuO+VTAEc/1YlCveDOiVt1yo+N96JdxyKGv/YTze1GowtHPP
65xGM8BxwDS53Je3ZTdFnAUuYDS2BT3/qW95I0Y7y8wiyub4grgWsKqEde/W+Lp3
uKztNzM3XWKDYCiE7jrqFvjA58Nkka/ZsHJuFjFSNmJdAYGDu1f2jA0/ZA1IYff+
q/eI8Rn4UDtHTM0PkBNheuTRfk0K7KmigUmQr1goYg3tBMdRSb1YB27r+654UIoZ
YC+DIryGGyMslehpk68bmgOyEbaCrgPhaM9rV3VXDmbKwNWrKyyu5GzS5/lBCchb
tqqxDB6WZzx/x1dVhdyHJUU2alH/lASBT6Ov3bXaSapBz/8hHM/GFqjxb2+W5daH
RCXLts+i6yzppTq1br3BhJaf/Jg0/y21jKY8lpZP+Ntnqu1rWwoURcRaUOSq8aDU
82QuNqSzJQ8+WbLJOsXXPG1sRF4c+whsPtaGEhqU7pXvLM84q224P72vglyAQaAM
2DbIvV5jOPJgOWv3iZ/j8jX524p6UylFP67jF24PfAe736B6l4soWE+dblxmvJsX
hBY73nK9Xtalw18NRplKkMoLyn8XfchqcZHy76N7Iyd8qkl1N2Ky4sYwpZhIL4ra
36kiTMlIScEE75SBFoM2Ui+Y7Mu5X5G7UFqml8AoPIoOvNTEebEn3aM5AfVa+XBQ
h4dPY1BmoOHuyTVukw4/sL+CE42xgE3fO+iTgBMTHbM3P/b5bxDjqUp/CTuPDaVA
cV8P/n9U00ZV0sLnKgVPOvoHMzOyP3kCz8Gcdg6+nxVB6uhDshTEWsXEVyp3YNNp
tGbAy79LFTOdjoFyEj1cvrMAGLrsw46ZqxPQ5EKPOPkXULHWF7nIvo5YotDKz7Rx
i9ivelezvYG38TByRhfL9dDFHjfcEVVgsQj7sj6d9oiNrMS891DIuAYYAPY3KITg
DgOkLFYz/6Q1IC0LoY7lKpH6qqZsGX2qG5kw4rlXg1FO22xR3X7ijj0Mo4AAccm9
dDNnmGRfdNlZcNGgazO5E6UgyktTxkPXalNDY9qx1EeQa8tK/om+c8O/Uh63qt46
WUrmwIa83ln2OwcdME0ukAsj6OoiD0eO9Im1FAx58IliEqmXE0zy+aBIRkkpHDsA
QUi4SyYj202UivEZsfiUkafpe/i648aqO5k0Xt7yCq1CApRYScw6lJ+WhdvRMev2
e/g00CNsLD9qTGLm6TDydSI1YMMwqEHG0NR/tJwreZmfyfmDDz3w5nVFTk7K3r6B
JNawasig2dt2a6TBGsj8cr81qVLdEeStObhQ47nMpQ4HobCCFBxvIR+p3GYpMCV1
0kuepGQFwCtjoXNVZXk7cxpZSfaR1BUywAbT2eVD2m/uim0jhv33A3Afm3QzWbU6
48UWxbNPm/KTmZPqcASxpwu2yD7R1k3bUVgISvHBCMOvk3+siuC5HRhoRDc3FkLq
pMrQNk0QLO5sLN2kDnY+rwWw9AJmIoLQBh5GyeF6Wp0y0hWQHx7KZwoRqKLAew0+
r0NXjfIPfmIG4rZMU11yebHUJRfm2NnR9JJX9jIJLLxXsqF7a+rlhMEvqnzOUoca
GPg3jsThbonP8eLyik0Zk7rtfDtCt0CG3zJHOdJmImOfqYKikagBEVR6aBuWmSIp
5ez8K3NYbEcYH+NbTXD3359xGwTSC7ie8P0n4X6H76ZCBC0/LZ+FOFecCphABN4L
Vck5q+JGBw9AahUUMTW91xw5AKL46r3VIpig2qfnFNVcS7kiPf/IgbkjizkjNdL8
WQSDxM9u31ESEKutaqiNOm84qO1qiiOW79QRrJCQ+Iv2saXZdiFJxhC69YCC8vDy
AieuTE9JhAu9LAzahFuNM4WamDoCnHT3XaDxFe4szUihYAdv2KFvtO27p+hk0YrB
XABwPD2g9kYmpiSVM3wL14kgBazUKcovqbnw8TYAd1T4odKUZbpsEn5X3/8Rz2KM
6F+KzaIhn9xv3uvtw4IiyzTHPU6KaTSGlvV//qJjSkL0yWDjPAP70vJAMvh97SMA
B+DqzjIf585HXHoxW4B7uJcbgWfMaQXeLaS3vA/I21T9GgqmGvqp6lw3Cbky0VWM
79i4bHdQZ+NSyfAv34JV1ZIizEXzSxtnPpZmWnwDfuCM49mjfNKE3QHIW5ZbfLql
nw4LoaT8opyVUX16t8LvDmaa73pTO67Tz15QWR+UbQlDtNE9fJQIjcJg83Ge/OyT
152pBDKxUfzGL0iK8lwFDK7a9gaBP/E0pHu6LeMvDKTVsFBOH49vReRMo+jyUQDJ
ebGo98UXyCq7uEefZTJ3QyTFwv5hACXu3PufK1G50h4+5qSAl3VlJQbsu3GUpimF
47IwIg1zLrNvBVUSueRSqMP2kM5+IR4yq3G4SuiFTnOSLgUHAZEv0MHB5HNj8Pe6
BZ7mAES7T8UkfN5yfe8XhwHuxjRk8MQeovYAMf3LqByoi+oNLJcjekp9nIVTBnFL
Dyk+D8yUzr3tov4Z9gQ+PHPY2qTcpCaWyo9qzQ+NTIiNFO0dLj8TDj0yckPdsBD0
/oGhZ/SeniYEtGgzlKqQjgkIXoRaNnYzS+Vme+BY1MJl3jwqfjBmP21Bq6f143uM
WM87miKITH5T2K8LAFlsi1rsneO7FxkJHOxtp3yiSv0g7wiHIzqj3ganRQkcHm/C
x9F34NmEFw655x2pq/bqsbHWqX5e7s/1kXQGD0RtGaAiutProm+yTjUq8PYqdBye
Dbd7/EjC+WF215pME6iOalQSOJTNshlRGtM63yws20p0VI7yfJAkOfnGiDYywBXm
NxfgTOJyjN7YZ9szsGPYVFx1vDq0XaFFDaJ9zg3Yn0a/Pm9BY0vJWzIqJXwnvvWD
1nohcixF3RNJYF4iv/KtL/XakM9vtSQyA2CRS5Cq6N9aYPDfTBTgwldL8kGTvujP
sUHL9akfqKRAHbFF6GcsaU9kjHqNWumOolibW1/C2UcQGjj/dS1RWUE+Sag61I2H
ZDxPfcOpmQ1qIiArdBqXjehwRrKizvV3bpSofXQlOGMZhoyuTaLNh6h7HNJUjumc
pMYpf73xlmsU7se9KvgJ99rOyxLD3Gt3iYqrWrh1IjL+nsg1GYFz8Wx2911MKThe
TBYBqJkvY/Tdas7PyHZAQw7QqRqsGq6iisKMSBDb85NG7KEpnxNKCH6Yl1qOu3RA
mzcSubPbSBjrw6ntZfXR3qM0GOinZOg86V/aA6XcWDz/R5z9Zfyx0JAhTDUlgltC
fh9q9hrwwyGszhnbAsuZBnlGDKLoq5/JPyo5qnP0HYPtPNR0Vr+L9rVWEP71Ynso
RlVx2P218gOSr/4XkfKiLqvT4pUbxoqvS6odW0fOPSyNRzmixrRQOqb8JNLgEoR2
LW+ir5ViNQrn/sXbAV4DPqNpvEwLT2K3tLUO+BjckQ/zYEr1tsSkFvmteKupeaUj
rROvDB0GefIgWRPxNP31XYtutA/4l3bfMIHk/2v9IQfvUPwzmCLIw+IFALRse+j1
2N7metzFsjbHe/nYrRPRkBJ9XIYNb9LMeDn3CY19tIOXYhK3keUNb6ZK0Stnj1TK
dqQFKcZhROdIi6xjgvVNiigQnsItQLbc+x8rPnRG16SB+dl5llSgVkVbYtkRkKlY
V7wvLupLRbmoeUdWqMY4m+20zD8VJUwN1dGE8p3g5tlrpKIpyscE/MsZhm4MjffA
qOn2WIs95JLRRuSPa8M5k+Gezla/3QPuj5INXgcO1/uJiaYt8O5RVS/PdiRwXIly
FuKmQCogTlH3EGiakGAqTYC4dW1siHVRaUj8xW+a5NUNquBuDcRxQbtqPKkuiv46
ITn+3vEJKHUIwByxYTR3iEn+aSB9hAMyy/l+vx6AaXOc6a0pgxm9A8DAC2LvlXp6
GAWTckqhDbTMpesPfQhKA42n8XEeHb34+uoH5WnNhIptzNmLC50iIjvuHFlrmIt1
BY69+TrbmdbUziPyLToH3RCZy2yH0IGVcaq+1OnKPdANvkfn/CZPXKcY3kf0VULP
QRbLkvC6HdmPV4tlUzWnZPeqxxDvfU5eaZSE51LLS+oWTrtLZz2+axab5/bIE7UG
nMYuBH14iIEblAItWbK94cvLN0hVD+7kPlp3773YuRaXjSxAA3z6MGAE6SyQBBKl
CNT2A8n28gJ5cCq4C/CHMAgyePLzfJZPvl/wsrquhIjNO2bFSTNUd8HI8yBGC5Kt
TtNLxI7sp7DcpPcTHFysAhe6VPB/sLOa8QMIpK07CXclTJEwsrgx7UQnl2pNw5LF
oquPrW4QXGDLlM2XOy1im3+kTLJOIjwU0Beuu1ed9EPXlFYsEfQJ1wtcE3WR5R75
llkPB206J4ZLNFlKhq5Iuz8jpE/DLwMkdFzcq66OlwYm9/CCS+zHZTBnB9FhzgLN
rHjUWCgQspnzladfOKAotR7Ak2KtVltYwFCnTPj03vqQKznxr6AAVbQNUL0pGXQa
26vzSYXKSgRS90QusIJsaVhp2w4f4o5flDHxvFbaozbqsdPyQOEcWORUJG7+27Lr
ED2wfwD5oGwGYBBds4ZwV494XdC6FJlttTjkbs6Cb0FAUxQjDOym6OMghDWOaACn
Y+CxLUcKnLJ605OpEV6522uchVh6IQO8ojAQWsWBYZIrYFH77TtaXeL7nW30F6Dr
RY+13989O26rwA1GupNETOoAby9MG/7AzQl1jar0To2XlfvVHDFrQ/PFk1sftCbe
QkXRK0FBUjXQ8AvuYr+W9dgySNaojsKKmyjRS0RN605McMsAIKOUbE1w9MVvEiAv
8Rg0+ttvCSPGFllBaOnzM1s2UW1QYFgniQ819gIBfIy8HIxCmGbSvS0qMHQgB8Ww
wiNWOUvvs/RVH99pJ6ydn752rgBcUWH/cWMEAJzaXYkldaIk5OrBs9Bskrc77wEl
DGsX6iGjyX3DJXLOTd34GiSaTgMFHJY+uxltnufMMvD+DCAuNCMV8IaYA3zFsGn5
0Hh46ztqz6t3AypwQUmnsIJkaw5f7QeEF33KFoEXk2eDuBOXm6iCB5CzlK2UgWcB
2/+KRL5XtrEBbyxWIixIOELxTQz1r5m9mgsACCI6aZwvjB0P9IJMf0do0SA1YM7g
gBZJ4ttTJmerdNA4+oF7zgdR415OnRIcC0o2AZL01Ie+oXgXdqqDUAMwBLLe1sl2
Xua2e8r0OMTYRAS8YAz0PHkDzG+wLYJTy/vJmCayU3MdhDRHVrz7qzZN38I+BpJD
TFFt81rQ0F0uhwCuT99T9ctjYshH/oirO878nMisf2g6wOHOo+4O3LUt0NefEZdA
eviFmsOfMkaoxF1Mb10sXSNaHjTWwpqpjyUrMfT2GCI7EHv8RWzsiRrQPgFiliOB
+UUizH3QYYlbYVPAV26jRk4NdgG2dWMkPhkGlC8OhdGBVNRfF51OovwnGDLtUgkx
aUCa+6S0CPexgMiwYmoVGR+YTZPBTiiMvRJ7bQiFICWOXUhOnJ+xkalLLEfGs6Ve
T/WA0ivPvu6LQOaOtYgUIGF956X+yZJbRjH5/JzDWmTSVCLomZNRW7hCdL3n+RH1
TQBG3jxfFq64EW1hHjArJE2bV4aku2ZSk9XevAq9tjR3BmOMES6m3sL20oVX1k9c
B3IZHeL8WBE471JXE4oa6jw3g94LkK18PUtgfI9eVTLp6P5sGhfEJHFBRW9Hd/Kt
qBJO7oYUP0GgudyuL01PuRo09jx6epkcLKziawVc3W8N+OoHNbp/r8LQIcrnAK8r
oJAa98+DOydhLxxr9qrBT3VaNI+v4J+q8WjysVkgGa9lq+itRspQ3aEW3rfypBBo
sylY7eRpQTVvObHNlTUNpEyQXqx8W4w+2r5P99oKppMT3GPZWhdbmbs1in+W2hzo
DK5cjVzoG/9cQ2C6k7Gt//qMlKbgJR/w3+RqBXKrZQQYliC2ZsUDGl7eb+ji0bjS
5YxfhqjAxUA5bvP8yaFT+/BaAEhhGQz09/Pm4y1LOJCgcN7XaPGcY+SvCUIEpKHu
Z2E4zxIABKBiDNg8OILfkL9wW3joztlY2WToB0P2WuMiPHMOjkilgZMTUXWsND7H
MOTDowNA9wlDcmO1I8LQxnKBkOaq32GvO2qMW7GIB5/+g+sVEF9kE1owXS8bTbt0
LEQ9WWGXRUmiVfF18ymnruO/uM9L3JnJwnxJffOQH1rR1a4gpmZeiqGugaLkMMjk
3sxniHqlEH1+jEG5Gnay8Jv9rrqelC4WUADCr2akAT+yKVYYtjsIrZoyd+2CIAgo
M38+EubWoHOtv1EBGj8LgjD/pOlL+ThIbF1eGWjtxAifczX3EiuqcK6bEkItpRfJ
2Y9S7aTFkkh/6TGqK8nKClhAkkgBv96zB9EJBiWWz6cymmF6QwxK5wGMGdQnjA1J
DjsZk38iAGVAzeG9JKqeXMW8eq+SPk7Z2/qn9uF00JqSn1oOA9VMyKkYJqeemwEa
ri08M1u/N1jf+Sji4jsxu/vNkPeHsqsoSgD9RSAQOuYvPiN0tkB+l/cYYwKlPXCj
1LsCX8GeZi8gAg6yjcGyNvSRrXVPeFtMqNFg/NZhfiuGvdin4YCG9o79k5WtfNTM
tSh8ph4AUG63SE9LTzg9hCLkst1l5YhqD0kkzCmQZUyg0shHOXZ66aCqfx7pJajp
lneEUweHRW63suMYyM8fkLJ2zXhitZqcgbnNmlEITy55Pwx2PUVH5+IL0oY8chXr
QDGaOIfhmq33VxYG9Ga0sGJ1SDlwJfHJnNJQTLMGjphk8e0gF3/gtrAH8DC5K2Sw
xw1bEXyJtesB2ejRP9Shv4P4jQPvWfVMQm/zO8wAcLQINM9vh1Z39X+QlAu95sEb
0WVopOv7qvaanZM8KLOoFqL3tC0uBXbNKc22eD3UGrglLgzvUeJ7zemx+DnckUNl
MCLIaInhIy/rpvARzWGehgoQo2jCO9hnejyMgVsSj4uPj8Q/+p2mYFU+3cXCsS5Z
KXSAYL9HLuhd1skD3CYSgZaMw9/SwMbxo9lJW9+BNKlxw3SvEU+k/fCLylQsNWxp
6xPIaYpqISsJP44CmZupkpXWLIMdegauX6Vw+Z186c9TP2atjRfd5IK9EAQEoRAm
AOSTXz8rPP8qHOUMgr2B8Lgcm8+rMq+zAaEiqNOwTHnBOdoUjdpJd3ga5xg0l4w8
JpSeN9k/irrh+/WDLbmZb9eiB91CPkVA26epjOCyZuzWFLKnNPLvTw8r50EdFxAc
aZ1sM61kmsKeXX/o7AXk8OZJ05L7JYBdKqunT7lAAAJ6KgkfP6gji1rQ60etgQxV
kf6fR2SKgyZaDVwBwKLNJSwdKD8KNpD2X7lDiOes7nzPYFRaeGnLIe8gJ72oO5x6
kvDzqYuoq+ZzwxVFpVfoj/re0BTsnyWGSDEjbhjeHa1jd0eKoaNEZhS/cdcQP5qj
sIwQ5s4sxRBv2nv0ghmx+QFOF7GRYIsQBK0J1H3Sc/E/znVyg6nDdQL9xs4Kdgc4
6kt6gUaeezm5yRo7OUCRJ0LymzXWfiQ5fzquqBl+8BAxsnyZPs2qlirmRRGkO1Ee
ddINuhhGKpW5M964RmY0ESg8xXPPcKk9AjXMPe8aPXr0WasFiHBdrs01QquXPw1m
2FgemvXxsBvYYUn8cPQgHzTgXd4h2bnUS71SP8RAiY/gu0lomSqh5BUHwaR7ngCN
q6/AJFt8ojhfHzlBn5P/qXUl3dx9154WtuVoaO/CpjqKzv3ChH6h/xBR50FxOq2i
PZ/vLOpMzjZWoTVlh0fjWEjIr1YTlJo1qOFds5I2VzDbMg74HfcVFLE8zxJWYVBv
kApgdHZ9wNGCfDJpbtWn14dsdr9p2FLa9sUkOJit2cGN0NHfwhLzGLA5eNvdpagO
Cm5OmQEx7Nt9TRjq0NByet/EFgMDYoJOoXbEwu2Ox4PHaHs/wkoaqibACOSxg94K
QcQl+iBWUcokaKxWLCseYlKAx/j6UiLnJzndYjXDJrZSkssAfTFN39HcEOt/XbFr
0BmcDacUfCsop5Jqu/lNyiv4AU6svzcWqIuewUEDuNILid4IlPTR6AYA4bknNFc/
/KX1PimQhtQf0zEwcViZBvIg7pdSk5DPWPM8NGqd9qLXVqrQqb6I7SigzhpumvbS
XtjHPg9P5RFwC/R/ElHArS8EPnLDdDdnSYAiXgKLP/XyCq5SWMNuMFXvc267hv0x
zzPT3FjAUzZYWbBS2uErHNTnsBXHuHs8SRe2TRQvRRlxr+S1YtDnb8Rfl2zih4Ym
liiiXdYndy3JHRY+9qt11KB3ZGNdvnziWu6131ar9hWGKc0L9nBalKO4OW9l3Z3R
+kWlR85nL8McoU+M2ntqI08kdhEW6dhk+Wbe6BQOx6donFjrDLkCpWD4Vox5uwaf
yEvKX5DxYUd1VKv+z+EaAIzNGODL3liBjTGDGbP8hw7P842M49NV+36KvAH57fpB
phoGdCTUofGWgcEiICQoCiu9O/bWLY1AB7FzQro+LHDw8gj1XIPIud1wV1z1kMMh
+eMfAx2YXoJ2CURRT/INuIdMon8F+ZBdX5dtG0kIepxKOe5oXSd7AARt9R0UQO+R
6vywTMVat/pUZLdlOXyww/YKi4hv3PYrQbgf0hgeRKutVIv/LDYCrZHS1Dllg8HX
uUdMcSEf4mUSewuLUeJBuanpW0Mr30AB+TObcLGu93CmJ8mvu+XP7gFoJcEDptXn
5TLEKsbSh/aA8652jz5reLDaOSk80rlbDibKSXvL2CtSLeFvA72BAkI1WW4E9GO3
vM2ENuL1YxeNRa+R5AVbUhwUrcOohGYm7Iwr6qNQJkNof74pSwdIfNT2OSSIL5FK
qShm2j/+MO2jRJqRHDkgbyA9wHEDuS8ird+ChSxFzpptOsHuhIIe2xdiD39gySel
+HsPGTMEs0F0+oCRjxYI8nU9xur0OZ6I96DjB2dM2Bw3Aa7B/G9YPgaTO3fLE4lr
j1/2+1yaTRRkOEK/RnYJXsWmHfJUe+D1MyRdKFEpsjDMlVz/jCUJPNdtqS0t9PWc
+WzBoJYMk3kPPGMAmwPfGJIC5Xzrn174Qed9tBaEA8iLrCyODMGmR1LEljPW5/Vv
TJWJmGQccwZapN9He9hsqGZbCZenCTjgH/RUE/+tAvC6IyaA7ItZhpKDZDEJieW3
YrZXI7jyzcoS2R1toUIlJ2lDW8oLYABYbTBF2poW8xPYs7FobVVkf+VAp0HBokgC
0JKwcJoErsD8hpS0JBLGGFWuxCsHUM9VchUaptNbPh929TJEyCAf2Op4Z7dnEscD
y0XxMkyGTUqTGenmxJgEeuZUr9K2PgUh8trnL/i8s4V0GVj1S65yMCvSpW0JYrfy
Joi4CiOgzRHWJxrnjyG0tUTdVkjB8C7Tff0Ca2cDUS3p9q7ZcdoljkxWs/0pW3a/
s3RnPqJUgns5CUO+deGtpvi+G6WqEKQlL251YnG2Vtt9h48RmSxJKQdXEamfrRgZ
EvYjYvWagI9roL6MgQHvvzPk+jZRJMrdmwX2OtZc7SZHc3fieX/zxaC9hEcTZy6O
yxSxpBKtRUN3uloTe871TSpBjNZKmaPUHgLGjNqaFJwefiEC1BCscKmw82lU/4KO
lr6OGwZt4OiyJxGm0kbjY2JpV0QHv0MLvpLyA6TnM2YJ9VF/ST9lsNhj8iG+72tA
NM1hYWXoTMq9ldnoJAIFKkUqKPNFuO/F2YTQ09bLcwYn0S4fOu+40bahpqRBs/up
DIbiw/MSdmu1kmuO4dPo8yUG9iryrJO1PjPe44jlmvjD5qAHE6W2Qkh/CXObMt81
1ox8fckVGJFNWoY50ZNz6x9OmN0h33ntWs+viIm1E85wSFSAVX++nJTWBN1gOuxr
kWawPHJ5H0XUgBTueMH1pqn8qtgCdsvtXzPO+Un+7+tEC+ES0zNkotjdpWqV71P9
A/bM823XJ8zSKNcQ7HoSzBHk6x7E4VmBtZJ7HJFf9I+zzZB6on3qQc0YEkYI5V3V
jT8WKaUAL1XCI6DJN40kB2uPCJGMwtewfbHGnfs2WoqY9HaOc4wtHC/u0to0o6hb
4k20dxa1zMCqGOi9etbgoZPQbHjJu18yjbHV9dGXdMYT/wDrY28fQ+YgVRQH7WZX
mRbs9Az6+a7rkZ0UlTVes62xSvMIcqwnx/GfSP1NpqnVapfzu5rBzZFvBlHCuIzE
aqJRw9654XoX+5sB6DRXHvJthKNmN98ur4FttHFH3wCogC0o+xD+SPCnC94nlbkp
HATe9F3RyVR74AOBECRbIaMWw0y0v2qXKCLnE7REYwNjCwbokRyd5dYxTwvkIxP4
SJJlHhlaiWMKxrjoDkpBN8yVbBsOBhHawv6gZiYRAUf114ATU47OqKjAwBfyTLNo
9imVD5VFHqp59r9ZTc6Zw+cbMHMU+jE1+prVRXDoseRDZwaiyTr5XGx9MZA5u/xq
4lM5Y/tiVFE0lIaDhRnXY26btOsUuygN1woLTzNl7fzeuvz4JueBMMGeNPSvo4Mu
WIg9ZeEsIIvvVEdP13sfMvOcoMX5H5YktH4xu6dQN1yM9fhJp0YCKSRwmNtY2OOe
lIGhTGgCIswKckpeHBt7RLsnoolECLilcOW0f1YmydBDMk+fGwULUE5aLjOkIVtV
vl+e0d9x1oYuNr1RPkL5i0NUPO7jBKhNTYBPOfYoicJg/kEocelZKhS1EWrkWSu+
nHgB6YVAFyFiak5cZhv82acBubSlC4qry91moCMlrHpFX9UqtF1tQX4Tv943KJUE
756ES8aNjPFW2XjU6looBVCjxOiQhdIZpN4cbjup2bZXNIawAMLm2J3yzfsfzip4
uRbaIKBPU/ePF5JNaZvkKg8JD+0O2lNMGg4nLVaJWeY8OAQiS/zJEhm0BdnzodmI
NLrdu7rRwwOkoGFilSFmLjWgorOz4QCkW+DCjIpMvJgGOEx4+KXV1UW9QNZGnrMv
OGYHAlGhcq2CMWISBBuaZFrTFKYwV1mJdnbipAAamhB5/DVr3HYJMuQxvOCVs47v
UBpELOyeXHHjIvoGOq8+x+pVE9mVCNmWqqiaOn2vlMvjkYo2MpjFskbQN7P68o7M
b19rpser8WJYdiZoEY67lz3n2qnI/wHxMRxk0ssp+SOj8/YCcKmqovKyX+80PwT+
nMXAXWgm1TX+Odf66YK0X8XXPdLmZ7PRUBPMH/Wj2ENyD6SWTVbTWJAOOkZ7UfrX
eee18f3jTDsN8oq2lHuah7d8Yf66GkqTV5KgVsobiaM6vNhWWt8SN2boUe4lCvrP
x0hgJB4I9Qrw8KIQ97K1od+Bl8NwItv+lBej8sHft+rQbGNmZeKR8dAaX9p3W1Yf
oeSowLl6KPYy+CXk3LN62oSLNv+dE10SThvpKApNxem09c4hkh2QL1iiR0E9O0W2
J0foqmkuhn7kwouer/4u0f+3J17ljn/l0j/25/CyKXaJ9CgBpobirvhcxOmjefs1
S1jRZr1zrWWAmUw1mPDicUTQlhFi1DUdQTSMOllAvSAxTFdlRawFss46OJFHC6KH
CBZcXzbzKQ2kjlPHoXJIYeZg7gC0a8V0F+SWDxg+HnMHq1x1bPFb4TjG/f1M/JXS
huKTGMMUJGLpAvDgyvsB1DWsF66x8UazWFrqQ79DVnLyDil+Bf9K2BcLgb4Hc8S9
Y5qSJFlG8EV1ER6tJtoNWki+rrBUCenGIBO7In7ALvW+EaYp4pzmKcdFDFhCuvgt
J6MaDqHwfn+Kiw1ig0Vj4iJN+OxULPObI+L2ryoB29SWB4Sr6vWtSSlcirET7Y+o
5KWqCLMLIxV/s5sl3bHBx6UZSs6rccZ5AQqDq0smZZ6L0bzg7gzcM56v3WIacF6m
vFqhRdwu5aOF70QzwPuI2kl201gMkWjDbwiavuhFh1v4bIb+DLkBbOu5wSL/4Qbr
C0gk6SDayffAhC4tkvSVE6dQvXdx4OEdHtth7fAdQyEUn3SMAnCzq90TUfdGMBJU
xt9WJAxnDtngwOnP7ttAdPAwfDXE5mtO3rDN3BHfyhIcrehatVZA60Dh/EKRY1M3
qkCYp7wEw3IyVMZTY8KnGQrRWrT7GZJVnu35N1RoOlEWd6HpAnqBWXuXw4wHgAzZ
fxGdA+uURO0vPPecFK9KTAe+hhSZwM+kXsOzQVY73XxKJB0e4LafJIBI3IUbVYKQ
soPwte0RBfVXhU8Uo88EgucnN36Yt2/1bQY4atq8pV/0oXVJnpXi/H/+oEs0GU9j
DUjGObfroOkWbyIpqm6o5JeorrW03Hbj/qh5VTpXgtvzPngr5Vc+BIpTlb+CYTrl
noX9ZuGWfqsjXifUMdhp42iffwPG/Mp9ZExLeGG3TymPcHIZvUt6mJy/9o+GZL+2
Rf+KgjGk9xItG9UGiy8H92jwFD5ZnFRkUI3+wzlq30y1dQnPXJ0z3QfcRHN+bSO1
G/g3lsFBto9VwFB4d+QLRpwJNyeZjtEqHRsiDnGZrs7h4ELya+FqJWFB0Z7mLhfQ
0CDVgj1+ruSHECkiq9sgzMWgjvVDtliFMfY2s6ri+G3uPIqiiqKvI7nA79HZlZUK
7vo/NES5MC8KTfawraeFr/PTylTk6C2SzxV3otmHDRHBZqZVXyRPHg8TOf5GCYTl
j4HYMfSrDiiUt+aGDnNMe1AhmFNJOoB8BuaGdrs5Ok59KhT7Nzo05TAEIxkmDU6Q
laHMOGsyb4WTw1G3hZYKixpJKgI6B35aWrb7JHMBSzihZATh9w7ft7gcj2uVGjoq
N5MJY1NZNVYjmvKaRyDYaJB1SDBGECe+jgBShaJQulr6Pfk2/RX20aljV5ruu2XG
1q1DxX7rs/h3lBc+KZab5PdVC/+n7HEYdCMOQl2xbWx3qLtuCcXBVkVWDwlNGVzc
wuT9pRrzMSTkV7e9C14R0LWWKj5vegx/GREO6zcA8qHLerVEbSdJZKEXKTyGHnRU
KTvDn+dOrcW7IY58S+zJJg9xQMI/8agTTOBAu+jEOr5YYo7icrAIl4JtFzUfzRGH
dZMvgftQ29FxuggqUsrXOUzUwCR8dCsotYjxWRd0KNizx09HODLCOYYkp2JTas4W
cNmtarMBKrXhC6uLULBkc/7TvDoREI9kmNK9gpMhJuFZhCvq2dk9FumkWMYiouyh
6KRAvJ+cU0aTxSqvQP8Kc1IEP8AIxDshqmSxs89/cmhMTt0OeiYqhinkkYgYChy4
apIpJsC0SHrcUxhc8AFRYTn+RMeCkCx9BfUO2eHguP8Lnd+UsnWdP2vCMDlgcPKk
6od2z9uOqDMH9Gy/tV72ICHnXjYwXoOp1stAhD6HP2OVHjLJHXVLvx4ibO0KVmGD
6s6gJ/I0EN3L46Uh6dnnbox9xU7b5KI8hIT0DtQsmo0hbsrEcrJfMeWfg88SYcUx
S2U3VrmEBzREqK1GFwzAlMz0QsO9yj7wdahRxXxSv4n8X48PZDQBg3Tr2dm9440J
teY/DlY6slYVyq5aY5p+3K5g/M3oKgYNlYajtnB1ASeyDfgsOMzPsOs3kDQxZ/Hg
t7Q/g+rWibp5OOiTTYePJ2XkfdV9vt02QOsyJhLFLaVjrsbggcl2wvgwQOjPrphg
occxi6Hyn8xLArSZDQu9uqxRnDWlG+vjDFxOtNYPWWeWwsPCvuH2TlPAOe8gNBhG
/B7K2kkQZNhJNpNw9uTRiHZhlXY0DT9l1+AmbijTVjDZTofJIFUwlTdxjZefgwIv
dGfCvezkCjnSTv7TwYV6JpuIe1yRqUDNE3SeE7z1F5G3ykXT9pjKfirzqxke+OaQ
TbIa9ynO1rTJmw3CFPUUOMFLiABIe4KIATs4ijqHWT1h0KJ9mvSEKLo3/vkD2zPD
iyhO9UUYPQdVSn87Sin3QdTDE38/U0522mZ5ibwxdIOtyzAlFOyEmd+Zmn2mrUoU
3K6YHLmKuEPAUZWbFEc37G5bBfDxHVi+/F76hJ8f1969Vx2CwAFMpMdqEM+fj4Zg
ib1lbHizcIN/rdptTLYuyyrvc3V5P30/Qju0OGkE5DqslRYix2qKLcLOBEZy95GS
qM5hrbxd4x5KIdxa+H2l4Ts5d+0VjmkcwRbRxCb4aDiBeYioi785RFuoFbuDuKrb
x+ZlnQOCKfbYBMEhR5QaUY2JINb2EZYtzTv9cKO/jgoqSz0zoxF3hbV5y7NYBOLi
5QTD7bzqRJhLY5raxpZRGHxhr9y4peWCjGEPqLpJoXMYXa70GywMnKoywl5rrbQK
v7k0tF7mR5tfyHraJ2IHmyXslZu/uHi80eGLdw9uZyK7HXPO9X5WriZB32ks244r
WL59oZdA6ImvFzuenLSoRrJ0UnEZQpCCnLCsL3PwcmUM/TjmSIer5ToYwXmbzk4R
xcipql30u4dJQsxgX4mCNqYhHVGG9xcd95QZczui+PNUV7M8+PRmZ00I0O60AX4u
EkdSqfwunCASVjRHI2fOMBv5Iu6T+2dVYYIc3Ft8E5xIsDzrY/1qeEuvkAWC63Pq
ZmqYVbdbsYLjx3zReLkvin+zTiKUbsxwUjK9ma+dc5kmU855wsxQSDJLGJ6WrRh+
2F3KnBd0kOfe9L16VwkHcuATnbAls3aHUlZnXAgmeIurHHgTMsLp0AKNfx3Unye2
hgJFHYVMakLYYOs78yFI7ybD3OIbo/8V+YrlqRHOI0IsZPxW4lDY0EEXzse9l5b/
yIZCLeSR/jJvwLab/6wnn6EFjFmCvcl/FoHTohcXnvP6v0145Af9inO/gmkrBpJJ
cinP99FST5GEN3mFB6KsyD5RpLFOW7YvZSfEgDvTiENxLy7RZjeeIseuDvNqYe7e
8PZWvr4uyTKrKNiLZ/cJqRbyslrpHZvtIJxFDtaBTMF5qUFD1GMt/ItIM7fFycLi
c3XVQ21rRoVX3ewLrKyJv+LIPY1SVn6bXvtgXi3Ps68f0kdyrUPrLAC1S1iR7RiF
OOJOb7B4yh2Y5CLLcrAf8eziv9lHooYVGnEoVYceGqjOaq18A/U7WOZv+WOufr9O
ikW2KdD6807/BJw4TgrRqXGvtABFikyxSV25IF/470BbDtUFNJzfb6lvzeZpKisJ
F89GS9I7To1n2Eq0jqmZuidDYOQ4vG4y6MSdVmQgi8KdTZ/lRZPRWKlcWNgF3MWQ
hfxt09MXcT4qYdEyia+hO22YNk6b6Ky7d3IKq/LfMPbrc1GOBSPTL29mbKFLo0CP
xj9G+B47nRDoEvNoA1lAc9mjWNymlpn3Gm4l+RG6+oNbAYJEKwOdOgg6i87DABgt
RvP4pKYMGn/b1HPGuXTZw9THQaqLmDt6GKPEKR6WBRs1NUHNbBdncpKvGQMd9pmO
M05hGTfMAfL5KSSf+igNljdglHdVA2ocD9Mu/diJ9cQkw3ywc7ShSWoQKnsbOYzG
gIDYUYE3NcrJb/00uqiweLqtqUpFX/4JUAWYPcM/QV6yuDo/HnPJ54rzQxK5UA4m
KuguKFvaSspAYxISgfGhUyWKIu2jM5kdu/wmHisrlfVDUJ3ry2qAO55pnaqw1lXi
kmVieCNAzxokVYSOIqA7K0lpLhuHFs/xgAyd2Um1KriSSv+M9okoxJjDZ6Bi4IXR
MdGhEMVmxieFmh0UggYIXJ695pAEa77bbGz38DCSmo0mJw91fVJsclbc5CcQolRX
afHlVy1fgaP4abtuxRK/I1+6WIXVYscju4EprZ9q4G3yOMXzBkw/a/iOH4VJVGt/
i1nAJ38XrUeBZARUtkQ4xpQ3CX0HgVEL7/cPDvhNl4Ed0J1GdN1u/wkACYr2kupt
g8P7B/5S4syDYXePeg9nztV4eGGhT8CUCcn7nXr6IvytmMCszGu9pVC+HXLTYWCx
QOR7bby1Pq67amO+76UgxhgrPwBn+iSI57cGcRF6LVfVMOat28yYZt9t6DBG3dmr
capkiLTPAu+zDM2o+newQwGO4nxIERdZ2xfzBvg82Fpx8W//Jao2YwDSXVsP92QY
JPCi/tPB9kYr+LfipSFebDolLEXIuhGvRIWb77wz6MZgwh8PhiO3UmF/Y04H4Qa/
OIyTRuHaW6toU54eTaDdQA6gWp94m5YkgUGzzbHmXV4aKeY9d1mpNhr6kPMbGRNr
cTZQWDcinOw8Dkcab1aWKu6eWcwJftaiaWwUDd8oIz5/WNyUpwBDA6BCmSyZYV68
Horw1G0Livuu5fJiAfoIsbTcQG5PZF3gtBiAjTvEsTvaPJ869hKkGwa2PcpbRfdq
jdmyTP/jYUZTP7RkpRsxWKidafyElS2Gob3t6uzZdihSh0slVy7Qn37pC1eKcTn2
j7lvmznRnhhPWnWm9qtYvbWDhP7GGEEglxn5zl8Bs9y6Y1RWrTzaZFr6Bi0mC7WN
n1q9IyVDxzvnKsddLbC3Lbc1ice2mvxuw72pa4hKmsJg5BDU7N0JXx+cnbagj5Iy
MrPG5q97NYl4fm/y+xS0eA7MODNXTq3Rrc5zod6tcPGqKDJpNHPlslJeGoulUOox
f7Ft3jSQlDMTcPZGvFVb3SI3iLXUJJwO8VOhg13UUTIamOajqTaeCaTUOrgUEPFd
0ISxIkdKHmhLGlOj9Db/PENgj0aLkqHG98pD8UqaeauovcA7vlRfJpVe+hzo4KZs
GzJLB58DOW0F7RWIeEP9mctVVP0/n4QonBxsI4/wgFP7QMIVM2kXA2ViEzhtRKkC
IjUq9zvgYE3fsTn+NgV3/WARdj+1RIx1V0h1wJd+7emPVhSzfaEf6UMGbRvRevli
jESw1APJwjDB/qP2yhZtyPSEOjrhxD1aWlXcMOx48x5jzCGuuKDvCwn3qSuLs1ZL
d/S9Uo0UPm3HdFloQeTUTacA3O/fvenwYnclXiNOgpfVTYcCH4QBmLcOO6o2zvWy
kGXglY99UWA6vYxT7L9X1D7jGZewHYkZvf7L5EMc/x55briPlhPn35PVpkFeMucw
a6j67JAAm+4TwWVnT2Mt8FlUT12ZAYwEkjUWR1mSehzfErzlUXXKSaxtvT6pnN5h
GqPm1ceY7cjZdTuLUODeqsjajpH8w5T5jTeuRw+kFX6th3gBy6dm2AJKW8F2vVJ9
D5R2w9VdYL5Ybs7T5dY/5MYIHsOBJ+gUL1CB8diHSvvjHRiCLkJB9D21Nty8HPzq
X0ez7Ff0+g6dxvsE4KtDEhVnxUPIQ+pdh5DVRG+Y5WongrL0LKzex3JVFh+PguOa
79z7lRAphbrPXTO/xFgUrINHX1/gF7wdt1/xPYNw2fX8j73Vy5V20YBHMlXkeh18
tiFQN5cxi0pDriBGU2F6an9sX4lDusXCYY20pPFHlVK5Qv3h/YbVqbOi7J5vC82X
JkPNkoi0ywZDO0Dx+qqW4VM7SOW1CgsyKKLsrntwWDn4jiPV6lcEDkPve4OLDbiR
5vf1KH5TtVKBNOE9OiW7Yg4Gmy1cXyqO8DTrHK0KbsqDzkn5x632LaUCceDy0yDC
IGsEiqgnrcp8D1VFRUFiacjYKbd0l0vR0nc8I+Nzqp9FU0Ppqj94plLxkevgHs+D
oyaxXKxfQMwwblwTyd3T6wphJhZUuG9FuVHl/9bP+Nlist2tBIvTk4duTqJbyxcM
VEk3Xm3HXX4UZEqEGVJHJqIoFeCeqS8lTTaKncgMz5VRYF+WhT4doL9aRfx01q3b
rFXdnK4QimCWcxGrQ/addZqhO7OeNlrqIY9wdnQsYStOVzxVdP0SQDePkfD5u0rv
Xbsg6299GnBPK4SQWd84c2t8WqX4pqoUCYQ2iNpjyhXtLyG9n/CaQf2Re6OXq7WJ
pw1XqprEV6d9jnHwUkegeayik9/vXcOF9gtjTOvmXusOpeQy1mibaAsCJXYbklRP
L/IU4oLHGASVTsQG7i59+pyNUs9YqvVQJTMd9VRtAECUkQ34t5Wk/C7xeghPK883
V0FM/DmW4fHTxqkT2Qwzi0aAW2E+DJ16+HG4tB10nRF0VHdHdj/w0kjC8BmQNDLy
zmH6VJU7s+ru0Y6UwF4QrJmJepLqdl+gaaiNVxjbEQBxILC9cxlwkC8PULjifw/c
RtJLS30lXpencpzVs3J9hoJeHkX3/ZD09bQOKIDYplaM4+iKzVim+6ooyDPYLBFr
RpPeFCeoFN/FZBpgR3MNTGtmsEaJwYSKkAZnJgGYP9Zv/7xKCQWIysN3+ZFCwzX9
s38tXs3Rwld6d8lgC0Nu4WJWijX9gxXke5VyKrZE4KxAhh+9O6BkekCUgXev/hhg
h/7TV2ddZ53PHeaOppvHwkl/3MRD1mp6qwLOFuJ5+CcCAxRz280P11bclps5u40O
Xiqu9dLyN5wP0Ik8CQfsvFTNAMufzReZqtLgBfcQ+5juBpLLrVUXUMdSXX8AQxaJ
ml/bYOicbHjRFCa+sG6SyYNpcQVG3ybTKY7n/zOAbflZzcM0QleAWMFjSC0XkQci
e/Y+1ais+FNkH+QN58MDDWB5L7t2EdSk3aClFAHqUzHxaOTzlRmEUzk7MEpUd5NH
YRh15hrUxipeMxCiEedhRj7PCwHFCq08t9ilgHFeX1PEQ/KpSPrOZWENImnfE8Va
pENEqSy8zVnGq8UGVyy1emz28BND7C7KjIlg4u8t2ATos8xUeatBhEP8BdSI37KR
ebrwR4jY3C2GB8rTji/3l92GZxgCr1jQOuKxt2BgFtvoUzCHWqI5xW+h+i7AQIWw
0yxmmD5C7rWUIG3aq45rsseqb6iiMzsETzMNMj7gcywoZLrEurzZe48nQmojrVC5
wSuhEhEyWmSeBayhTI36P0gjl3nZZaQ5Ko1xpgS86FOgOwiLISa11jnavhspR8k5
W3ZMEQqtrn1phiwf1iCQGdo5zsRQJGrPTbGvgp1sgGkDJO/yLlXwlyS6ibD5IcVJ
3+Pf4oPM8Oxn5ULhsFxk63OzwqLrANx2CC/zOeHQGmEKIM9u1jmd7ITCLq8dZnQb
cyxIYhuTxRHnxIGCeSrz0gSfVqJx37v775tan8jidArIQ3dtPfqkq81IlI5nxOT/
5K2YpnrChYDZ26lIKAxwYFLj5W1Eicf2rbCdcZxyNy8YSkSirRFsqAS3MjOifVxe
by5n5z7ID7URI6XSS2XxWJKuHWSEF2v8RIsDXoqQr1i8hDDnjixQOh285iXjnDO0
MsSeY9yKBXIpylFg7MS2QhU170/7Pgigy1tCqQsQvVG17sZw1OWlw6dw4K6o1PIP
Do32sXiQ7uBkbakVpalmqpmfZHYWHMfeeihpo3C61s7kWHfi5+NTb3YpOn+05IL9
8okTNJYhN80j1PEegYuhMdh20KWhbRNMIEm2/X9NVKzqdp2rzVSdblcekiLzmGGh
/7xetref9CFqlhqn+6y74+PiROrCWOHrr0zRsh+t693j6gDPopahohpZUoX06eIR
JWIdvJD9mQkouP43E9UxOVkYqkeif9DidyUAzF/UeZVuKKkI5ZopCT82cuDbc1Nk
euOmuqInt60oM5mbzpJtF86ugHisQz859+YnC5DweLB4jGT7Qa/3OpT8szaveIwV
kOfjE+xLMZb4r4Kebi0qoqOD721XujgI+azAvwUW1cTGRpMNuwuKLoEnf8e1Dnaw
A1bzlNoD5oQlaKUCUadb+A9FDj4rnj3Unvo58kRa8jFa+gul8TCeAd5Fi26luAoj
1iqr9J2mPM8BED+XwDgXBT+6KEVkJ1BJTf6uSJrpJiiOqS6EDtXd1FXRQ4qwBJXJ
6dFgWuLnBd1xyxbBh6JBZb4EqED8UDO3H/sf1a7OyP4YZgEXATXhdWjbXUHhmwwp
ciRQxoOmGUpk118Yk8PJQ007zolz1HZv7Gh7M401FFynq1j1BXC/rkKMrKbomXRy
YLZcArdxG79nlfWhOIyX1khU8DBRal7GufR5ajixyYsnJBJBXO+O0lmqhkJ2OGHq
UbcF/x5OeHxw7kQTjPqVHgVwGCrZx6iULC/+KD2oW8un6pmHhCy0WKKOgCIt/gng
yXx+j0hWr8r/aifm+os07110jPN/TPaacZxsmAktBJX4HXX+6R3qQaahJI4eZIIT
cHtq/5x71xpWuQBGOgbwwnb0QjPmRZGE785hVReX/SD5U+Q4d4FjrBUZrBzWIBvG
eCWQaEfscoth0a/Agdp+rLDX+WgDxMkTqtJpH6Q/BA4dY9Dkr64T6cDu/Ots5yU0
4rMsi8iXQN7W08a9L4Qj+rivu5+fI8wKNdJbI+6lMD7CtzxIUUm0lcbsqrCBmGfe
XCgaWAouUhnc9NCpE7qtRdx0US1qRJLBIOdEewrG8yYRs/wzoMGEaGScu0jL+eiU
QTmG2bn4xenKgp26w+35il83rFVM+BaafqoAPjPGWeBfTVeqe+MS9L7mwdplxM8z
/L/3tzEc/6445SIaJBF7NA98wLwE88L2D45Ji7Q8vZyB/w5JVh9rqxgCzEq1WlmD
WTMHNP/0G5ojyA2qPmsy6P+MA0cxnefYjioZGXVvzt1+NCBBBpQdSvpT4Bmar0XT
yfo4JXgHK60hKwlH4ygBqx13y6pUNzg92u69pJYsy/4kGhZUNeO556Q4Z0WmGwlT
9BtcARAEDl/ExRDbiurFBipqzX8E9D1uFohd/4kwAmDwZuBvV/2wJo/fZo3k5p+r
9QtztL8yCfwqlOv7UUumCVw8cg/dxGgK5AszMptFZtQMxPBbI+kKf4UfPph53vgZ
/erhrnURfwHvI8eXFuXSbxyQO8/wDVT3vwQsz2zE7A35W+EyFrhvu8P1ho1UlXY2
xIrv+BxYyrimozo1fPe8cTA8hg3QU4/hkxLSCIXZI968h5kHnK/u52Ea9IxoZ/VR
WhonsHTpXyQ8uoJcGWdEx0cbOThHw1YuXlgXZd/TEkEtHjgspux3bF73FbuF0gmk
FIIomACuzdd/yZeKVAiTrjnc9ftxQce/JeBE2qnn45UHAJv2atX6e2tuSbr89GnV
y13qDyPNQ4n4GIEy6k8zE9pNvLeof21xTE3r4W9slFCC214smQQv7g5obI0+0Pzx
iB4cSQaJS7raBLiqWvHZtCUBAJ86h4ZstOYJ5yDuB4jrxxmxmAOXWzOOg7HR6Zi1
umgHHAXToj39xflf1VnK/+YDbZhXzI7jgaigije3Ul/IWbbku6ANqWHASvnZOhox
9PffqXIF4JDkpHCxdTijiERvZAEKQlk+pQ6YMP7NRB2wMz51Xk9OzccmEaMRWkKp
+32g/2Yd+YQIkTDfkv2vY2zTsPCWzSd6/fDlzRjld7LI+fCJa62SLM8gOTtlOQPh
qsw3O7mDXHPGh5KjguoLkLaMvBZZEf6Vg1usNoSZ6+NE/JQhsSrghtMkRo6T3Uon
xMvvs3vvSS1imEc3I2Vh7Ajzr4NyJM6AtqH+8liBoXoJpaWfrRGVn1tpVl2MduTw
6hSFxZivINKWU/3VL2sS7vEX8uPsqcnJ1iUsZkQbkfK1Y1ytbbxBh1UUt3iFg9/J
L4mCjle+C1dHUYfUp+IVNiuAyZ5/UAQfi3SqOECQtqmGzoQNWX9YVG338XaeWfVm
oUEdJ8cY6VIP8FX9yCAMh/rCQ71HzN8dJkDSO/5a2l1BTNZaL7z5UpAevSPWIOjt
GvR2cLJPnZ7sYScFajA35yMPBImDL2WtrRTnsLyEclOmljkil/FwbYToJn68roCH
SgUIBzvEaHbwbmRXvuwHhjr0AnIXOnhaNG+YI6JXQcEGbhyPeAJJrkRCn/Y3JvFh
Ta5skb0L3gPHHEcAfgKB9N9gwyBl8xssRTeHaLVp54CNMBss5Ae4NadLOOo3rT58
48svuabVgG4FikteIdWdS9JF3XyCAaSWa9cAwK5VAQAbpNh3qdxdFNnJ7a0wnP4n
oG+wGtodVrW+q8NOeYSeJaABeoyyvtgL+sswpr5SK2GtAyPfHcBFIhMBYJDCa6oL
SQuAEaNgB4w4ngHboyCSsZf/z0G/UFXP44HJ+OjDz3gU3Of5cILlpTr9mkBOxAEV
INeIwhGWTKmdB76dn8rp5hzfVJpfvsvnzMCE20MH/WNseh5QQBqMOsig6QbbnmJ3
U11p20BhxZXWWq1GfFBYjPNPVv447ipJUdv2ViUjLOZg+ckT6NtxXRmDDrPcZPX6
uSbWYSw7CMswD/0tF6u/5U62Ujrr3tlJ9vWVcaRNkuIBLroyQSteYy3OD3L0pkkQ
JwejveGKcNq3mw1pEyBBnmXu6gIqXAQ2qqCALtyuNra9r8K2xgUf0MHEDvAVFJ8c
TcPz5XJwu3t4TyxiRy7ZqNcXpwUhnGLYafloV1RHCbNHe8A4gREj8O23U3YDlzkQ
1Vz1VSty0o8Ht5AmLog/15mj9vQkBYx/lYFtXqGvU4Az4e+LukQ3ujsK/NBAyk2U
GpM2gV79wGjj0s2Nkh3o5qTP3a1PB9Y3tYpN18CGULIq1b7ihRzdMbVBQdKypWVd
Ho4gkl8xMC7KsC5NEUPPH+19LcEK6yivyfo8Rvs/89uLdpnMjp3Laqp10qglNawW
qn/Mxm/6F7wegsWt/jt/dTHi9gyExD8/IfRB428p+BfThR0DIo73AlnYpj8xUmV3
IVsnpDtzPV11CHOHcpAB0tpq9sv4xfIxpw0Dl2PX6jjo+YXiSYe4e+Hg2KGeb4xj
4x7TaraFZ1/Z3SbbdlHHhVHqg8o11yxVvL9QASCEzwc0bIBZDGmja1LfjCgQJJQc
v5j0D6rtvfdIg2cAh5GLiCcEoDlHJUoOSnAxrftvcGk/WzeK6v+o4ZjHKwy77Qmp
HXfWU5t0pXKIAOFq3ZnogGsNbdehp11FxcJ3J69IxIc9E9UlQJGvZ71KbpRD+4U5
dOKKzSF+JPkWIfS59sZDRHXeZ5QiFmnV/i4cePNgg3DNFvQ6B4f7AYIcrurqy2a7
0rSDvgIGrI/18yQgZ3u6LbY9IDuT1dKF3amVeXsnLHsHF1ldK/OmYXTDUGoqmG42
0o7Mvs/hVs3GBHPyaOjD5jIEvMHm8Y1jMycjbeWMhbrpPNevJpkpcjDuKOHH2drC
868s7kCYexr1lJOxovXuwbk5X2zhvWulxQxi3NAtewqhjP239iDRej3BJxwlY8+4
jjoOUim+m/QGn1wtGph5fUGxm1vD73tnLEQQl0YCH/ig2d+gs76LN3IAy0VJtE0K
M7vHWBWsTrUYohIBKfDtD6uENxQE2GPJjKdx1ylLi9/X+oidkpQJBokeE8tH7cN0
nICVI5J1SffVOYTKi1+Ie/ZiFel/DCVrLoJS+fZiUKoa7ACwNbQjz0DTC6WYggmX
BGN2Iw812by2yckCn7v85B5iWTk5vIshQmyohbRjQjGV+Vkx3XYXhvUUC9Z/ZjTh
DD8rc4mNZo5sqCT+xIDj35gKnPFrKLdof1tCxfPU+BiyXJkQcf0+VdWTyTApI2IF
zQqzou8XULoaF60r7faYGZ4bTAYbxH+5N9knaqi2Zy2ySmUDXQ92DPxLQ6WicMiv
OeE70/Ixz/glkgAfdtLGDE6tioV4ycrDAeZ1OMRnjRf3ZaCxImfFLbApGXuGN4I8
F1yVrHhgK83+EEEJaGvlRa/hpPfo6kPGsEvha74VlDViNx2nQK5OKLo9+hqomDp2
PR5TSZtgoiixRlFWpSJR1iw6H4IKcOiLWl6Wa2OMyxQGPD9D0b9LldnN2wSKo3wg
yDAv9kdjJS1qkyg2ha+u1XWbFgxzag8tRr1Wfr95MEJu4CRCwtsWm4IeI+zFs1jj
riOWLfvICXv1j10DC00GnXzuBiBvg1pZMev49zJ2KBv0AYnzUFUTo0zjtYDDErBG
cF9sUjx4sMXuatdXYOzz2iNXJNB2/dMFUirEL3mbBYeRB7nV+s21u1Qj7ix9JbGY
vMDEaaempXMz0VHUecsW6CgXclSe4R//jNwKInrx5glF5cPuOqpIohaAR/6KyeH2
axARbz7wbJ0i04iq5zRNTalj5HdCBMgRmRb6f9sPCq62niN8q1yK2QsrVMkroYJn
CDPVV6bkHcFNu5MuHDt9K2tlDxocdK7JSkBqN0SF3Mmtar1lUX2PiJ4XIHHQUpvd
i4hVzmzdQBowbnxhG/cyRLx0WkatGKamQZaBhjS1NqoriooZCyit9mLJV1EtPdGm
bfUuWGh5stgOsEBZi18CR86hOXMxl+eAxBLXUD/pNeO/xZYD8dvPgi/ha/fU37D+
iLWihic5w9xL1B5a7tZPW1tPsCcthTUslP0Vm1aLkSNA/ZbkKTU4mGI+SN/ACk1/
+4MHsDLEA09fqithb1GUM+2/DELve0H6cNpyN/BRSG4x3H1ywh5dm5ehwu6dqsCx
p/rQ4B9Ox2+ypqUomFmT5FZcffOm73PhfGqRX6LV2Nk2SMYoAVvy8GWq0t4RnrF0
AMXRh/vS17EYaLh8gjDNKARa6bvtE6Ou70udWux2ZRBJeGYxcWCalPRt/YRU4GF6
B/67mA8R449Sy+BBJ9lyX1SsWvtiBtA80p7obf39Lrc02lDnn+wDmBSm4RyUFZB5
WG8naTtsyip4eB4WT3vy7YFBvWML9dgGAs81u3qlbz4Un3YDW4GuHYEwK0ZRrXdQ
MDxAkPkkr8IkEGB8qH4DRsTxplKOiseDB+zhqw5nTqAnlAsMQoiLERwPNUtTkOoD
rSORdozoi0X3BxrAEYr5nfn9TFtg3dSDZOrHmaKl203QaP4kmFuDs9fm5iAxVnYY
lFS8vIUJxzEgcqWELTuar9IsJA2v77Ekb4d0UInf9Oh/XFXLenD7YKthGV5rR4px
+CoP5ToX7pDjTAxarbFomtt6QiYFmChJqsRDwwWRqInThbHROcHHRr5RmZ9keW14
Ma+FqxR1bEKfJECvBAIv54X5vQn1kavJeourjl8RQUU72Ia0jroBvdVMsYDXb0qT
KKFPuD7yyWgjdVtPAQ50Hrek9A0eOpiC28cXZ2k8TI00p1P4FpfBtk0QaA8EXnUs
6D1aob+nLrecEewVAFNsZbuQ/tG3oOP+Mh7KnBe20p0u87eboewoGEMqM1SbkyJ/
24eV4ZVXnk1D2AwVIHxJxIdrgE5R7/leqopqbN4DxYf+L+1sVCDB8dP9RQSt7NhF
o/o9Pqmz/vUDLBwv760fESDEtvXATnFSYvBgXK/NxDIyJd8R/dyDhEsETy/XzWei
tEo1/2AFfzY7TXa5+VWocuV7l4ooIvHLg7pEqNDM/cyAfc5Skq1A+sGGp1Jsk51/
Cu2U9LEglnVnL1ST7VfWj3BtujpxooJhX9Vz5Oam8/SQ/gQJofuCxL9Rg0wFw3HG
XiWlbYz3Tn+hyhQtyf3tno5LoZBktS1IcUEnrZHr44KGtk/QJ7FOrNMyLt6r1Fr1
72l/LDjF/jgOneYIYZCyNuxyfK83aLDrp8p9L7xlHdcVl1i4yvw1FlT8tRf+RtSM
LIRNNsOfddpHvfcRyXpBUunPeCPMQBdqGiJ5eWX5MEb26RncjPs9vfKoyhHs2/BP
AN5bHYpV84AfQbDyX8oA8lvi8EyFpCIarSlc/DyUraNDPjN4q1YkjS2QDdmNF/Eh
7Q9jyG29U4M22fYRZLPklfiKHcVqp9TnjXtzyT/2IDSw8vlgfcJsdWjEUoODrCRB
Ame25ZzGQLGyRUfwT5ouQstrw9pY9eCPObQnXdeHcdTzrQLF0CB2daayyrvHF7Ei
7zJrFN1QYqihwvKEBi2XQ2X5S2qBaCkQmry0mEIzPJLg3AaHFntZtkz3tyWV/Fcw
AjyMKlvlXKA/Kvk8seLts1DArojXT+Yvqmn4yHhoWr0uRivONfqjPRnySod/CFV8
SftgOR4n9NRp+7r1j6wWKVZbV1Grb2oWli8GH1fmRDA9HeyUysWQs7e7ulAE+HXj
xmeOBc/nIRG+FgCK0p2a5c/pZP3wJavOrtqz8o7R55jXxHFHC8YGFiVPriGa5/dg
qvaJuXSDk2vicFcu/YWh01tFdKI4c8J5QL8xUfgkK+L26OkzcxDIT9rv9bV77p06
W2DNyHzyBw9nfByZ4ILDRYgXC2Kutuu1sx2KOjy9R5F9XRMhONPi2lNwJsRP6aZT
rGKAoOt2eE8PwaJpUY3itU/lVb1W3+wBCV2t18VgxYM2wvQaydeFIKj3bDI3S76G
KirVeKsUj59Bbooqp02J7tofIrsH5Ha9KR7n5MdWJQEXJC8uB/4O1cGhZSVTFeCZ
tQSGf9TOEFn7JXzCmnnoLSOqBB4mECedhCExmauXY2PRtqSpPB2r1mNGz0H3CQnt
V9yIGaJufH8+v9UpLfbTRqgcLLW1pdL21aK9UmpjF0CQgy5vAnkHWKZO4+ZTTVjG
+am1pyssTT0Swd7/dto0Amqv092hcn1UsxWj/zunYE5510OlR205iG6YXlZdc/UK
AS+esEyANh0nbGUkvHccyZunsoFn92sIMnu+sciYxZrWPx0ZXh07z3v2DPn1J2PU
1x7Am+SGW8FnmXvIjR8AShwPdf5rfxfRnTwo2+8XM5tjZCDkHCV12gvxHzRnsuSR
orZHIiFjIYe/RxGrw9qKu1CXR/ceUlsFB4PPsL0KPSzF/aJlSDkuDeGpzolBJ53i
xkyLptt8mGYup1DC82JToAtfMv7b0cLlHmt/tYmrOeObobcADSS3F9JMZCoMLoB5
Dxf4wdqIqaacMo534qOpcfgdguCWDhLPg1pfcWB260nh9k0Vb3A40Vi8rk0amQRI
iOg84LO0yq+ZXO8p2FrbdNaIOK6ufrslKqNeU0ew3K15SZZC75Y9VgAce6ARLpxj
caaUuGWJh7MmFsG5KKfuRPcSPm+otyCwyoaTkb7RaxQjeSkhcbOZprX3gRQ5sbJN
8IE5CUE1E3ELWv21G7eQ+ZJ2X7gBcd1yIGu9vRbjc5eLQXFmDZoS0xsUBJnWXPPw
jUU2O1a4S+i6JKBrFApqviMQIYZP864VsJpkQBw9CAlso8/UmcCHgEa8AtKuQwlC
R23mY1/75qudjjX2riqHvtlMVJz0t4cboqRZVbU0lOMcbNOmlGmccwQjdjAIz9gH
78qnpcaUYowQzQL0bmFx2yejxd7YTgfAotHjJR7vFzovK6pRli4YfzUrnN8wWd4y
cQPVA00+HfDBFVnWBtDLOWrxT54Fzm7wzwShJ0HPeeYM4ZyVAGNF8GknGZ3Pu4nB
0SjDBsEUVyL+IvRcGdORjRAEBGmsk2+1yMWIlxhVDuaneBfonBpOOlXz7puiAXWN
RwysMqu1OryE/XYj+XY81XNd9Nd4Zg9Yl9E6ocABcOm2/H2adUIrNmFOE9ELoQ3K
3qyU1i8Krqtf/ziCgfNxc4X7cP8jgPYQcX+j+DPXlUmZj9d7ySZjThOrE7cuGZQN
yOhaANF4qOCxi8jqHF24A1wrFeOreBtoazW0eDXlNzUNC8mnLqO2oj9+LAT5O9R2
tQD5sTXxEIFyLXPpzzlZuIOm+Be+1c7pIouI0RtVOfnYv1a4ALST1bEEKpyyTLjb
VWagQ8JakPuceGMJx/IB9jlTg5f5eWKh2i+vl4jQsCkfq+qUYUmMHHgjbqwX1NO5
3lXwoC6J3QudqP3IWfy4vyEgxiztAcjcOuHjKI8EEv2MB4tz4uRpD1GOfgBGzi3S
AsMxpKte3vg3S5wAoL4LIIFHtZ5cmAuUoUGg6Vjf6b/6AKKiSR3RrSkn5f1Om1Cg
BMIxiVlxibho7+9TU+mE9imQyCMyvhCQU0AU2Fl8XT5NzRjtT/lGpuL4ekapCONJ
Qe/m1XtkLvmle9UMTyAkDkbGH9v3afBx/OYcbNeproNHkaAS/X6N4hjHcH5EMrY4
RdfgjpPWrM2Dbye1wwrCI4oA/tLle4h3mE+blU9hZlxhT7ttxGeYxP7dVYL9dAli
fwyIRe5IPQXbEwsSgOXLvZfQCKbY74mnrMUiXnDof3VXC/dwECalb120dtp/idDP
dJSJSfRCp2XbJxBdsQihLxIi3YbKA4MFzsvsXP8niyvlQjp6oy+3RjaNBirRlKhs
0Nd449jZOsEM+lTOgdqk/seJW7wN4adwKCrVVFABB7Fl65VInExu6sjp7vRFXmpR
96vtAMzIV9Cz7A7iiRleURrwhkp82UXABOTDMuygO/UBWxhnPHwRF9Oz2zUab+hI
An6dYZagrjCeMVBQBqn2cxxwNOBiJ6HnYIQBkUiWW6hwNOPwsuaXSiBV3J19Zc4o
vapQJAiRI88MGqL95FchylmGRHR5+HDlCBAwS+yO89EiyOjWg/BdNGbfuxK9l1sY
A+5tKLac42UB7JRuhfIgNTFCn5tAA3aXoIIdrEgCPY/rHMlSFsGqr/negXCVR+1U
WMwHGHvDV7MSrZfvz6IgRzPq9SWtTRvZ2ywHTNrk7yrFgKKBXvpBFc2GDK9E9wGd
0XgAGFKoGQN74TwOeGPiNRISynY0BxpR2X685Q6b8l6pOQ9lb+kMERhQwyBp+3h9
ZNuCpBvvsON0E58UaKVyBpi6v8IfnuIbup0AvxS215FXrbrzQN0a5mOVk4mWIDd7
JvA3sQqy5Igw5Zg4rp3PbqsHBUYrzmIMfSo1Bb81mdoICjl//z6JuE6wc1/W3o4h
34bsbLWMIGB7U+KymKi8Ai+kK7j2rsnDqnikdRNguTI51yfFiNzlVKMMvMkluK8B
M3+VKTwFcSk345XIQtglKgTJWHuT9Nv+0qIFW0fjwwCr1XlOaMvCjctaTsJZNAOW
3zrDqRYfxttL2NTJ97ft1IYhqs6NCSobHS1IjrA+da5TUoF3ejJ/gP6hgn2CtvUf
MH9hgOXFdTaEMKwlu3TJDAzpxr8PbN9sK/EpgnGmt0LQ7CToZuZvOUMrFbexJtat
zcFUdZ/+WJ9QPbW8xh2vB899m/yuNZKAR9EZ5B29vQtMET0h9muKiEkPuxxH+n3R
v70VUjP3rgMga86AJjFAmppC6+pX1EAzxH8ANn4XrIyLbCcllSTLQx05FvDL+zFj
X4+UdCFQnD3rp220oxH1E9Hf/txbPfbEFKFFvSBv84hSDWjZTe0QUALLlXpKP5HN
He/fNVmrrRJVNAIjh8JComHl0yL0T5JwpEEozmudECL/FgQ8J+2GaNsiB+7qfDi7
ststzTqMhaw243bsiNx0mlukFjgSDVv1gVNSoLaTtTfaMQiDbzY/KKr+6Xwedmur
dV9ez+3ML1fyIAVN9CG7gt0kR/v3uHG7r0YW94Q7zHEvWEj/bY0rryCHkp3Il4dy
53+f8sgCeoA4idsXL23JFQNVC9eHrRE3jmZM+6tOpYhk/SsrIs5HWErRvFsRi6jx
/p6Vo4epOjo/+9fSpKIaRY8V9uhl+DyoMW4j8JzWrafZ6zJTDY8i3+1ZdUH7v356
F5xeoeMcfXrkn3qoEjep0KFoQ0NhmOq4JdLrn0YfQ+vSv+ycV32QpXpw9Xf5uA6k
8EtuJk+uzhF3BNxrW4SkDEOHKhGNN9cltKpt39XdUBRFg1CBIQ8sqCIDQXaNOpYh
1e/Yxcg6UoAHgsRZmN4jnJFzUKJNlgvTArBjcqR9Kisc0QEhf+oWFQQzkxTkkWG/
Id7Wn+7CSvFM7YTfiYOyoxuyldlqTvTCZRFCoqivmhpTCe+2k1MGGr8J3U23Vc6U
wRih3lLYj07I6w04+7tanoIybw//r0L634O/AIhJHrMqTPew54bRZad3Bc6Rb9/Z
HIFaaoXv2lIGVCpd/yZXmNxFCtsnWiYSg3J+Y/0VmtbbtrCf+309iTnauXfpqZP9
PUi/UfCvIF7xnoqglNHjzpj7L/PVJCkOUm6jYJS8uVVdbu/oAK6nN8aXe+6uaifN
xTZQFq0HcHd6QYTeMmBEFAJ0fEF4zT1uRRc51YofgDsgGE7QhdM30Yxhgs1e+KVt
mDO1QBOsc3BLlL8RiUbIdP8YMHAdO3JPJzMlHmrZkD4BHHhtk1Tex4gM9x8Vawq+
+amw14+P+13/u7Z2cGNXp1yVEREoFJPsh08X0LBVKc1l5k3dp+gUOokJVbCTo2y+
p2jSm35jm9qdRsCkBaCPFRGZlXK6n5vz5e20yMlnvJl4kJTGj+Oqb2eGKmkZVoDc
O54LPXzLncXf1b0syR8NN5k1xEYGjuTxSCSknkm9XTZbl8MI4kYaEpfslzdLs13u
5KkmtNxqKKhHEwfuj/MzMK0G6AHL+AFw/9Q41kOzmZbF47DuUce27EfQQUIJZHHO
MKDRDEuZ1KfR0vOOoHb3U2SeNXYkfv/zKasoLVuWzDGFVU7NR8VJ8HLuFeir8N3c
WYT0Jb/fgRl8Dy+82rMruA2uj1/fo+cXTqwIoaYM1lprCGU7ZPDe2A2ki4+AvoFH
udNQTs1r1LOlbX1q8A5teY+Nid8gdsvuNywvPZZkG0g0gU5ZUUEcyaZnHAVy/lHu
0mpBJDHrKU77Luqaxd1g4XnZxc84UPgaIcBpxFS+jAzvL5lDn2rXMwWiK/IKaCX2
eRKreWoaj1v4D2SP0jrXIzkUO8y2N9MP9C5JjaCKrou9A07rPk7Z7o3n8pRaYs/6
1lDyWovd16szUPwEIOcXnQ4qT3wFtgBdkUTRTKOKkbJ6GuH5Glnw2CqLGx+irh8/
M4B9+8bU/6UdyzdZQJs2fB696N8aK2TZdMwn+20tUfrHBIO7k4Ry8MJeNb1+s32j
iu0i281JUfUAWbX38NraoJZDaL21lGERTtv5ofscbSEP4MBsWV7F1qhCmeg1eo8R
CsoY9u1bAk3toZwsIgHe/l1lpFpexMi48rgKTerw84eG/SxGIgYZYwMh8ecuEBfF
vSI0hXQ+QSMB3qLOO1D4oIBo+b8tbwI72hg4/lM447adqYIMmdUy7uExZMSfWe2e
Coh3W/q6m0Kl+MlhRClyN5ML2PvtGnSuSmTFXFXYeO9IhzxFsaTPOtMLR+Ufd/El
Q2In/gTEzyWB4aRhJCAcYcCW+Luk0bXUwsKEvPig5jzyWMqhonJb29uvwNmTP1vp
LLWtL5wc5pYsnTtmVyLbVBd4F2/orG1eCuSBijoIDgGitjEXeHhY/TJFIB9w7xYG
lHZjxhAckmOZz69X4m8m4oBBZTXvNjFiJDwYJrWHMkotaIozPDy/ayMs1SPm9TjK
0JpQhzJHHswJ6ciIMgWFv5Z7N/zky3Qh/UxTT4W28CqGZEbb5kIH2d6qCwPXzoa+
D73iReZtHNKfeLsLqyklsspIsfm1Xz2sqh7N6FZOarqb1WNsv/tDIVK5ZMmd/SSu
ZwZneoCagtjLNxOAf3fqk0e4c36Q6DWoUEUWNO9ixopAIYnVXyJNlN88VAw1hHur
bTkmkvIlW/0+ensh/k+od/aH7/ZTg1bRfDpMBvgHYPTidh92OX0KC4KfQyQ7CR03
r5ZNAL+n6+7394kYJDxDP7P/6tjaBlcYYl0bzA3x44/hIXvYpBiBm0v9ZN/ZF87l
jtGaJQl5loYmOogpXlu3CXDYcklTDjScR3A5bcCeBuchM3POuCdIJby74YNQCPwI
y+XCh1fSzkNLwHK+hVygU+v4g+64c/bzESsHjZoRQvTSNJZdtPtIs2lxe/du0smg
js+0xnRDzdA3UtDTHI0AVF5Z9AyeneU0eqmvrw3W10EZUO3J9YEja7KpFnoFqIjh
3eqTp3eqBBpXpQvfDAg1p2oGz5FqWGPgdglA+MlyWuF+zfWhpmct8jAC+iHDY7qg
L8UpPcLB0lPGPOvyc9bzaj08d3hVPHD1wKmLvY7C481g8iGIS+xiaVP3Jo5aw2iK
gKUrxxeshIbEzLIkEnbLIOYqWHJBwAu0GA29A0f5SlUI6bhLtnZbQxtpwgwTB5XD
bWdf1GTRqMN31vewP+/BZne9NNuCrgha2go/Cyt+mMEbK3os7nvYynsQB6oTIBiX
Kr6FDL4K4PRvW9zFnjWnpDIzMprWIJBiqKPKWaPUuelZjiKa+WwqkWP+KcECL/0T
QT34SPUr5VfcY1OpZRHgwrzmjiX1uuClK0TagRN2fT7Zlcp01SwF2F8QhgtDoiSP
DdF0OkLkxAnf4YUpVklAl68bEYreS1hkj+EJ3ql/anR32/ySgZZHas79VJHRvfx0
AK37D3u+bIzM9A5+sivihqlZkXs/VgiYVx71/DP8a7zbt9AC+gaP9/4n3W401rE4
RmuieZewsrnXC03ra323AJL0sc//mwrIqVJhSu/qM7M3voW5g/LxLGtZI6cFynoT
GkhCadCiOtVgpQWhwmOruhT+VWbBQVlOFQZIxfVBygUBHsJktvPKiRSI1lvPoNFi
ByN6uIAPmy5B8tl7IvQV13TiXWelmcTk/+SDBSU47LaVxCdEp0hHjSE3hruUspDY
dqTW8Em+9JO3dwnV5Hkw9cUUXC+ug8uz/SjlbeuN134A3PNN+MqZXw0oAM2a+/Tr
9W4gy/eUwrbxaqAtYZmmMMp1oOBsNEhVFeAW4vOL1JHVgxXXpjJc863ylS/aMp2n
scSgJUJ/SXfCsICzszWb6FK/fLNf5kWVm1qdFJ4a+iHTdNPBWmOLziOj7h6p2UVw
eHYvvCF7gS8vDaUwEvjxQouJ0VgUajYruNSBD+GMEBh3ccFZor8MhQbLvlg+ZRaH
fL6EvzgRGNcHlIQtm/b6HiaLhHpGyPnMBhPwKi2IwYqi9q5ziGcToxQD+0IInNpz
jnoWg0q+EFZQFRQngaTbSub70gtQYf+61j8vvyu3h8QUv/U+QVBK77SlyuItkDBI
YJ6P6Q1S/K9v8AIq4z/91G6TOnD33SMyp+YOWQqXPmtpY852jS5MHSl8ELongT+l
9afYkDQeQDezEZ2EoOAOUoH8GSxdMS7zq1xdaD/CFbVqM2r7SXCI00Xaxiop4sTA
5E3Dc8TQYQnzgISufcIDjPPAa9uLU3wjhF+4HvyF9Nl6V6XkvRhhsvR+InYzdfi0
z9Z5AZCGgAcwuiayXDOyd+fZMFV1PyXW4wh6+OQ/c1//gJpPZMVxUfIHiYgzaMNv
oqHgjcPeKBHNtmkm5/M7RFGz4/oSM8KxO5ZlCDJsIqgi398yy0oI6eRwOy67SYOe
vMbNwb+920JGV/LO1PlV8knAQ7nnVpybt2j5LZYU9zh0rmF08CykSQNa5UU5bFIC
WDfQrDWAOqEWf8q02Z5oarzL9z+/PuPFSvQnCI1G7jHRY9sggYpy1X3xTzHc0V9/
O9uAJylmJEqboWPlCftvhD1yxqMWicDtO/GvqDXUw7d1xJ5Z+TCBxQ+AetT9A05W
gv9EDw99++ce+3cZIXzRdBLdB04w+WO+odprs7LOnAQEcwnJTdcagP4n86lmS2Ml
loM21dcccqz7QAv3Aukelxc23WdUHUw67qboxl+BmHtDE+zNAmwwyo5yrPhHJkZP
S4wqFo4AjKcLxry4e4a6tpzKXICKr7rnOn/2bCi7gFoPLfpShFoZCC86C8I3wC9F
ZRLMlA1dJSHFZ4cJytru9/YeE8W9VNZbbcVHP8H6AJeCWQFBly7HI+1+vV4iKFvZ
ryIpbBFxWlWj0X+wuvTubdpp0wp3ZDV3QlH7BTtXo+GGrczLNW19qSALjZaLHCuL
qzi+i6v0OJKlrku+zSEq6mGoiWu9H5Y9wegXrd67oR7jTIm8yuUGETIEN/RFPzQ6
e/E794nIHZGQWhisJk/ILa4bhtmPR1UNSyCEXJ9uiWFdlzrwt+vfALFlsXuDrS5t
GJNVKuB1GaYgg6sw2PejVGBO6Vi3WsQtrDVHhN9koKVh+BIPUEA3oshDuaL+XRaE
qR7YGAoTbLu1dyCB12RXvMtJKGUrjDWXih0aCH68kNHDdOe2lw5qNHHc7E8j3Rv9
EwJqCpBTyNLRtHv/7vJzrsZtUIY6c2KlDwaKkJJBK6Yhw/AlFT79ahLLCUQbajr8
udJh+eoU/BDCCGbmHFpwy+atOBxrVTLb36z0AXgYabevxyzI0cum33zvn8sKYD4r
mWAniA8osKWf2dEhTnincSJ89B6UAcjQgLJP5U9YakKf6N25Wqs9ONV3mIJqMnLV
0gZM1EK/oa0vJuJKDRVwZho5q7L0TuBC65Me4tPQKsQ0Z33V2ReqycQdzFA7q8xN
gBO2pG3nq59MsC3iaJWTIQtKc58I5MWkT9Gm4JTnTnjPWftPdPFbE4VJjZY3hJ7H
DjEbvEQ9BTfp2M7WQozzCckxMZvOM/YK5SspYytPxWPR5J5mQsrwChMSd77Bstny
V8XX2785+Rw8l1eE8Tuf4TMr0hIwGLIsN444Sh23kSqyOYWoI/MX9Q+ud0fwUqRa
zG5mRFohYuzkDHPDdee1x22VFrpGkBJ6eMQBrL6y5skyAmmKxnAjN4ZfMck5niet
nIgYLLY6geH0DJV/9VstOhRw0BkJb8ZcvswAo8UT8pXoFf7jPrApNV3lrp8AvgKT
IfvwM2fUPKXJ+aCuNxcOJpomn6PJqsrXWufejXwCsK89ncMiarNAzjmfW1c19Kmo
O+fvDqvLd41gGNjZHQjeYLryg0UAHXKS4iHsfTzjSKY7Wi0xMqSqMv+dLSeiGLSh
otNtlpY/s8xsgOq2Ef731g8lbjiINn1aTMJbuYJWgqA4VgfEbo0pjZ4Qcd4Pz+yz
Rag4322KaL9lUczdZP/X6A61SpAaCUrcGT4qyBgkCmVnOktbKOIR76OlOnUXVpBW
HKOpmiLyu+Uxn3K75F2ghoMgE6WKMJXtGf3Qu121Fk/PGoebp2T7Fdj6xMO7Xj0p
DsdGAGdDr0Z1aQhCP2ex0wNld6P0QD8pCyacNW43s/qQWfu0GjCuEddke7sOJaMN
AR7PwBKOUp1PjlgjEPeN1ugxZ9CfnEajgKNuyiiPlQhBwEUNqHbZ3l7yd7ZLcQEL
hL2k+ka08UCJmOFKMHYt0Gi0gTNlN5dZPOztAdoG1d7g8aUcgSU8yrSNCYQsuAqG
k+f5XuOTpsgawsF58D7Bl5VNVIf7wcVUNs4rK+T2YUBo9ev6S1lCGfLwBSPbHU6F
04bunmfIZa1M9oElwlWoChYUdPVouI83xjNfSqoebrzH3Cn/FIy7LuZOguGb/hVr
LSWN5EuJw0vrhI2ClpP1Lmrn2kl67P8MQ754YinB/0mQ9am6KFbYcngkC01EjE7e
dD+CPZzPRM/u2y93U9nYdouiMINhepbCzk7T7l45UQd2jGcV9K30rgTPUBIpd0+5
LQl9D2xZnQM9c+pgfvdXRIf3SLvs35yxZeXoGzqvaIqyNgiSn0vQvrfBa99/5Kp0
82LOKAAJJzzV8UzXduGSWVw99Zuhy+VcxO1Ic2Njp03ZjDADO/ifmZ9me2gnXrrz
dwB9umWhCC7q/9F0dSsShdKbMv5tYTCkOd+IwqkF4lbrZsHWpJuTx9Nt/enxVamV
1GcxBAu5i/quLfcDyYrGAYdGgRb6kvWcl02Ik2+bRGbo1V8ZfpcnIRhFXwhgT9Wd
2qpUtqpjW67fxyqT0/KhwQTSfR8KDid6DH5hELND0M0sRvfLBWqhKiuGC7GOekjh
S5PgW1I4G1YTOiQzueFffy/174+eHcKpyLuPKoZPBaL9dF7mlLogaULVOxJsspOi
HiHrSHRq3PP5Sho1Oj5FNhUl2VmGkE6sGzC1jqdnoPO9g2ULvBRJycujH/4n1Aum
IUvJ1nTgjyhLVOKV1Z5oCV/aaF84OrrK9RUfkU5rAdTatpnpgXdAMZ13SAU1tU3y
Kccq2WTLDOgSAgve7wkCg3lNyAK1BXMSLVXLYfqSE8DtY2eLDeIO5pXmWC2JoEsy
YoX0DRD6D9yvyFJKzBRKV6GU622TGosUHP4NAMJ5OsUdprVHcYI+ck1DqdkyCn/j
WGFJiWvOxkRsXtS5DBV1IYVlAa+dKy9vqHt3Ho69cT6Zhhu60kQpI0/ewCXgBvh9
FvcI62uwD2qq+fQSgbNw5cwlTOOcjpHQ9NY/l1tAlRu9Tn34wHNlhvW75luiP8j5
Id3YklXuguFkjdCqvTfacUzF2PkIHImbJVIdVIVsrniUzRUXdoHZu9ocTSM7PPkT
xQWQUS2Q4nC6SpkWq8n0mUN3lUFY3RNe4mwUnKzo9aX2dhIQ1TLLRI5xJ2FHp4cW
NnLXnZQeBURdzOyfYj8T+f9KmvHnuvNSL4NpX0rdCTEXDh+XyowHgJ75D76HsKRg
cRCYjpse/GRiYSCQ1S83EwOSxiSpmBynGMpSrbB1KCd9CWsX+TuMHmJjH8zQzmrs
NSADNzL4WaO4y1ojHggZS5NuoR/zHGw2EFrQ+g7LlRMBeqGp152G+PwEiKIcIYvu
p9bgcekvb70HyRUOEa/rc/mTRrZbGvqfjBXekQb8/6YWyPd6WF9ZE3EJM/UDl85t
0euTeEQigkhLvXeYX81/rBvsh2JRjDKxClK43BAQrq6tZzyvn/HmXFxc0asxz1Un
yDLkDfWlc+jRqf+yvoDJk6cnDe6wH8s8nBohTgYQDyoBjl40QdWHmVclaiOkECqv
9JxMNlA9vJGtA1qkvDSHrsfK83rT4s/wOIohhFVkBN2AlN8z9QCKyazHwmKOJ+sz
IvHB1HvLIi2+AkVmscXiQMl4l8Ef0Np3Nr+H8M2XGfZLIowTv05kVy3AIXrTj4zH
HKShChCEuZ1ZUZshiflZs3AMih+X4nNfO8GX8A/bVGEs1mlohrpScwnC5jtOoTAA
2rEHz+kb9UxvooIm/6ztPNhMI3QusaViGeOzBU4dX6YTdXMPDH4WsFSAfYQiVosX
KAkWxWOnakxX8APCXLcanZVUPTB2518frqQbhcTJXtx8ZK0I1s8NmZWC4LYtlPRR
UwHUFzBw6apKTDBIiOA8HNjAKZ+e9o4g30oeLPNi5qI5ykU8nXffbXZO0W2NAom/
gwWlhsxC5L6CPFyGg84y3ILTWclyIyiXV4MtykBcpscHjqUil+1IOrDE3UQ8N+r1
7yHHnBpd8bRk3RF1Uf/oDw59qPMw8ikWqRMhgnF3FwQMVhNsxf0CKr3LeqjkmefH
dR2MCJ5kQdWYHhlXKNSM3crGbHOnYwiOnvSAVD8LAd8wnvfw8cT+UrJegsaMLWs7
5Yt4xVGQb2F1NLfM3Uehou8LVtxC75pf4ICPFDklN8n/j2dttFEeCv/A1osvfP84
w0ekS0f19j0rE8RleTJMSfHV16AEHFN0cN1QhitM/Yl17hfhc+hGQ7piXtnPuSlU
GNiNYS1maeiorJSn6PvubaNT+sv3Wj+yG8bEM69yv8ZXGc6XdR0LcSwQ+AU66thC
/p/WOrIr+jKLRrfVzwA6ew87zZz36NoH9WkR98Uwrmb8X+qdnm+6LsQ0Pz/A8W1/
XzNMnCzvdiM8EJxxZE+xRtil2OXjR4jD//J5wWE6N0rKLf0W6pRPIVV+qEBmUGWp
ddlDeKh06Z0bOUC66GlL4Vr0QUi/VEMxWHpsTKpNe8UAZzqjErynLJXqZlqFhq5R
2Wd3XXdtYj/l7B1MDBVM3YGIHlt5WLSRKB1kMr5zaMkKzSj+rSIg5evimz+dNVFk
yB2zvmUqxmBsaJDshIAXpLh9p/0uwNQ/Ld1DG/CVRGbDOG+zdyr+n/lIr+tuLpk/
pWFW+zR33iHa8a8+X/jke55bk9JPSZNrAjFuPsCz6ZGbQb8aSsbWCJe86vutxbK4
hiUy3FTw00yTkTlcWMJLC3VQR7hHQgQvRB0ww0DPCQ+jONzIFxym4X/pEoVn8V2r
gLuyTDaZsbP9ASMcyB5TxgbRp+iNYs0tN5H+FRR/9Ug4zWspBT+xR9FILrOa/i10
pEHgnRUhnS0XeQhPauSv2p3j3YgETkyh26RfOho1SCe2waJ41Xg/Sr12SPK0ZxPR
9y76No74JCfBGembSR0GL/u+6gz6tlbT8CfkKRyv8Pf1FPmC9FVeSr9val1tWhnf
O6DaI9NU8LClcFyNyLRqBnqt4RyUMyDCaOHspUokcN06XWEceEt8C7w0LL+OYWW1
ydmMhIW86n5c/LLM2IqCFPfQV6MIvIIZ4HtSuSKyr+NyTcLt4ix/9hRkq4avEyWW
uaRCl2a/Fd61EvwBPSNBKW/tUAGQ/NP+/1x9EeVde2ZLfvhxQTorNoFbcL58FS+e
r9MLxwsaWZ7zJMJppefAtle5IEGRNmIL03fygRjWV6pfCfWrV5s4UMG4F8nQDltr
54/yF5KxNKCiMok9ru8u7qzLfhF4wHd6cNpvpD9wqkstaiDHmHYN5FQKH1ZXiuOu
hfrWiTqAtwf+/T+md5sY9M4ELImKiayPgiC0m3upSgPla0SoT4oHV0Su9veNYN1K
++V0QkTIzJEFo4MLmUEezmaj1ooJi10ioOOnNG2bg9QQv+N38S6t1zG6eFwH2JY3
eKGTP2MLSYen4mhmeQfZgHLddlHv77tpcMSpzAN8LakujkwmMYZ6geX2zdtkwiSl
hKZpqRTNZaElMdFCM6sXPIqunri6mH3PnZGXtC00HtVn5yHbP1jZqtzgE/wP3HXg
aD6eWLZLjYNveVW6kosGLHFca5LChYtX2SjlzKvHtFe71iIBZMONXGn1IB/wWRqO
0O6dkVXxfBVTDQIzpuOGId39ah8m8CP6lPmkTpWsW902VrTvTWcgJCwnpid+SkKB
stvvAPWEbpr+GhIF3nm6xEjnxDU940Mv35bH5jCLJaQ96mcKkpYGZJ8mkiNpltGU
bSBey0VYSMlkiQcLlo2f8qFdGVYBAh/ak3E7uagjpv2jeICCEj1C7fmfYimHB/34
6kDpxEW8oPCNG3ZbQlpoTWyF90To3ecGhmj2wF6YDPTYqyO1VtY+QSScRD/0/rKo
wssiOTrMBE9HJinDRaOmhsbqYlHSQl6M1WLrNmIYVBlNRXP21OPl5HEztf+J7Iu4
3Z1lX7C3k02hSXIz5IbUA1bkSrHrAFTEbKEgFzyWfEG6F0/LAfoa8wSb8cFoOEqX
GMZGleATuNlarFraslSSQA+usMATC9h3sUNmUx38wAMevwQePSqRNpn8jm5B+Xzl
yEOdD4jNUL/iI5QkOUOd7t1DOxxr3qmRtsX8yhWxClfhHQCpjpdB1HCfzNBepprh
q/TDevZHeuHtwVxv9mgKqRUdzFzFSQO94vuWZW/eykXDDPcF+cn5EuFk5xmSFf91
qLW51DHcgySnmTguDZs79rVHxlUnLPNVmqqTJfuRRMIIj4GMwrEWs8aRZr1tdhpH
cBkMiaH8w8bDJHTmxDRXyB3mwMLwZEOffRlbsloij/XX1dp3KtPDvBB5aPI5pNE8
Svb8djjKuLdjMGz7dMKHZQBE/a+CxaNERr8jlba6WcI1wl26Ph69ciC4061vnK2d
ROFOjVw2e0y+nqLF/HF3dLGhvNVsheGeBHiaKQQvVDJoPuTeJ6uf6Mjjaz5lS6KG
OrGYZaT5hVE8E8iy3ZDG7gGp7eK/Z5Zd/8j5JfflcOrcis0C48Uqbp2fuDsq1EK7
rnUrLCtpKz4Tht2h4sAFNnmxGAWF6Dcnr2MJ71OXs8J4LRWFUkhK8+qmT0SHc7Ed
AbjTnsLhiAc+oHpIidi/9d4Zv5H1zXdzgOciNKZz5V4Vg1kH3GROuu56CaBqf3Q9
xBLgG4MWnAWjPy9W5lgs0BNKANl/vIpYlAZSiK7QhcVlQMx0JlNDk00HHvSlg7+d
18RM/2KeCRKyGiWyZZUrg4R+sqil57y3aHAEw+00mx2pBaaLlChYazBmT/Xs7G8/
mKrE+UAedOtm3zfw5hOeWIwXr3g65FloPDDn0n9wa2EU9ziR9+zLyg5RVVdCAcaR
EcSZjSSfHEAI4MN2MA3u9vSSS48r46WdcSEnCDHKCW3bxJ6ruWS628FI0n5TaLr8
TTg9u08of0BnNe/EWHPDdMPVlGI+KFs9TwmBgT6ntvzJzyNIieMsrC/gx8+JXOim
gbPbsUltVHTNBjAKEEbw50FZEmDhm9+FbIy2Sy5ZjSX6zMP10xA4ZUkAl/SGxqBP
rm+en/W2IJHT807I5muU+KQH+XRLqXMytlPKZAXn0+r2yYF61gD1/OzVIrSXF1WM
05sLlxIYd2l44ObmMs4n17IVCk/8eptvHzpc1mTGiRBRNrP5xqxHQzkfgLiOILYW
CkkGlQYOzuWU7d+IU4xMx+W2t+hC9wWheN18gqiupBe2JhRzCx69bKt1YRFVh5oZ
v0el5nWqkVCUEIT/fCYqnauDCTmfZDrFlmkX9KHbPdEVGcwAeR1LVqPpW/cN5CE7
z8AoiWW3yVUsnXmbbjRfm4tEYqohFvqpMPP1MiuXxEpkSwMDzn91/rOcMSeB3XmW
YqKYbHKIsGXTY4EmWlO+l4WvbLsLNvgmXEkT4FL2GJ7DMKXjzZlicbRh+1LTwefo
BFG/AJd7eGgHWAATkDEmC81Xs1j46XPr8e9wpEe8bTviZIQMY4SflK14F+0RIl1G
6Ne15qs2ldOXJQchiI66oks9AgvlRZHgFDv07M3hpkTpphlxhHRITBAF9qdojGkP
7PKTuMSN+jQj76xCA9mr+gEfm/cJozi3++B3eur9tx+Xu+VBTTyixZn9huXU1tcq
Gf4NobT1bp1hMiAp9RIOBIHeKy+UU8dfVFBAPNDtI30FBg3DS8MH2WcLtztqlR3o
4mr9SWUDitw4ggMANHqL/B3Ej4y3IBsLybfTdH0bMxi/A5gRJUE+P8wVJ7liN/er
53mU6nkT1NqOvN2l0tdg9UjLbuJOrZ+SrosnHpowvv0SHxndtpkVB2gGDaxdxBR8
UjTU4hk2uUHAH8ZHPZKY+LmVFNEEkLuZIbEOw0/yywZkRhIGqFf68h+EDoW2UPBP
20I0n+ocrG68t9kgkJmRgFFan5wyfcMGKDcl6/xT9KSz301Ey9v3QGVrct2N9evg
AB/urwvgOZ1+/+Hz9FMaY85yrHlrpG85xgBQl8hkHf3/+FCkxTpc8jgKzJMop+dT
IwPgslLOx0Vi8MyxxZtXUB+mf8XSZTywu/5QBwNs+0uQBBh/rNareKS9B6FxbkEQ
dFxkSC/ZdkPqAqavfs2tu84fcwe6C8/SgcZxJOKdnALRGpkOqARHh+AKfQBKhdhk
erJ7LqktWY68mNKylHsZyVReviriaeTAawWkr9Oxrjx9zMpm3KWQmoUOGpfbSahq
+BxT57AnvPKRGrdUndNY4waj2Yv0QAxWsXpWT5/lHpE+jLDfWQzFxSbhe+e8iBmc
+8D+GpjUD4J4PXYFmMW6KGCk6gb1VNq/jDVP//1wsrnc/X6sdVKyghlVP8ecxcmG
iv1n9wBP+T0XMO6xgn0LPqPZyx4lkmS2H5fcwW+igIQbqjKnjndPCFZMNg4DIWw/
AV8S5S9b7lb1Glu+2qDU+jpkSXw1RR1WU33efLzQYYWXsWl8rkSzyo+H8wX4EbiB
sAoPIOrtP4GTwzOv4oOoknT8nuRDP3a6g5Aj3vnskKeWM9/sPVNILjwYHcT8U+V+
IPRoxdhW+0E0RPFpdJnB6VhA5NRPBL4M54X0HR+xCdEeFrnF3QNAzEliC+Ny1TXV
m/KDCzYXYAXKIVsGYTnc3IHGjdTby6Qw87RWKcwMkVFHcmNSjI2lX1h8Dk4nF7R/
DNN/QqUKaRJvvvt+1gHrijdx3VmizuDP95eGwMF7NxdHnf+MP6QRCAnX+YAs3I++
54Yu14MlGEZEqXWmAthRWRcwHKF0PEv7ABFccam5kJR99RsUMc6GqTzIbfVnQb/V
gctnwJzoyYsGsw++xCAvcA73ptnYFOuNRRLF8u9YpfKjDOrNYYX/HeyQaNPStzRv
ikFnMiK7gnT4ugmTXaer7aq/tq3zN0FIDFE0UqokYOeyS2RaiS/pT7MxiPJEFL48
gcgSSJZREr5ss+1e21t+mbdwNRXBtc3PK1bLBmWqtVSMnyBomHCRXuFVyOJoFKbZ
Y2aPJGke4GBBT+uVRtYCreFkZTc+SH1mcmFYxyiidp1iKdDqd64QEs2WStXInhAd
SWwXlIoUsIlUexwobUBCjGajplZ8AKRDLg+6V7A4/pGEWXGr0eB2DPKRoEWTfNn0
Z9hhepXiuphQsqgfmEp0NLz7cNJ4O7E3zPJuD45I3BQH5VowNBg387zxpuBhQ5tm
2mDuZYvJTtk9UeydUZ54GamzZfFK9jgSwmkvrsJAv7nzdhDuQP1o/5gmqtungQ+l
3P6JMj75y3v94Xq6y7iAodOItwXrY/cT+u1qejy2bFMTPzmRGR19XA0R+O1L4sgx
5AqB+HlMf+SqWwpCOpZpiuMjvqCtgFzGlIhmo0bMywDUmDK+VFFZwD7iZBHp2vE2
CWSljK7f6aOxQRSi4eN6QC0mwnuyfatJypA5eXSAtoI9zTUBaYIaqE3n4lsS9uXt
9G7eqsCRXsIJO7vdGQTr8gT0MtoGjE1FKBi8orCzyH9vCyyJaAuZX7UFUzSBEbUz
SMCQJYA83BAn4N4MklRnH6T4GGZSPqM5mRjAlw6Ify0ipoLSjisXumhlK/B0mtrV
DJwU9EXgGmM11mOnnMKFAeXbcpgdj2l7VTGRALq9+DsMb0uhQweUF/Sx/Tw2Eq3Z
+lPdLHdx0VDYK5HacwKBJuznFqRxkFxO2TQlPYtlQ/6YU7kvhP/LfHhZHFCN4nVI
Ga3h5Jp+MimAMX8OhryWsjaObwcrmVs0fg5XbShc+H+yEfWzrJG1qQ/0TkhiZhrK
dYN9TB8SvrO0xo+rUTHoODp+NIYiSkUXB9H/VGXNQMo84CyFhvnkg0Z+eBJddPHY
sa9I4ZQDxbxfC2wfgvpOeEvuEp240N18L2oZ3j6g9ObYneBoFNoVDIvQWRvPjsj0
aaZXF+Z39kQDEnxy8bb3+vaLiCCDXGp48irt8w787uSDJXV0gLfrIIcSvm0DIWyT
3xNqikO8jumGgG4lkcEQd55iK/sIdX3utNcdO5uV5QGoNTW9xtxtjDDhf1iGvZzd
i1iN8go6cat7FBvoNeSMfAMUExNAB7FM9J2klf+2iovOW0vBU14SBpAeDlkjt/4O
7WO3iJ3yWJy1g1C9oUeo43EPQ+7PWHM2Q8xYg5Rq9PxLlTDugoTiV7WXrmYzVfTB
xh3BTeIv3kvAaKsqdEXjBXYTJMuA8H4z4GsN/D4C3SUL3LDn34KIzGE1w2Y+Nteo
Ulv75SPA+UKkMjswqSU+haKFvReyJueBQc2QdwONTbi6YllHrigpLXC9gAFOFFu3
N+fRV2sdJxbuyRCiCVn+pdg8FRmywRii3T9R6qrUWNCNzTXuor9SiojavVfgp/q4
4IFEsqhhB1tQx8Uav8Je/CXuk/0vmmkMS1lUIEEFUh1GXK4kQLNXhHhqtyjl7KJh
uOQ6b0xmJrVI9ApX7joAPiTkBoc0mmFk0fXahAp0zwUovi7uvXAVKcsJpiFj9MZW
Tk5W0yD7DtLuFf/ov4752IFNFzdTKuMkQ4HU04IIt4rXfV/wMRWNNlXZWXAmogo9
yHfNj4OpdI+XhF54j0mquXQVN0WvhasVDDssuEV4IRPFcRe0iQMIh9ioAtKO3PBQ
P0QbOdQaFDqgab3RiYlU3ldTCBiB8KhId+ISfbtMXt0Gob4WbcTG2GJKoY7g9CXF
5tsaRsVF4HW+139KmaZq2dacMFQNHpf31Uo04tXhlqXU4kuDuMRd9zHuYkicF0y/
/ooRbN/eUgRuhHtcd2g0ohMubwJciCJngfovL5KAhgoRNb+8J4O57TGoWG7Px670
/SAsivHaZYdj7/DfvmgoCj7wTXTs4eD9OcwBWLYW8r55RA0+m3TgRNMImTvz0KpF
HvUmSYLYSh8V4NKcDQ8Lms3AAfRMcJUR/9ENkFJW9QjvBKgB372ufF7SY1GbLFDT
2QM8s/64TdHWjCUwqiUs3JI2H+QQPbJjZ5NSN1SAnV+DYnNlOSw+eXlR97EokykQ
pHHoRxk40YzMzTGhjepBqq+RgrX/b7EDqytQ4dw6A6MGsb4xKFAUgvho4Bz/+0Hn
INZjUadrKAWOgrjxbjW8VHJCWddT65Bqn/b6TpU6lqgd8KTBv3coESFbKuy/dIIf
HfNByo4M06nCtmH+YBd6tA9wPLL162d9qD+wXL7pnxrIR74eKsS0AroC47dHPvqq
ma+y7sHc6Oqr7aXbwu+Yig2KAusAmOlpw6iSUzqn1y+QWUQ7+1nK7e6lIX7J8sqM
FZ4E3LxXw2BCdt5wtpCEnz9THC79FU1hmboL//wq2YMQABm9v16Ew5fJvtN8/etk
FQJoIrTeBTj5P5dZQKy9KjYTwKkl7089oMdw/g1Uud9R00VfQP4LzHqyAVTxz2BZ
1vlwBkYnLQkKeIpWqsZNkfugJJ2JJq7qrPgeAARjsQvyF5teEGEbAPTEAQozGQ+w
vfeiZwKnX8Rvl79rETII3ndPnr8v2StpF/B7YzE3uhWvxejEXPojHlGdp6Rurnz9
NboBb6KMFu0CONEVTWRifbHWdSbruSDlWsGNhBbh3n8dRNQCQyiiY8DWwwXCdAsb
ECiJCT3LoSt3pwmfiU9EtjsWBJMKfqPhP1TSbI+ejDplIz/XP7+sXBeLiFNsmR6J
jILQu1m2Q7iequYgxMn6X3ILAhRDdCzOiOLpHtiWzliao2kMkVaoq+7nEggdihYw
pTAMA80xh3TpnkupBa+yUrIkBbihrgk4HI0bumS59emmf4wG4ei0x/PSv4DaWbRJ
08ea6o1X3lgw/wvFV/57LSN+MggDDMYIdowQT4nPo4JYSUKgLE9ZakZYvBIBdCuZ
mfyZ895XBWlxQVZTs3pNlvmdAdZUqoCun153S48ShqYpxBxtV5q1NFhttuIwefsV
YK9pRunuDvMlpjsKcXvpTohTQp2iIGInvkbKWmNMK5Dy0EHt6EpqjKBkZ4tuGRDA
hI7EdFnc3UkegZdUb+TINcx//S6NQH9tZD3VFk04lSoOfWjoPgSl0F2qbZT1OWg9
uGlZ/l1YV2Y0pz4MFcG2ZZY3dAqExgq0uAbTaaFKbwmTBk/9FuWOJDxp7Qq9DKfu
3XT7h9/JaN1wMmhDn8pOLw8oOAz092nc79G72C8MSN5SOwEyLeyb6mPQs56sXL77
F0LQdGRqcj7BceunznOi5Rxmd4RjuOnvTLmibIwm7EgoCI6lJIZg4dvYvmQdadgx
dirPx0etygxGOlfUPS4WSVDnH/31O+5Cgci6TaeQJmVaMLzf+4DbbFKyxBx+Go8A
M8c56t6w43d8bD1Yr73+EXfVh99I+Xdzihf+3OHvbShzdzM0seh8u0si8v0vmB9V
Pist3VnNHlTTuo02rtEXq5Z3f1LWarFvkBMrzRhPieN/e52aq/BcmxW17WbmYzsZ
caiMhmGUGFPqBVJNnGACmcK0dDbzc90wdIAbscMGZ3+mDY+4VWOQ+DU2q8tjCn89
rE1ladC4ryMnqeYHb+NM7hzvrKYZNTQICk3/ZUHWZVkLtf0HEoUgkK2M1LrcAq7p
fiV1PC0pcQpr59H4hFcuUvBCq+66WuWJv+c9Ke3ZBdE66XY8zW30awQ1tBAf8J8U
pRj4hqAAJnVpzDao1dEUK2l/aitPZSLJjjM9nHSfnt4ysKJRi/E9Lol/bs7Elvab
SMHRYJNYja4m9v1F68tf6gdDAHXf5fhuvGOnw8+F2Ld9VGQw3IElQlSA+RUlezDd
ufcA+a6maI6ZjdBHe8eCn+4Skxag9LECQKEywXBNad1RXHMtZL5SkQAHeqLxXyBN
2yBCg3EkmFnJlrhOh1YjQRGB8t0MiOKi1U88d2tjpSoykmrdK9AolX4EI3KzwyHJ
A8U7lbvJRoBpuuQI/t9yfVSVIA7jWaGWjEo4e/72RsshHaG40lEBGkXYjgTW7c+b
/xlTCWe88igPw/Fp8Y6xpzZO0c9+/K+9yjvlZHu1LCIqBTvXAKe9+1Pjq/74QQph
Weqx09kc1XnGfrK8mCiK2ANyTbNEy66Psu3oO2S1cPk4rA89KReODkAijYCMmlPa
SW1SzBtSyYTjuf9q3VUHAmppiwYbksRUVlNL4QebVj+qrAOavrdonkxoKAov5LPO
3Tr5IJF+TxcJK0fe0qfVQp2KFozewz4niJJksfaJFDdjDmaHqAinO1UCVnNfomjw
pXJVL9ReVyvR06vzrXzFCCdSDWFmW3ZUaoCiZqeVXZLVHIHALzIb6XIefoqwN3vo
idG6xfxVUZly9Du2TGj7SgQKpiolB+852ELnb5Wp2zmlVc347YkfRvvEcKYbBMtH
G8I37Zs+v1aw3spBICth0l8Pw+kKG02ZIT/RZpch8zUqnOQAmrJYAzBeb0rGRpWU
5agJOBmdmWuc92I+NNbQSMobzIraXVf+rm0/QxPGuG8cB+q0cqQkTM6RG0GASmAc
4rBTz1pv7Lb9wI2U6zA4hL7HMZg1ISt/5Enq5BzkQXl1DdKryV4VSPcQkTuyFNMd
tRsTQZs8sAVV6rOT/RtM41EUqzCDtzaNL7Cux82zO6WBn90bTIa1ct+lIBDFiCpy
H8dQ/2afUtbZQND94I/SL3Nksr1nIy9HP6XBdHggjAECx5q1/gBkrdyp7NZU6aML
jgD65oQSzA6Uu2OpWuBJdOpmttP2LwLLdlfPSzP+5c5q0wNGRlqUZVjQYCtOXxzx
1JiBTvOROAXIUT+Dfs0xcVuWPvrIJzhU9os7CltCI+8QmpZGR2SHa5e0VY+JQzPY
e4+ngbt6cgrKTIAikW0he6zJ5IDzyW89+uVSN4AN/dTJVi5Rnb7P/lNrW3uK3sGL
SLP1nFsBzRL5W4BaOoDEFHXxbjAoGlrqmLtZ56pAFtkLaIS7rUgEMvTHMoBSY/zb
SLlbUz2jusOzXWFhkvc0Hc8fDpzle9fzs4KvRIahLjP+P5yBzrh8YqecuK7U1zAM
AxJ/eioItNM4/8Cq95hQ6mHzFaWVXuAYOFGtxPKICSpgAJ2VO79gA/maSSyms9Iw
JUGF62Ho3LeyVuRO5tSLt2ED3bOJHi9khBbKwtNFxnZOGK7nAfTHXmQXS9WEGl88
FnzCp8X7bGovnUDszWVIi7Ld+u/w8pLGxVSe8ybvlZ1WkNjXCeygKAfJ4baI5pAK
+Zlk4cikTwDEbnMP8km6pmC2kmtjxyM4n3Fg7ugwuu1B6jaVyS36iICG19aZO+rj
ipOOYDbtsqwDGcTuyLsqpO3bfmQ9vULCIy5e6hr/mNaSogaUbLKrC2uXuOk4lS4X
AZfqwAQ4uje98fDi7De7vhPGWtWcUzETAFGxBXAeJZTtzQzWwOQrc932IXDxbWnY
bcYHUtK50exqmTc6c3N7W6uxrJS7ZS6hD7fxcEUKDR3pKZRcu8IqMXhugIvlu+/e
F9nL1R563VtyigZ/vHpjdufrAw0v/QW4dUFX9QTG/GE9i8wiUPymGG6oa+DBDcv/
IwBonRQRBlyQZMmZz8fS26W7nk57Y0hrCaPj4lXTvK+1BvjW+GJNuUnBzB19SJf0
n9S8x/NdXJZ53kS6KL1daC8dpOYe5nPykAdsWziO0lW+bJoE+qDDTgXs4WX5PX5j
9+szL0lS9ZoZor8VDlL+t4Yst0eYWkKtkkyaDXhycUTvVfYvvjZB67t3fr4oDJNY
ArQkTCml0se+r3lkuxNAEMqjbj0iFolLfUI1Oc9tyn9wJKM6G0EgBvDE/lFt/ih2
iDMEoRpq3Lid8QLgeYS+Bo71U1fhfW2nHlKrbVOecVWT1i/CXxbrgEZ213TSj8A2
MgvEKbyP5yKroaCvChOAApeU1z8jcrcpiJTDs1oJQtjabgqXGwnjwkre/nO8LeTm
+YN5rOMfC9M8bVjG4dtxDZbiOWJ7qqozMEgetcjMTD/thymVjIxtXdZGsKbAH7n+
c0L72L9d6KdaXk06J+PUO+BkY5TC0HYNpa7uqDgeUnEui/bLvr5RZUeFZQwpxUdD
KXOi7TeoxO3U9YsBgsYdDxaPSXRF2mQM2OpaIzukgC/FtxsYWqwsxpKC6aSBja0f
slVGUpjAZi9A6y0R91KMTo+mXrDagpeGs2BVRLXsTwGkr9UMr6gexKPyIJTZIMgF
AzAU5i2+NatZIXXQLr1DZphseE0gXpXD9En0fquGdV6ZZ9OoO8CBMaclyYA4y9jE
2WtAdgX10v7+e6kcX49fkj3XjwB8eKIu4dsEauOkQhpLFIRYDlLzjjIUZZLJpQuT
ApRnDtJYht3l2g4y7T4GWFkle9hgtLGlRseLukqflVCe4pDmkC/EAIhIrC2WvT6M
iPZm1lMF08pPrgCOE4PI0M2rj5crST9wPT0GYy70w+LFlibFrb+r1OMIxy+t5D7b
UHbtr77lplDIFJM3kZat9Eds6SOcuXDc+KnTBOBSuvChFgPmQbA5rf+HFrJuhpX+
2cy71kUCueaqiwYDy0INW+6IDBhmxY1GU0IHOHLOxGyvs8lc5xcwOT5/2TjNHSF4
Otm6NIqLY4yv7IacvwMWPvN/CnnX28J6gyZ6XY9PR2/UsjSRSwS9SvrtRSfLV8z0
I1Oi+1b/hbzirIqAoJDbe3xqjzhrlNXixZfqR/2Lx0rWdspewD/FAUK8eCl5/HbX
imlhn817zquLcu8r2g2SOgAWQuvy+K0aZJToPxj2age5+5pK5gkSNDgmg0NwGbM9
B4/KedEMxx/BC/TxNtQH3vuFDTatG1IW38mKntr6FF2gdjWp49peZPp2p5AqT8Gf
tO8JIaTF1eCmwLqzT/sImzXLRZp2fUbcXY0P3lUDr+nDL9wepUHn9VTVlVEK5UO/
a0AB5jM2tkKGl3TAylTH1c+7w0MrByTm5x1EEZ8gqLXNQoMs6AD3kXkMwd3uoBAB
3KM0AH86m5jBJSPitl/vmCTvhtg0bYvVp4XzRh65ChMkdd+IAgx1jWscoo9QVq8N
9qF+Zq/++Uc7Dr2GIMkt09en9SPzMKQvbRS0yJQpJ7TCyhvCz96DKNUkekeUX7jU
w6lVJGlkr2x5CSrLDpmegHrTNqUQbHToxjFOI3/Jup7RWUdhBGT+jntbp/sxog5N
ZLHLCW2yNmCmneZ3OkCK6wD0X+WmlJv6Co1Ry16oPIrdSIMjYhsMG/y27gZywIDG
RZl/fsXtw3Rvuv5yt4wDFRChAhyBTv4AM2HzCOkMfhwJGNRTou3sLwX8lCKLEMMF
TsBmijV7u7dXqYneYW++nIjI8xHNNurzZLxF7mOt0m/CsQ0jiZnmdPS4EB07GKDe
sq4nfp1XtZI88atcM8ljZ34Vwkqgl/dY/HBoFygg35wXajSH59VqoLL60RkHWHSC
rKVTOxJlId6CclG8aE9CbzoK+uDSW7lE1gMDPuKD5588keJi82fidNBYmVBA62p5
TnR36NRcBmLNT4pcW872sdaBmSWe3HbRkJrN6mmf/i+dE6wRVkSKOYuUPbOavrte
VipoJHL5q34Ouum7U5J8DGQu6KS3IOn5ZrraqXa0vZEhsXURSKIF7VHngpE0pTcr
tJAEzm9p6xu1c/rVys+KjIulqX++EHgHFlRqBplhAjq7EpXwcCw+HN66T9jJDUoo
0K3HK8h38AbNHCJ6+hyQUqmCHU1MmSziWVn0qR3wqnNOCpgqcS9ocMcf9x8nel0V
ObFAgcZ7NZ6F3XM+S/gwliMlesn+gXMixT53Si1omhi5yWeF9tIfrBWndNhHYD+J
8F0P/yzW3msYekqVnfJ90tfMsAOVEa3YQVNyifM4MWgWAUGq6E97JdT2WYceJ5eL
OfwAGPghJUSgOoD+xfyUcdRvPaqfOIeThDrKVJXyuVxfC0evJCaR/TyHdcRyVO+B
7oAymV5/F2bkFpzaL+7UtWLL/CRQpStXIWUZo/1c8WseD3Ltqyrh1jrplzE0lvfb
KIhnLkpnFRzog3UTPmgWB/Qp10sLuXJwSrKFpWsZuTo/3DNk2tH/P3uo0RQYKsP3
u2r4QPRniDKqZ4u0ij4SNEEDuGyf8BsS7iMQvF0wQ2srX/mawT+0YQlXVJupV5WX
9jNt/R1pU1e4hnsh9UQ4c+FubqMd/g0AqIXoatR2AXltnLdLrIYQdGg3OwLudTEw
G5VlRHJz0T536wv7ClBvOje+FywD4Mt0Nx3GKAsNnaJ78WtMLvZmhZfkI+z0JJ+J
xrbKgCtCrOElgY7hQ6j5eeP0oFjdy5M7+oJLzK92EoAyTrLgub3ziF0ivKoW2iU8
KVjrj9U+QSPZZN2Meraq7An8U4zwZxsxBbNrne3hn+isLUqKWHTzZksXiU3xLGMH
EcByA6D95zNd3zUaXebXlpMd20J61XPZsXDJEcukcdGSzIBcLs/gE0jHVVDBfl5D
uQCH/neraYn0Ge2TnUICQCaETd6m9uGEWt8xT1ZqsYnRW28nKDiXSwQHLTnHO0qV
mwN27Q4xd11kLK9pe13aSVbTDqN+TsdmKnVkRMje9wKck2fcKrKslY1VxaiSXPgt
WVHf66gZvdz1pUU6yDYMwPbUw6+5BzJa6Re9OjMrdVRw2WmdszuHP0B/XqSdhjbI
z9P1i4tTjN/7ZnR/EcssYLZ+SmyOrdgBr8PSlmPYR09MFXqUv0qGHK1/MGuFTbkP
csRGP/sKIGRvUvpAW2UhiwEBr6Pe9GzJwZD5fFhErCe1z0Ju4P0myDaVrqvhu9gj
S8gf498rMrSiqgTqsZeZRQT0pbHD5X9mK+Zi8tW2a4AWXGiy/Szmp17s5aWnNfDC
iGSxWBi6qeVKjEDwvMyf7XMVeI/o3+xh+YEmV+PaQaRoOixBl+Mt4SB7NcKR3VPG
NID0vD2Lk+7VhD+vnzAFwoS1pjdXXiC9jquNHB7mw2iQSrjJ5E60CSbsZQM6dIoj
tM/2DgxKJuFy+2Uq2ddHFzyCGw81HMn5LcmEyGDnM1CN3VD/bR38vEWyuty3VvMj
C/Yog/Bhd3a64gpSZZqtJzeYXcfbxPKhwedCvvqJOjVR5ud4+srnTIA3TphrbgTk
8favmRszqmBEFY0QxjxDzOiitVTupbsXBkn21MKCgp+5QKeAXOUYwZUFCVmiYWDU
KdfTvbcWNvfASSRjkkKQAV9F7SWx8Yj/MGVKq2MjNypENFxHDiFRzvBgSc0W6KTR
jizCEIgEyFdwWMMRtOkaC5nGU1tLdtUJfYhaI62dbxGdjdQcVNZiOootwkJ9HOhH
CixQg1AxzY8iaiumubqzEQalmv+NW8hkau5RyuuQNTC+nr5b6W+hJHdwUpWfPXDx
SoVsGc7cuoLTn+jEoZts2rY4feX4w2qOVpkn6r4JyHNrRBWxhGRNAdqyoT0fExDI
Q35G6xYsFWSJlOKdxSj1hLxy0WCKheLJHUciI2blSfvrCUin0EyB85uK88VIG0JJ
0af4XCIrm3QVOPo3K/w7ABMcIFUkJNT78S8shDVbxV1Az4Drkg5znrOvJopupKDH
AMkuuO6QpmZIMUf9eifd00JnzVeq4GlD+XxJTByro10kw2BE0sczTybzgZ6JfCOt
yhxlY1277t4JzMQhdQjU84jpHxamU7SoOW3vJv/JkoNGmYzuE1cw2rNsQUyKqnSX
ZNNRe1dDSNKXGXipUdDy9wCI0sdQRamT1geN7mrMDyYtXjbxWhlgyDPI6hL6nXVa
z9KRPGbseM5c0SOAi22TvuHY+eAHSGtjZYQ5TysyWwhInL19VKBqZpd3h8LyHFdA
7DQqT2lAcWVGTiHUzuJ+xmqk+BzHxirV4Me48/W2VhZXBnEZgbOx8ht597y5Vcmx
tt+UhirZg+Opr4moKsw6x3OeCPFYbLqgBf3p68tdgL8oV2QjHZ1o7CiVFguj3SVl
DWME1g9oJX4I8iAwIOfgfbREYdSjBWiV6wa0MOOJdkjRzpPicDS9WpY6PjEPntDq
c1bVtfXaQ1FNb3rCzRCHkXpIpjeZDv+b/0SkpQ+9tawfUiRvYHKT8ZRZEW2lG87b
on6uSScI+8KRDyqYhaiSseXdVyqRGwqEAdlR9JTEprnkdc6a3dnb8fn5d/2AW5Er
Jwyct8P+ROkSJTlgjZa9D4MkySAO4Dc95BdRrI3N5e6josAZm/qyO6yAdtT0MZqx
2qzDugv4ISI4MVHOOEgQg0Xe7OMDVm9F63Cxy78AxtZfrK/uszirlwBmDgeil1Ba
TyCxi31DAqoXbsbGTs1ULCSeG2AT4FSsewsK0Obai9ZAKNL9MxRf2/Tgz/YUj4RL
Agh3NFQ4AOAc0koucCvpLY+w7STrgt8knrwxUc3bxTeOQpgVIyk7xNJBvsRaBepT
feuKVgrIMu+zaCrmfFfO9HdJ9Nh6ndIENyAR69r81ew4qDDwxMk8/16r2hmoWLoE
DBXle6FpMvZFOrK5+UBU0mMlwXSAYMWtaztSVFXluMGMOlu/m6MeXETGbdi58e3y
iP9Z3Ju0NV3DN1HjZuiiHqdQqb+NN+aSKgJGAidDZWTDM6zv1X2BOyBJKVphiL0B
cHvh5fhaDHRAbq7GXCxMh3BN/QyAE1QKYR+tZSdsglcTXgXFtKEi6LwcHM42ZHfp
MXgp1Ca1XDULeERF3knJDWdH4B8y8q0Yu5WHgjK9QV2rMZSA5vUQrsnd0AnxIJQr
hHCKviRWBwLVMQQ4k3C02vEnJ47lFHb37n7F8V4jot8bAR9GWes3j0Bbs/knckbL
a6/6otp2jMo+2BXPELvX+pqCNfK0lt74pCOjtnYTNZgbj0PRIc4Y7BWhwS3oWgbh
nrvHMkkCxCSvCQ55nnwr8iA67kw5KVX7dak8ML0ds4cpNsnBU3uVmsoeKy/uRYZp
XZDNzx3EcQkTetljY3DZn/46eMkcbs3dCimYaAFOXaCnNzdmTJw/bEmZ+3s0ht3R
3dNcdwshOj4hzWphpR8rDlSRfq5pcZWujJXvvnyur8RSUtE6Wge72BxbRjVlFb6q
d0hCTJHL2zsGOthSSXraJsDijp2TQmSqllrmBBs6cdMeQ/yFQzIFQWmFtvD0FSXv
UCwhm1xvuaVQiPn6hmS7Gnn2usEhJxcdVi+fTtdftdpS99H8amFPaqQpzItxGFsy
Rqp/SofkhnsEkYhLCb3p/yHa9Q4ZHt8W7kutqwxF1wHJhb4kRi31ClVF8UcBzQHO
+ooHPQ8p+QLlDJLg/O1LJHSZx5r3YPibpKfEa5ac9EzprvstkPRDMQMGryTyeXS7
+ku+3hF0Bcah2JufDKruFZ108XUdEQDFkxuDBHHxJe/vvWtLuuIKQGYNE0N1+45Z
2Yu7OHTchVgl8UHPi0GfNsDNjdHDFlsHfbKmWoSnOwpRKCptldInj8KsrxzzcZRD
qTo+Wyv9vZMZpmFxTjGtfueaDikOk4DV+t8qtDOQJ5v1nKOl4fOxpbDB10Jy7yE9
6Skp1CECi0G6U0QBwoPXz4Vjh8Q2usDeTCm9G0MVK71JZn/crndA4m3RtJRPOag3
yvTFVwUvcJLLFEO2BNtbNkv2M5TfbMgelf1Knl7dBd/zLPaIlT51rSgkZ78ev6UT
Jy/bNaypo2TmxGZsnLM+Wto9/V0b467iDeUvKsCAOF8eYEPNFHJlkqflyXwm3Y7G
piqlqIqEz7uyVOSuSgu4jXbo8Dniu0QtcXfauDdTronC90TJZL4h4zC3NE0X473E
dn9mJfu2mDe4sGDx/9KJGZ0VGjqeJMZlOm2Po9y6uIDR3EA3Xqlk75Q0NPQDhEqO
DEZMr2i2sthKq6y51qMf9sWprlsqE0rH7tFNkRyB7xS+oxUskGpO6fa28Y49hpGI
Tfb5BvT95awkcoKJGd98cXe5ioZ/xmXf6BhntmxEJS/4xuIb2XRu885ZF07er0qD
KTY6RFE7NlS3ypOrS20z0CN2nB92ZuZIBN86yx/SZ+nMaK/eHVB54+ceUO68aLPR
EzUpxCDfvSVOcKYi1JMbK2pAZfWRy/2q2KrsKrFAShLtE9f7oMLyG0hZbc2jopqR
xHtzlfT+tD99oxQjW12G9rghszju4eTXLFF+ngVfkkH0Xcf3UbMMFAIUxP6FVb3t
7MEWvu6J27ebSJgOMgeuAc2PdKK3rDxqpyaO2bhCSP+jWVoZ+J+K+wYoyvI//b9o
mHhXPSkOsJNHg86IZBgnsZ+CgEIqCQuYd4O0UCgPRFqToJfUbeMwtdMmTyb8jjat
Iin1L+e6iTGE4jAjJuu/+O1y/4NYzpjmsjg8n+NDjYGMrGKoQ+H0nQPjsigNVjUO
60eyvdS17Q7Ntr6sb7MqwDmux4QvsBZ5uqcUVHuCUs6D8++H8sGi46vVhFiJIWz+
+GcazSyzeiB7XC7vYLZO3xrplQhLVqQqT1MUsMy7svHwllrBwbsLXxpTX5sO/PpI
QFgJmnoTtEnRpRIEGYAwSMwZj5TVzT8xqqeCSW9LKJqMEDRxewbXuGQOBP0iGhwA
0IidhNsup0aMOdy9NHGNerC79ty2EdnjuZLWapZ+lJ3tsWivPeVqfUCT7nmx4W8m
yVurU+9syF61M1LCDSym2ojiEJ2eQS2FCnB9QxMuaVKtwjConzbvGzOA3HCiQYtt
qQbMwpr3EDESjpfBCLskfNl7rlN/SyotUe9tnYrFRA4igJUISvm/0wJT9IECcHzt
gboxq0wjvhmnQHg+YFZxflCQTL2bzJrY6x7jNcwb8SOQYuhghOAuBFmUmHr212wv
Ui+MYVSiTl1aKX3gRFxnx5gPjysbs+0JBAQLKIGUW5x5RGMvP4G0f+LjaTktSgUc
rNdoj5jinpx3LhFOyF07UXiy6E0d1EXvpbKl1+GAL4iOWl3A/igR556D1UA7UbA+
0axlJM1joG2eUs85bxZ9lreTUHNlSXhEAjHgo6Z4Rt0katI1nukzvYKTOdnq0NML
kjnt3DOAXGRClMRcr+bvnf1GsHa1CEwAWD+CSI+7PRlgYrCHiZEmM7RuhJ1zLwXB
jBfSe+ZOsr/4WFkuaMq0j5j1kCRbSOoVPHqASQIrqcBy4mpYPtzzLYz1nkrWxLam
oqZEYa7HSxavJvgVn+KbhPHmMemyXjhwlThUNKMxqYWhfV9xUTT7joL7kkbxwNqp
HfZB5Wis0bnXQuMW8hUX3ExMA2FE1eIdaozz/IaBKxOZGMf4XMnO+6l/ewANWPRb
QkFVh/8b3YpQ01qQ8Kf3NKOLlS06+Cdv3O2ZLvIZ4vC0VVPqLHmUcRS3Z8T6B09b
JbWxCLr0M5VAxbCKOEu/jtZ7kUrgRjSCLGrksskzValkeKNfs4e+fkSLMikfA7Nw
Ew1ckHaFdSV3M19lBYYGm+MnAY9+U982LnKX8FhZA6IJVHHcE119/Z11vAeoovhD
+soy62ZpBjYJ4w+GGF0IG1XDkuW918LwBk32NDrV7y5cZUgVGs5MqnSV/Wvag4cN
5tKfyns1azvSCwyDsgWaSF7OOqYMJp5fQ+omkEA8AagYa9RvhgCF7/6M3JPr7s1r
usVj8O2CEDIjcz0YMa8P7aEn/L7ARVeZMNtCsPhqMYgwZkMnHqSyyX/kU44e0iI6
p0ptVSLFlyO4nNfck/DwOyGSrcfwLMWgFfEm1rKc+5R3IxR8GbRbVJSEOvCI1H8r
my9lcDWa/RRnRLal3ebS7JoZv/kBxrQ/elPfyHN0MiRMEN4xGgaajyvQDzA4P1Lr
7n5p4jL/zaxSxRyWHH+fhCc5WG1CetIteQThHeqFq7gv5gknYdKj8fkwnNI+Tyqf
1pqjJPqHtWhGFNKCvh9beHMlDVMYxF0aLHJFSlmTK5NEofT7+jJJ8oxZ4SubWJc6
HLw1PA/94m3WVQIzuErTtc20LU5f0zcoV1ta5op0s3Ne3lA+vdzOz8etvvFZoDoy
fpTYVrYNEgTC6eZ86xi0YgsCredOwEJoiwv8lHLSBL9/gLVJPCjfg8awImoG0IM6
WwOKU6FveuGZXxyW7NcHvNFRNRgQrLOFQ+DSbBb65Mdey2oTAmFFyc1XpuMaIigJ
23/L/161jQ8G/ccWDjXyd7i+Lwl02IrP+uyEV+Su82SXlJc3nTzYjBaVImuyWJvt
VrFpEJEnRmjJLXkjbYlf3El5g7XYddJquuaOLQSRQXJm6c9bWsdgYA72p9jwo4k3
+IY2h/k8RzGVdyyAnQSkzw+uquysLEUFCuE6RrrYdzVWiAHqy4IFPaSxNHd1+55O
q7mnSL1ycrNFd8P8ZhzkhX1VYp3GzGoTF2MQ8zZT+CgV2kmjXrfwguzL3TKPB2db
xu3IE5lfK/N7lyn297grKrd95w5GIgBwqOqUZnuLplD38q7taS9cyAFO8qP39e4U
m+Gg2dw8T3Q/ECfMBc4tLHdBivYPNa8s5UL0WD6s2bBAmqUzJmEYG6E4K05BMBfP
PdXfA6AkSdXo1B61AkOtyO48Y6lD/AQc3XXpMTC5c5IKrEAi7BCY6cdo9Cmugg+h
hniNBfzfdP995KmQiqfE5HNPRr9XJAo+YJxh7EwjL87nr+/CSqBtHXTn4nTPvOKI
SpYdpVGFvJz8QbIHqg9Zmp/BgM+bfbRKmxHRQ0UCM+7J3F6/WOFZfT2o4DiZ+s/e
o6PAkbMs1cTflEmpVOLh0v/mtpPdXYDf2zjFHneGlK7XuDHQqQ8n2xoCenYy4IyR
aD33dQRBDWJMYXxHNSMR8IJ4QCT5QfgDozXXKWZyjIJNdOIXe7meYOB7A0mxucaY
poDI2jmYl2DMT55XrI+pMCmYifhgAShTTxskBZoEFX1nxbK9Z2a4xFTAQH8p/68O
e3rsauAm3x4E9kH5wqDkMXmFMIkUUSahSNOG+tByJIgmSfAT2lbY1UJWigGKGiwI
tqUhF/mfrD9GW3BxfhzkL7m5kU9dAThIVPKrNSzKweGQk9JZ9aYd8aMgYUXw6fqz
TVd+YgUndWhh+vhRJnnEY17M3X9vGu9awwhVYn1bKuH37NoHum3KssyHO4j91PKq
uJTwGa9gRxQYvt5/rVTMEcxS992ZBQCwumvkiAr65oad9w15hrJt9t3dUI4PTVUA
vyxXIwk7751ZVrYjbJbEchQf3bQ3we03GqzAp9ELYFPHpmDz4G8F53HHQwtBmt49
xZh59QBxll/icG0+uiP7MTmg7CkKHgSbmQzlejnnbmlg0uuH5ERav48sY0S/ZkBJ
dZkkwT73IHiwl/VxsNoF6hTfboMoHhe+hQ2WO3OWtOvg3TSEf3BVNJ2eNldO1yk4
zvJ7y0vXcDQj0WMBV81HutgcAwNMIFJOaEX130wEjsWVVW6/sa4ljLy9UgZOQS1J
wSmxAdGl//kENasH8eXvQZqgQHdqsyI2qQZpOK1K7pOzr8t31MRx950RfX2mBNLn
Yp6EQfV0nWvv5zjkedernMrI0YgjnlgYpr56CulIzHuRdP9RLtw+0E/GKABD2txW
EqMeIcSw3Mjy0gHiCcgrUb7Q6v1A5791w0M2j3F10rRkT99gG3/+ltIvIpLBQQtu
2mI4cXRmHgWx+UumTLyStPna80yB7+M53zibztgXcWSZEaNLtFABjUWGXPoJN8LI
c01S7lhsiPCVowces7BiuYVKnOk6czrrkSyyYSVzKvIPfdpbMRAhZHyHpkQ5MW3y
Ak903wmqQgwvjHuTBUXD/a6vApXrxq85SIDZOSqo+JwHpVbPeTrE7M1pyRryQs9R
nF05AcQOIuSetsoeBlnpuLhwNu7cxGXPL8tPa4IZ2Dj4Dom5JKX8abFjKlbz/pwM
D0l0eox0IO/pnFvx+ifvSkhf6MkoF/+lvrPW8Y6qljP+e3Xyz2PNioHdaJhaCz/J
ANxdcly3i6e32vYDFJL4iZYat2qBJhYgJQioQvCH67DkqXhnu2us3UBPXHkSyDh8
dNk/dVxEIaWRIv6ilFg0nuxgktH0JNNLeiKknl6Ll1C5Rg75QkSWfb6b9qADesFE
0rD3sLMYcuDu6/Cftj0Rb1glcgnLIB2+YfMq+DzdbzNafBYCEypC8L6i6B7MlVJT
H0iMGsyUEOXapsEzEAgA7HJ0lb+pKWNT6y9uCk/mZ0ckrd9rLWLVlD0m83JABtXI
XEXLPJovYwI/JwT03gU/sMR118a0zTSKiZgUAmLYVEpYGSallCRnWP58z4EVpHOv
k2WjXiGnocnN+Wbzn69+9U46r36xf1wFn8VcDrw7lEdnQ9G/6JmQ9TilOb23RH3K
/Vq5Km00m5smgxV6NVhBHxuJODfvWsrRjoVCoJGFLA3FxphDTPSZDnk4O42jeTlH
tZuMvkC78NDM7P46jMK8K7kPzaD/QlBwIOCZBkFd0afNYt9BST9A07/Zlifunvf+
JdCsS82ou589q8Vx5S2Z8zEKeaAoSJyQPQBIshlMjIgHQmk47+eiZK8pfr05ciR+
6UBiBRTmZR1ow3XVL3iZGvtEWgIdwnS/2VntrBJ/qDt7MkXrLInMM+Pei+2cbLV1
e+Gipeb2QXjbvz8syuN2yryOTGT/vMjLoOfDLH9TsZYLOicn6At54Wjwu7DxbEgI
/27YQW/YPlYYEf8GXvQfVTQ4IHPQ/PG/g7DfwxOAvSYomLGOGi3/IPtuaD8WgNTb
TCShrSxX2xD8osrh8LrB7lA8xTUsamhqgfC/9X5DekTp/g5CNshu5+wlJPI7f3h5
M9LvYHue6Utj0RsTL4Rbebqgds2uia1Ty6akZlI5ZcbeRFsZEVr4WhMGOKjzwWOi
f7N3dxsBCpKn4ztc+WyyvAvAa2NzyUGS/luY0YmDoLpP4FO2eflEk57XRH+2zxzU
XAFiZuHXY/nVyjwckjGuUzAUwxk0q8iK3zLyLBfByaogtrbDZIDtmrYIF8O/grSR
5aQjI4MfIHaAOc2IHdnEYGSGAd5Bb3K6H5PRJbNsPMQSalkS2L41Mw+bkezym6HZ
fUPOffk1UwSsD+4NWZN/a2LRSg84TOp8X7qjFsS8MuU8ZEirzcNSyTjLqS3YL5rl
b7SB9W88AhDSXWFjkFv8gYY25LH6domAyiA9GPdQsBOsyaAEUzBq0rdvs+cxaTlh
grxQHqvHgi2+9lyHw8nGd1ZQ15/UOFIo1Jn1SkSTj+xLM7iiYAg61C4gWUQ35m5R
ageiwbBtPMuIOGrguP8rGl+Ic7hBdLdUw5vpVHHkum6xYcb3hH6vfJ6qD41GDC/T
S/gJh0EiGkG6S6jJNe3MbCBtVPC0jZJdT3DoyMuWA5QHyVgZyamFDcT65r+qKWy6
UtTgmRzRAaLoBq4NdFc4Tp7GNOdmcGiUsWayA33sqTKGlMvTpzHrj9huaJ2QlMma
HSjHpKm6obNAQhBXcXA6YfnbWLHnpTdNkhI6GUPDtJlI22yNinS37bswwScwlXnY
DKxhWRSqSjlLNXQvmAVvNJRouUCwK4YOr0IvGfuGof+A0q3i+FNypHf9pBm6ZB4p
tkTr5GMqPGdaamfv2RZBSUKUuhkXrUmfRVK2g1e4AlwaFcHf0R9ryZOF8/cmzEYo
q+OJqxHG3owV1cxdiZ2z4uYlH6o3E+Y7CJFqwbAgFmSX8PceJvX/GdtBvfeUalLP
VUW/igLBiiK/HK09Fbqtd0IuTlcqka6NwgH26lL/hWmg2c70wtmf0VpOwKoEhLk7
Q4zjymvdLgGQo1SEAy4LJHUrZUmVK7HtAI0eQBH3BmioVHG6cceOsRFcymidsdxh
WnqVrgaOuDAArig9W6izWkNOjM7ZWyRtEDgNuXH57cRlZUg7IPJ00cWlgFEivSpL
puNtgoToVsLlYlvTpIkveqsHpx26pcRq0dyKhMNGZ9YuGFnz22eKIHYo9B3oZ4ff
iCtRHCmeTTv66vrkdyWygg06/uvB0RrEFBspNCrSNM/w4GOTbeb/LsOE8kjWrb90
dXC2HHqWIUvK1niOs/oilQdZX/qNUxKLxTfi7ecLd745x2EwIvkP3sDWYrs/9DhF
OAdp3n8Mvtj8XFrfsasY2GhblQX9p/du/YTsHpstE9w237fHjAiqtRdEZqUBX5B8
pt/Zirvf9yEwJhHxB1005Txv3oUVJ8v0+8Xec3Xov/msmg4XMjTBswbIl+MJD1GN
gU5lxgvXz4jvxduNNWX5+Z0zURhtIPjn9C54qMxSGa3782DKDrjFmV3ysR93TdYv
Ojzi3qJWttfKyC+T0ewhVmyYZLZQTSHhi90pc8+WHhJvSaQRPtMXB2/BqP5Dzp72
mahYTUp+k7MjsXLXwjgBcAcl2XxYa8LP2mPS2MU2zM7Arv0P9P252KDSvAgszxyt
2+EQGFz2HlOzdbo1l7pRN5EAFi9lzq5nQfbBoLdPcTsiyS6aElEOGI+MKKvS+iee
ppBLT5DY529QKmpZ3qlXZ5aPt+3QL+lJIT3Jt9R20RWlgleSj/rhk8NC/hsBJFjH
ZU8b5GbuGTsBkbTv+lxbFI3i+3bLPmRxriJPSHZWwxeRVkB56jPDYAW501zmAO5S
hhKAygnG8Us+v73PfwQCjQ3VK19NdATNAK1Rt3qu6LlS5W23yJB34Ik1hIHK+c43
frzELYaepdinGoRxmxPOwJxDofWRxE44PsgZFAy4PAfiZcmEatj6VFLGSTHCBR60
/shYB0J2T8wKXmpStYI+Sptz9bn8QhZJULtz7IMjIjLNeQA7IE9PgMbxOjQayiSu
oIX0W1JG1l8+lhBD6tpu+njVIGtkhYeOSS7X9lanQxS+XWYnAI4fzEHZDdwAyxaz
Ao4+/IJuRFyP6KtSitBeN5F8NHd3oX2vMkkXrq0osIVhUAw4ciFNPl9vQGpezOy9
gGPk1ba12VTQIxV25S54loj/jb+v6rnyras3Yl78hQKQcAkh9tPW6bxR+EuFmsWR
ZiU/7iAaUGqR8YBQZ3N22YpTM4XnIk/6Oj8AsVenR85dkU9zxhC/TSJ6jJoYu70u
0M+os1YGcIwsdN8GVHZNDvXoeRIcqGOILvnamdbRQpPGdilUV7xqaKFqrk/vXiDT
vijvZA/W/dPTjvjMrGmeJQjM8tfy2sEAgk26A0g9NTSWS4omQVsnxKSS0ypqxa7L
1G1vWH6W0AzrHFVC68NIMJIWHy1sC5EMDIWx2SzhxsXXnSEpY2nG0Z/4m0SQzrDi
ew0ANwZyor+hlFfHQJE3ZHCukfeHKSzD4xqr+YgoKd1iEuLQAO95iO04P8iLH0cU
tO9Dq9kLoM42mj5nYKnV66arvW+QDzWoDz9l4Izr1Xj33qy1HeENZbqpmhXo2BNy
xyzq88iMI8lsZhrD80/24qWevrqck/F0Q6TgPdk02aIQjFf312eqZkstJyiUq8/W
x9CLhin+INlvlb+n4YjMYDOTfKDh5Njvv0Of4stjBKPOULgrWVxbmnQDSfLsBKoQ
yQmdvRyikw0e3JNL/youW8ogVP2dnYiCWczkVHcdLxrbMtK+7eW52LHWOi9K+KUO
GUzYEyVRrYjqyTh594OCYD2OZmlS77ZngCAPhyu9BPKij+I7l+G89ssRPnVL8Eck
Wtk9TDzAaKI2GZlFXo4Ev7fVX9z3mP3oNpl+GJoRrn3OcDvA7vyqJHfdNEM2Bw4j
KOh3oBGwFRv01Swng44mvS6eaTyQDVYqNyueLyq63l5fqO6IJqea7fMjws/4GB3T
bDiRCcG06Ay60VCUrqJALZpkN/O2kL1iU1qMqtdq/di91P1rW/X+ejdlu93Yj/Sj
8mgTa4oaMA0QEaTGJ/xfLfDS0pTWFcqOhPGDmSOGNt5l6wpV4a2uVvabcecV3tOk
CPntj0D4BRIP/gB8ilWMXGF1ldQ+nEjis9W0wmk6b1XPYkw2tO+KGOEydvNZ1Tmp
p5988sjuJJA98eOSLot+scvirSs/kMu2r35f1laT5Iq1luDQxYqckluECyjx7p7+
pLytlCYw3eqnwu1zcSRFdwiQbMd0mADJm6thyu05W58yYsjtPein9Ek6Ibl4Fep8
tWMNsxPXOe76Ae9yAiarsjPQDMp8PcfQvXWkAyzhF4yX6Oj/0M1jAeCT8GfVHF9o
LmFjPoXULmJutS60DxIbJ0ZOkxlft7csLgpI//0dlkDUpfR9Iu86Zp+6GFkzVpEM
J7iZINcWEyEdBCj9LamJZRPnBu644qqqC1cbxGDcECPQ0atGJP0ALCwXJ9xrnUli
IXgx/Nru7afOr2x4oNmzBvUZhMvQe8KPlRpeJQPhC65IH4/iA8HHLpxQWf9uStc2
BYq2sbIyBLBYd6AtMrpXtDjq/ZvRdgI1cuGACdviGUbzxARzLLWZ5xRUXuT1P55A
boVXAKPA+LjK0KEf0VCKPqwTQFa0nJAySbGvxOg/7xO/wEartsBixDu3rlIk2+LW
uhJ3OG5jc3y2uSGnzLrsp2L9rZTxrPSAZAoPPCchKexi0CmTMIGSrE3dqrOtAWjn
UK/9OFTwL2mJPI9pZ65ZwjoLSHO2RDUfJ4YKpB2AbjTmBnJ/J0DxMSSpeXD79h/K
Nl8jurCfNUaph4+5XVDpd1zostuII+PVRvTeFdq5ySKHDXqdDeINbHNoKv6qlD7q
WkMXewHB4PYA8y/yPWCOSmzrzbZYtEBUNqC5SvCl8CLNoXqdbgM8tCo/Yq13Noqh
OJ7V7qdAGROcY7xEW4CutbN7GtMQrWoaeQCEAImAO9MeAg5XAb3QecII1nn/1S3G
DCxLK2T+MN9wZECSUQnjt06W3WD/eTABYNDB+/I0lyQbBf+JKn/A9NurjRzv5glG
rVTIATk5tABKtAjQFl5h6+KeqYvJdC8ptHG048hb+4B6Huad7iFFW1gklYnaCi6t
XBjzi8BsPTZCqwpsuOoGZZhoi0PGUAyx2vsxMzoQtE1BWbwODr6dZRBqkAI+n4+i
OYNnJ7AbQmPDKVekzvKHJuJ/U/uThU7JLXvsDlRyrLHPGCmwfWWdcoFOmEXS7Fal
tZjaiOr9AEvRFIQzeDDiM/arfvEsu0zI4D/ybY6zD5Qk5aAWo93dVKZzQKTHNFtb
KWVlCFyDZpOt2tlE1hOVEJwVsgabs/leLcHSDdkTjrFFMZBMwDHEV0tdPjNoyOfe
/xxLaVdoFRfQij8ZMmefczchRrQh4T88I4QHesbpa+3q3H0oxCa/b6PwZScxDYWi
RDLCDXmD6O8TZwt5nr2o0wKGzVFfE1Qx9qZ3n+nRDYqhZbQQWk7GSRV/urVETYdg
7WpoCvrl+wmI5lUueTp9BH30Ejkwl7Ipy8SIRgH4S6RKeMJFeaxsaY5VYcLnfU1S
+iBgOfWPznUKY3qwFnvD2YpCCqgzYXOVtOflqXm9LxBR6wJPptSfo1HDY2tI1n97
WbQBmcxE2VEKi0PrcTPouujpDn3hVLMBN2RJ0H7UBbX4PZKUBcbc7k/LSZbBImlI
FDmvTYfmv9I9+uPdIqMamqFclSzKzib8Pzo3RD/cv5lBTMk2UtEmy37VOcUuKbtg
aKZxqIaHIlGyS0apSCeJFozDXscJTxGVjgc/IQnMrwYPYWDLVPXNiiQY/vkx6dus
ZujsiCqoHluiLMuT8yDlLQcwVNN3EaAwHSkZD/7QexaSo0F0zhzPd8LwXx95/fNm
2XJYiCMnQrcofF2dKq5BoR3IXv2zXdd7r+lXsrIJH4u7GXJJbsUn84+pNmaRDt67
3Wjkm52cAPzn4H8z0HmNmrpULOycmBmKFfxiwCMVHz2hz/hbmK6FuOeN8VRuAO3K
trsRAlu1wELOTRk0Q/JbKpfvddDqMVmuvLmpGHNRIvNKDliYJ/KnF1Tzlq8boSgq
PXBV+mJkpKdo2Q4lSHyeM01tWcMgLwS6vhJpD4y9vRaGiUmAMYldS2hBqXKKCVLy
vH0dd7NWWssTbJl2jUkWzxHm/sIcCVGV6L9VQcwb3lyjvXYC4VZXCW5zuKnYUVWT
bPX/SDg+9v4bm8W4Xv4uhSlEg0xIvQjvIePh0Qoz2ilkTUoFVZAsPgJlshAgSL8Y
0KGQD9FYEeRbIkEQyQ6AF8xT+hzjSNqtGXOkZS7VKmBKbnHHvqWkR3zsr0gIpIL6
4PlXEKrrVabM6ZqByOS9Vp+7z3vXYOgy+KSY9/SpsA8DX05p1hjl516rahqn19J8
zFMmGKzvAOPsoS4XjIBMi9/7+jgbCjSQvIv6UR7b8t++wDk5GY2pLiVuek56f7nI
zkj4jV0QMoxWayRTJsLcf0KIXRFzqa/QyXGQRd1GKMRZsz2hmyv1HPiMoUlU17Xq
pT4DibzUGD0SLxsSrqLGcO5r/rpdXB2+xFM6vLYVI05lvn8GDaGx8mixiRADMkUz
x6plhy75VOs8Awwb86j/XINbYevT4/+CO2B7X4vSWrPkkQn9GJJGnGjEC5ul7y53
OkTUb8utGY7uz+33r4BVitFUM0SXea7hQ20jZ1j1jPu7OTz1uHTU1NSnUnTsyOxv
8BeZUB5H1OIZKGm4Jn1Ivd7LD3z+9xRXOlKqoOWNViC37mfbrVeajPosx4BTBFP/
5GZifLTKKYQ5KU70Tx/5+kqFAbCawyxNfbONNl9mJOJAEcnZaP7lNPiJ+BRTOoMq
ox6yyk/XzdBvGxQHWwk4Ip7j32sqJgSXfdXDsoPo8447pPQwSeGWH4HkOhtepZbO
u04WLBgeI+LXG+IB72POND2YN94BooA3zCe2uQNR5GYg5V4GuwbYR+wLVRbodFCk
HJpEdpmDymr50ZDMeQgsfNl+IKTXih7U3T+8Wr6f3r9ohinPMVSzhtJeE32/tNhY
op1QILNBjSBq1VCdIrSFUTkQ8y7sbAbxxkzYKumaBGGM1TE1n8DUFeL4qcc4WtA2
/QuP8d9pXfLn/9afZpDMq0yv67yWL2H6FQZRn8Zk6XzSgjxhkSqIptQvZ8owcA9+
8xb6Vwhg7npv1/yGv23dPZy36YSfxMv2R6h2dnfMwK/a5ucCp1jWP7inkrWG6pTP
eoPbY2CBbygAMbShTtA7ZG4/NIfDrxKgcbLq1IiAi3sixBy6VjbFoUGSFiy5pFn0
S7N7p3CdBMOKtw6l/+mhTHX3vY6QQap8GW6bymf0U8Onw55xE0X0H6HWNq2AisLE
Jzt88nVr8B0/uFb+alIybBUqBGo7mfb+STMgC0WTvGen6e7HA1Ppt7I2nGC5Yv9M
7AAYutxj3dicntHMCkQzLs2FAN403v/XWVIU/ZDYSLB9HJsalSlc9lAqhXzhQrFM
9WtytwzSN4KmAoB/K5njjngJ7DwVfFHkjJTz6Dc23xY4zLPAupmNGY2N/m2iGnZs
KRMCPCj0qGLaT9lpYSW9xqKJjewJFa0R+uxElyly8jql4TtKSiH7d0RDOT1gjceV
Mq3l3LO51ZwWqAHDmGOPxyo5KUYeejZRbpKH5qvEv66cuGyZthIltd4BL1fVLSCr
1rZ/xkFBjE32Tv80kDMJ7bot34etArGXFvN6+XdEWWbnxhtxN25R/p9gYCoQ1mPf
OTI9b4ZsHwzVSCPqXbDPpcm8BnivvufdvfoXln6LFiXZ8l+lRzLnnLEmA6V/VjKg
8YSfPPHWyEWEOAV7XGlTYU/F1x2luFtiQJh+sqFPiOLc+Vw171yHOn8qKjQBeJRo
hGhIiW7tHPpaIMKHG1hUyi82AI07xm7/aW2sp62Cq7twE5l23gU/bkmfNHtjqYQa
DTvHG6RW4VkNxhJ6egI6ZqNBL8qQ7yn6nVXL66ahPnRaRHaSSdYvvc3eQtZCxjGS
yIsVCKYZWJN/JR4ajU/rzZjW/wkP9fPwNhS6RxoszT3CQFmNL+jKAMRhHxdtbOmQ
tADtzMTK4YGBuZLpsdOAry32ImRC0ETs9bs9RlZOBmyyLOYe3eD6p29w482mGSPF
QNpPlZ+jYjteGsvFapts0L/uHol55X0vyviY+vipTnccdCX5Kb6V2zz6kEtwYuhj
JwStIHGUcb35hZDN6XL4vyDlGQAuY5fTFwHCuLzTVGwd4mIudSp2PkPVTdUGIrGW
ynL5c8r9061ITb8icurv4XKu5AhcgGFDK2+QgJDSmq7xbHdk3IL7kciQ7VvXUbrE
spEpobcJVBYD49l2leTMVEz2YIC+zDrEyzAv6nZP1SPdhcpZMmk8IzCGXFPY2fT8
XZqv9e31/dUKQv9SnAWfVjKz5sdnsCquyKWV9EaIXhH0KKqTY2zFzTTkb5pLtWF4
brMIx+QnyydEoZkN1ZB7d0ymvGzOFZSWfWdbQ0oozBizR6+HMWrIN+9zl4/t3wgj
DpEE3ol7nkBX89qljkY1dr3x3CXXWPuHSCN5X97wqmoZ3ODgrHogLolSF3HOVD9N
q4kp0ibt+cSItR/FSC2vZqsH1PPsTYlbtwEHZoq9BELsespikBMNcHC6SV24nA3K
9NeaZlHQRz+gzl695Rjpxpa+/Kz6yhYCIZS0iB86yozclbHZYs864/kKgeaup3Gz
B8NyJL5xd4dcCKvTH2hZ3EY48CF360dDNh43S806RmbqKgOwzuoIcylt7MTpzYFG
ESpoCNRSv5L8aoiX91u2pZmC9xZGiUD47K5SWVqAG5Q6uSYc3WkRNYXwLbB/XXiC
/TQmAXrkFDwPIyqaZ4oBEAlGxZfinZp51mSb/Ew4iNXaMydxJz/jdNbP/Een8owE
YXp+4BP3QiaeA+dCHRvzQg1Podl5RNS9uz3tQ3KgpsIRhjgz9DGUyg8Wr1aY2BU0
5tPDzejzUF9kqhLiONjzec7ZUn3OdImkqAvmQpXAphWCc1NSmldvhy2MIiNJB3ZD
4zF0M1p2+CA7WDwAuNyoeHacf35cpiwfGgIuLb+MAZw3uVCHWv3VYwMPrB/OPjl3
V1tyXtA+dtzyT96lcMNJSyeJYumXDdUB8xy2XHVzvJPktIzXQPPrWRdpGaCCx+K4
qDCPAH19fAOUhygTgAvW/HPeInoZlcQEFqymMghwiCzzfmJtczzRAgdaRXshRf4q
q9Be3VjP+svMCUWMfa/KpLH0jnwB8eVVBBla1FkC0YlGsIZwsjPWzk29sV26kxiG
+uw2VovH3Sc5S2fTIAM7pGMeaWtHTAh7Hr+USOd/dpi1wpQVIdyqL8fU3WZwu1/r
/d4l3FnFgp0gbR4GQ0MZpwM54Xq84giPGL7sCpb6htShzH/3ZZTnoXIYFgGANw8z
JCavQP6/7nS7Sl65ktcx29u4C/VMWQIANl4UaYNSW4z4TSXujiz+ny+f1uIHurCy
BaJdKMNmXtH6FBTzPvc9Wb9nmuvn5QbEGxwb85dIxtzDzvCf+Ek5lML5hVRVQ/kx
6y1ce89oOw0lHWTwhsM5LjjYpM51/uE9hUW4gYgqdjFe0GnT7zzbsw6JaGaalA6n
x5paUAQHLj2aKfMWxp3Oh44D0+7258unkCIbJjBeqxW7H1ICF959mh0EIhPg7RX1
31OMdf6r7iqFSEimATUBu6p+jCA2cF7rxAlMt+dm8Ga1UQziW0fwtoNVtdBycANP
P5PD0RMSYJn6BUgT2naXGeGz6gH73syFntP1d8RFUYOvZ/kof8a6+Wx6t0PpQj95
YzmA9ubhIrIu9L6VArOQVaw2WGY6mSB5yHyHLD0GvC/aux4wQK8SFd6qP9eRkjR+
NDnhWGoSBunLxmR0IvXMQTvS670MsLl9KiHhVetIWZno7bPL/Z8NWOgu9Og2opFt
14i8r/MP7q9Mb67QCzrfUipqrlcH765e4R7iGU7ruynBgzgtK8dRvtP/FC6eG2B8
Vo7DXpOkVi37f9KiRwlxyPI3EUbVASFnjSsaDjcs5rdcJ3g+QmkMey/Ec29HNVAp
+N7B2UG+tXZJAPLza4BD3SplXYFLfqZS+S8NYkxaaFQSCSNyy5NrrN8+aRU7Bh+W
JQ7MzOzPs1+YQ2dxgdsjz6t5THv04gGo1SVHNOQ71zScqfEd4JbdoDP0DjOuqyf7
BymjuyCbiLpRABtigEZj1ktAWpyPNVISYqdfStcluhcD+u6/JasvgaBE2Cw5qBtL
OfbAqGCRpIG5fRIW7ERAen6pAw3oiCimkV2911PR1uxDmmw+HB7lrgRVLtC9NA29
c4Koi8rYFiccerQlMT4Kl7IeKeb07LPoaGNvUrxGT3DE1Q6vmbzKSjASWIxIxJR4
hCxSTamo/3rnnV2JLobuIf+D1JixOBDSbZer+dISgT0Y7g38gVmJdJSEAk+CO2rC
TAODRsjGbf3XHf51/RocDOjyu6i8ejEZ77yRHNKi/oFy1d0FWoWN8pbzrQc07pZV
IoHUxhrZstBOnCRF0JPsIt8eFjD/YVlj2FUsdarJzrpXv7Jyj2lQvO6vJPVL4R75
pogPjBoq68QlCATxgK45qksKXYU1WQVcYzZ5Xnp5eufHeY9KCf1Eo4c9OXLB9/zV
gxIXgV6s+EJFfT86+EULlAjLqrxWZvYiI+U2nJlm5c6eb15xgF6WEBFZ1vYjpqjr
UbcPMTdLalooOTHxwUdV4vWN5BS3aayfYRPvydWy0XmpB5izkGCrCC27VLtcF1oz
OuCMbYW5D+7zGJcl8XTEPAou0/rvVOaXD3e2mePqSB1VBLcdcmJbgcJEbIYUCcTf
QblyXDQ7SJ35ghsT5i6I35Dy5lBEyPFteLgwgY+vwMe0Ve50zmjfNXHcJ5x0uzRR
DVrs6AkQK8KV34U+gjeFeg+QNJxrZMo6Jhs1fHiNzZHV7srvN3NF/To6JQ/mGrpW
xl/8gXVhazKYn8gZTRXhdYXAbNF3DHeEtr1L0C07JZHqtZNsah+CoNPV7/XpuA9/
NxDOyaY5p243XtQZezml/71SwtyvwAbXGy3As9k22rErS/jAUUDiDw8g6pvsu+k6
b6PbrcZ4dJEKxBgtpsOx8w7VideqsMnEs47vwEXq3g0pbQjoagJtPcXwFoIzHQn6
+alR5iXcM0nLtnJfiDpzPpo8LxVB5ZogXUDOmB94tddRRGXV76FegVAloVtxjKac
a/S48g4VF2QLdWlSUImVr/q6NhY4g22GrOuAp089imKT2Pc4AcucwmEZB4a3usp9
mKOQXcS9iAmUV57V7/ui7Gg0Y5n7v6Nw9si2XVVQfvC9zlEHqxX7lGW+u324kI6n
tQ7mFY1m5ZDRXVnh377sIcObBCj0+N04XBuL4EWg9JpRzQgXe/Vssnae1bqP9zxt
wAEVrIGgbvMwBr4nD0C3lWP94SvJflLY2s/MjzJTKNyDZDfbdVfZJ8aqsnhwdTBp
ZTKwOx6/T6uXmsgFGwwJler5IUo+O9BsoHs+567BsmdiWGoCCHrjHaCjrdMrOAjP
byLjpVNJOXrbqA2gYdcqvRHE0lrWmC6IGwQGVeOLF2qRinZQx9XFyayfeZAok9jA
zv+nTFo2RYsqzlLClvuPTb3J4UMR0cmAR9AJrk9lQfc61hMmCKoU6yzYTvoBZqzn
gJBxgCwBx7iyEsPq1xhm88rOygCuR5XMH5cdzrvTtTWPnFUC9UVKL0mq7EX6xCVY
np6pE5iPvX+a4G27+deOR1OpCIgPpWAG5kSUtTSML3frRMhKjYQLgBnhP3JvluAB
rSROWxF4QDZKS9ZCb+WXS1KQUfnlv+MYujq4cHBic/ZfC9jwejFs4E37Pu9mVNle
ICS2HHgPzej9ej5vvqph9ekm6VPUpR6p8qDWKGvxs36eUgE16B56Of+MPTjKXvTS
2VP5BFD4VWoIlyqIoLOA+aVIb297vU1c2uhzlDk2KcNU2A/XL8N+yyLSpSyYwHE6
etxUAMyTahx8blKO3MLct0uEke/Wl+ezqCIFF7TFtI+V42lUHf+3dSbHSbdmQd7Y
zoL6uCIkw0N80MOjhcsEE6p54TFVIgB+T6a9pYe5+lKaQsB6uhsXE6/2jNhHZ3CO
8qC069LoOaxLAdbIDp0Z/TPt8FqlSjxlFOazJ6ezYE6rM+KiVeiiA5waUzcmRVmO
fqxTZjrawEahfP0REVmyIzm0q9K7QfBel5pDPAErKBk8WlttEd0eUdl5j0pCNBR/
lWPoOB8dStNLVCjA8KV26ibmN2oGBWakAeYeHlEt18wjEFnibaT/RZu6IEgiTfuM
ZzQJg0lJkPL3offOnjRGgvb/M65u8tb4BaTORisb8lW/0auPCKUeX61f8NilqSS1
c4vJu3Pg9z7TORCIj1M2gPWUV92clJKxNazqefrZlzMtDww/eihr8ZeeOcgZqzsh
JG6dIDj8iV911mnAlrbRBLjeIV20ipwc5inow/TAqF/6qc/Q83OTSliYqE+XTBjJ
IksmYrefCkLu9FNwuyqFHTLFKdDwtyaR340rZgtA6cMS2i9PbAHX0EWBQ1oS84OJ
BbkIFlihSiNbuwBY31mIyhnNAs5OUYuk0jYF8aiDgtQOtINup2xhbY/yCcs+tVhd
om5ySGty8999nzM0SInRhStg4Ea+gbZIUBv6M72pay46NzBbWycgaI9ZlPuDpp5o
xVutn2MkbidjQrz39Qh7ckza2YhrGAOv1+DbPP8Cw5a1y2WyMUI8le9ANzm4+2UJ
nUrYTBVeyf8vwmGycRbytkabx6oOC56IxwwMN9YGHlLHMyeRw9vNIQgyOuvO4Oyq
7xh76mdsa7iw8roXdLGGZ9ZbMmJttgQxOded5V+yU6bHBWL419Z4ysvjezd6I9xr
a0ioJELqoRqq+6sUP5sRwqpvI2e6khbo6wK96QSEs85sqXmdaJrmrG/xpiDTlGrK
wk9q35OHYFY6FDml529Yp34yIeHNkoDf3HMBqm49Ap8QrfrcR5/P2rdZuYzfNQtc
jA0xBxEmYjGhNQzlf3VYMQNO4dqWuyLIZ7H0av/A692NBWjFg6G7slu7MPejdWMl
Lyj3/7isrzLuxh8NAYI6uET38gq8xCzbW5W6B/Ao6JNFfFoFN59U/9+qTWjk10v/
CMdmFyfWNy0dJiNyhEmfzVRyk2LpoR2eVnbD0EW+pJum7iu2xU5sf37A3006AqXW
PDGVTSg+ABmnbbkCglZxnqKwA6e8k9qDW6gkGBj3b6vqantAeeippWPCspSUehug
BFnDUpQ1hrMZxqfJDQIdk2fJZ/fcl0O0inntmwc+/+8Qdu40qjThYQUqWEW7ZEVH
6nvZh5c0G8VjGiKv0wabSPQgK60Lhu3d+1mN9WGN9Gec0pJcY+BgrDGxn6Hithu3
8WYqtYKwFNxRB38fvGJrG9GYhP55DYkjVJZuKqNd6BgzLlzUs+B029VtMS38fxQ7
lJ8h6zWT1JUKWd1gcb1FUq1DoPG1AeRO1iSeSy49T1sTYOb7hDAtyaJJS68DEFi/
dKHJikg0x+Z96fQZg+1bYgBzClZghkPq+Qf/K7/MxeIlBJudFaFTXyUt8i3fPP38
99TrIT7PjpPRk6dARWtQZ+TPjhtfUXRxyy8+QfDzKiL6Gk4CjbEvn+o1BL172UTq
R9C/VKoPyP8sH2NGt5ygmsfWj/PryAwL6QWnW6jcYEwSdTcwNWBWNGyxkB5rWba+
BvnQse1HKec3R87qeYR2cAEkfkq8aybMIuzpAG1lJUebdw5iZLK6Z8lCYiEEKZVl
VigneAewzQW8pehvDJ7NQjqEAw8OASXOyhMdKy35/KapWTg88TyRTz5NM6BB/rmA
gbacyHHFPCO/OC+6XuE9jPm3g7nV8med8F1NUCRaGSRUOGr1U7wJlHxfjtbFyh0W
kYQKvEXxxdIrbykARYisAe2gJosYq9Dznk0I3KdKZ/I0HeDCdfR3cl5kls3eavJw
E6IKBzL1yvDvZlmjh1aj1cu+0mShDaOPp4Qa766AEyplbjTHNwttZYDvj5P3RgRQ
jyZZ78fK37SVoUenoCoj+UCkEEgU28UKovCsPqzkcPOAeGUXGLFA6dE706WAwwI6
4QElKl25GOCC+DzdUGK/3PYqY5r3BRAyynqIgdLL8+8kIa0jswPKXZO9WZwOu7Bm
O6qrsLjLihJLXVur6QR6QxqFLhS0iXrby4Oe7/EVawauhpU7RlPCf0iFuHvq6NiA
rG/4eeDWl1xS1asiKOW6AttkYxchsnF0+/NQPZOi+2XbQR5niPhSDSgawucwtuop
wwmmskcp6agQYaKa7zQc7uf8ObsgKwO/dyPIIUvUNTwnjOFzN48Zef0I0/LlfJqN
k31gyFQargH/T0vWecK0loRG7BDCL8616goGw8LP2TBdSsY9w5YOk0F2FSUmnLxM
EynwOgJ76bsK2dFfqKW4tUaYPngPQkiQQfdopLX7trajwk714QpWvXcmtrZqVOkv
KcV9pX1IfcH3i1JW14xOX16AR4An88JUU0HNXRk0sJ09qmi8PRfZCQdoosbaTYsy
4MTpiRtY8BgcyuDMxEZ2+fl0uglnQ8MlaAjXW6bnf4nMYcrQJt0ZTN8gcM0Q512B
9tdB7OyLlKDnpmMjcWsUYRmAL6fqQbJ7bE9aOAGM2x5rpM5EZeeC71TQtf+evslQ
t5WdPZ5+s/W/ueWhvRG24lA4CEX7ioldHCPXPxHwwJyR7Y0opnXBTtM6LWCtGd90
QXWktQg0Xk0SNtDRKXHGDHHbYcp3OphhztP/en+aaTW8cRQm2t+sTJtbI67bWzOn
3OMezkXiI/YNvc72IOumkTklx7y2OKtCXp34NN5D1UqMcZvLjA2qXmS5RjyD9+Wv
IEJV6AQssFT13HUOuGnK7sOSaTTjA4JwIfY98BHq0osEZJtg0m9tDWHVvE2ULTp+
U7YaiSajaPfFYkyH7EDb0G09d+/32iSRaGGIyN7/RDLoBBdZuQgW8e47gtHP0rV1
aQZeJAxh+2dIIAffqQ1sdbbR+fopdQ6gcAf6F0zGKX5F1GbLMtRqNX10+fmF6H67
xy1XzjC8fWJhghE1D/hKeNGDIeJnKf2pWsHGI8QBusB9g7RYtnLzZ6xBqoFkYCgg
kQR0tNGH0s77tUt/0z/JuNjs8cVxwCRjt/2VdL17ymVkxCS5B1HC5oUTauUhj4JK
n6GPm0WnV7pzegJYc9UrZSVzOKH+wclsEcLIp9/51aHqF7g5RXDMYhiPJpJeBiN/
OCOjxqRi6iGyw8O7tcJ90e9Hbw1C8rDswn3EDsnjxFViyvx/uyNOmFNibTm3v5l/
vP0AdkuUN4y7egbzrBJL+I9zWqpfjwmM0NdFr3Q0g1YHzkJehsHT8ybhHvJaUx4w
eEiikhxtCsPgaxSN3kgmnj6b53inG7c2OqfCC9tyjCA3ZxufRHy0stUz7/K+tJHy
vTubWAE3IxIRUIdjxs2wYAtbxWHgOGGsfU/LeCrbem/SqzEspXfSoZGmnfTv5kDy
jQlk4uBAv+Cg411W9dUvYYTptD+8JujwLpF4vF82J/tdOE79vfnVFPyuhpUcMM2k
dnTFucEb4yWjg1JiZFDs/nrEWdKVrrd8TaFNHsB6C9EWrtaxTl/2+xDf0IPD2z3U
/fTV2KtReVwWm6nGWwpGquHFWSn+6kK7fov8cmek9EJtK7Ts8HWSO6Z3EGVHV288
qa83SjwFB9V5OZh5SFmvZi0VFW4ZtThL0beCbLNXvT3nSRHKl9gXzmxpmHbvcz5X
rm1SrqiIx33QxoKNI0KBUkTfhG11jc3ufPTr3daaBAodZOSupgZOhsWAO/dCvVWC
GUwupHXvRkuFhUaHLqGS2G3LMIecZUd8OZuhPN3Q1FRY6Yr3yNaBQUtKLGfpYFcD
cwJj7su06YpdYbHGbI6yC1iQ+qO3YJAxWOxEJo4985jo2n9QNzjSlsIlOvAcCsuA
PMs3kuOWEFbx9O6IyWGkPNrR74zWamZxZEhYjMsUaisEot9V5LWC6BPnmV/AFo5O
EuQuZtH+TiKecXN/I/ssQAVmPPgO3IDMUl7aytdfwTKRzObc75bAhilVnpzpoiHD
wMHthXOPvmENJbttZkta9Rk7sTkAgvxQgaZ+HwhbZ+Vjy2HHKEwJkrzdwa39OThC
R/alBKOi3Kc+qVyKJFyycwD5hfN06aZAy7WLILICapUWtdeu5i81uQIBf9NQqwb5
aR3uiLJFiEBlr7bUAaNc2VmRTyW3TLHp0ST+AwMOIgdxCNk9CiQuLabI3VvqY3Yc
gGiLW0Mn1cwTIoLPLN+VsZgLJBLhIHAd6KZs/BZvMDDsV6td0Gcb8rTTggBGGPY8
xcsQUIBKiliDHY9r6meOKgrbMlCtd49MO0KRO2PLRojtWiu2t3ceKUjh2oCk3pf5
DbtEU/YzIKeei4Vw0HtCwwpA4sylAgOChy+j3KcLr7PgqFEZ1Nyh++IZVbM994Kp
5lxZtlCZp9jIhmtA9W6fWRGbJqzy0xuwHn1Owec4dhxBpSx0PkzT6nTeqdOAM2Eb
o7Ur8YeqFi43//hIgxU8pHdLM3FySmA2AzeLOmNLych1HWn5s/jRPbfSDd0lYAFR
XA7NDAyZsPhAu0ThAEvcdiBcMjNjUnkVzAsE5Gr3PCHWUeFhIXsjG3YW0nA5iH9g
R8Z+tBo+MAW02zdxZ8fQR5mzhj9VnJMpohN9w4zk3EIwE9hy5geX+SKlIGBdej+D
heX30y3v2+gvL7naFljf6h5uk9E24rPx6qFx/KHlpBM7yMsZYDWp17lttWKQq+LQ
hnUET9Uu7+hc0xHVTosEIA6kYOMc73vUyrI/8+myjZ37a/hsQaTsg2FUwGpKdVMh
369pEA+Q6F5maX3WP5M2s6kcJ2LTrX/j4OhhIz9PBgHvjOiOm8zfY9u4ZDVBAAja
2HnV+n6SJk4Ci4wz3GtLI2pesnNOnlxSJOM25W6T6KWvG9Giw7jGzWZ1JKqbShvM
oqEwRGOL3gnGcX+0BUetbwNIXufquiY6nYiS12loNhnv5PL5I74BTSPE5KnwvFuy
gVofzbzpR/BNZYB5lFAZD8OhJCiE9MWKAGo3WnaZaUzv3LItqHFhwiMGMW+zEm/V
4BAoKKvHBmzgwUUdpf/5Qn2H/HzK6HAVevIaLetqiU3Or1AEH3K9BfLKy5P1d/od
rvgu2uR+XJYeTf7ci7rkKPrC48sIUXw3YLTXtmy0XNkx65jEKbrZFCaCEEavW3/H
JpjcTEvvNBSMNLYmuwzW48e/vU0E1wlrzIHtsBnOwkdCbCb3gNpOLuirSxX+9KtS
NJxCuhcB8FcIb7P3JsLsmJVEg4SAjkxdrAGvU/MwxVGWF1oy8doweOkeodl4oej2
BG7vWPIjyAntiKheNVe8VDrJkHHMqb/wZ2u0yKmYeSTISpSgFFr3ixDEsURF9DEf
oJTct0JdgubJp3+tqeuT+3yyxKZlOgSEYskKgekq6roigu56FnsY/mGFucRKePzN
QruA8gLcqS3j7E+cy8fyrqsIH/WXwhSxoPIe32sTyq400kJ2dK7Oxpu0rNQT0HhN
qhmpWdTkcuZkpzcwUEiZ3amg7jJySmMIgCBAVlbSEOZXLfTfkTxmDngT9li/GB+2
Wyed3TIE7K+D10UH5wustcWMID/yf4nbOmsgbNwzSNN3tnqg7sFsFw1tUAVjo8XZ
gyYjV9fCaV5NlmoqBIilyrXUwAVtEK4NZYwrotB80ztiV74UHmll+NDikcqKP65P
DW4pA4dnE9oYU1yFgZKo4DDLxdy9X9cYFELoqaT+bMc6ZTeskKsIFJeWXZHsYshv
kTtzDNPENDFIij4gLPedYKps8iK+3sA/ho2FR79hmOz2+lfzA3g7t6m8eq7Ktb8O
VCx5CalLQCm34BQ6f5DXyAIyLGdsMYd02JSOHnqWc2Mhv9L/J97UGRM6LkjBB+Eq
GhErljqdEC7qdbYqACexCO0DKZfaJqmw1cQF3gjas0aKz9sT5RzDZuIwSf2fe7NU
a6pzPz0gmysAFA/UB6uNvouDp9vptObflp+yzH+D3qM3InuBQeNYYFiP1aDBcIL7
FyOCHrw0J/nLaJnKLTDW4bLg2zauLThFgzm2Gpi+wmH6l5NZ4G4FYyktQxLE8re7
g/np6oho8l2qCPLoi/zv45sdHp0nLLTgk+N7aaMe/MachY8CcpBuwKzxzXmKiCg4
t8KQ8ShD7iluQOk+o8j0EnTmAFF+4m7kPQO9yfmuwY7RxwV9pH3TGVrDgQ5hHrwl
ZM0yciav9zUrh3qWyWHOZhbvrnQGbgLi8qUu4JH+XJElb5vQibelj5xd27O+w/An
XsONXWHZgY3fH4bZHmf1524g4y7GUyIob6RDTViOiZb/CSmy1To2I+UtlhM3bdCM
DIQwsGzAq+jWJDqgFpIw823RH4zIA2x365A7IX6rfhP5ycmEjnNbfQu2REzNAOCo
Ylo2sad1auQ4Xfp92QxcpJ8rnkDApsR64qll/v8/5Yv+0F8dn9wgO2AIiuStINhO
s9KUx1zgOFMBohFSIazxlKJdF41IXLV9Jy9SUYlPb5UmyxZ+Zn2zsdlEek+OyxHp
IXgdTAdx2Q3+JsdgdI2Vd6WBgK9UmxpGCmgFZe6ptl0KXZdpNqR/g2j3P4vHFXR6
HF0NN/4LDUCoWDHKTI01cg7Oo9afezeW9nXxPaH9Ph+tTjEgzn3AGRLlYVdKryDd
bj5ndH64uIxcDGHqhMUzWhe/aXh7jcJTff++c6U6FCReBtN5CE+ALwx1J9/TVkLC
Sa4LeO0b9Y56AyZThw/f7MsWKRL30IQDHqnaHvoflkMB2nL7XDcpYPwgYQ+rB6le
IvXhfvhSjkOXv4HltN9yfTXKdg7QMRsUlbkevYnPopjKM6cd3GrX/IUgG11Qd+R4
ImsX1SEpqPv7ymJtfY2Mw5z2NnBHKOdPLKs1k/BgJ64PF8TRnxUKhinx9LAqan3w
SIIs5mNZz++A43B4Ao+NqXmhosCRioD1bRhV8aLQeiCZpsdGicT4GtMfkL68uCA2
aTIfzJCr30TClO1fB2VPa0zn0vRyDd78D5eyemoq46PYN8qmuOVKf7k7oRBhia0R
zmlcwUdIr5DJrnznpnBozEhrBBiK0nlGKWQA5BSQQHJQOkBXIFtKOZakHg06E6F0
S25FoSaFKvGmV9YbzuT/QARa6L5TC8iXfV2noTv82IfNDffM55H/cZZ7DOOWnse5
jCTQc1FOgLtJUyMICtFl6jdMlxNKyRx/OobS1bTJkU08E5cPcrmsSc4lelKBatbE
BW2czG87Pt74/0kzv4h/HhS7ImMHEAOS8fOmroUO/+hxJK0FKrIGfgoAH6xBRUU0
ctUXiLTR9zoj4b9ZjGohClgiFll5Xmbv805ysVTMeTpKtPBnyjL3pcaawAWicMFH
NL1WyufUoZ4MuWxZSZ816A5LtnBizpow4lFNPNlztC+ORNMLa9a+NBmJyY/i4d/9
J2UxhGKMs9LhGPwhPNshKN9tdvw0fv+6XEUdnmf4IWvFw+b3YLzuLVca6jp1jD6X
g6UfKeprucGjWo04AyhPVYDmdYIWYD3XIiOyt50WI/HpInP4H0mqacy2/Of1j3h0
yrfoLEZYrg2lFaV28kjF8qx+x/rERAFJyRcz07P/RQyfc02juoaJt1HiqAs5XmKV
deBzTzSoV1QjsRonG2UGkaQjmFYL9+UXc15/cpef0MJIG9AdCCnH/SPoM9fuLYxm
NtQ5POi6W4enmaRy8Htw+4oVCH7pjEg7BvRXzOPohPvsh9d8QKh8DksSXIFJIVrC
ozfzdl0UkNFWfFSZx0cdHupMI5Igd46Z+L5qRdfZ6lkCPtlc7VeGz92DBAe0G7EQ
uA4aPDgarifXb4GaRbHR39/MYTsBq9UPPcxtmsH5OD8d6XrZlna1bJxbVtuDTqlk
lcJHQvUxSsbpx6Q4uIKUdm/TJAk5Sfz5ehnXAjymBcjXgP4th3H1Z8H5Z5VZpoc7
o26cN5bT1L0yYee7Bb3MkJfC6KdKCgRH0jfqOW8qBoha6JBaZ51qjSfZCo5HNrP2
uJqeRRDuZZ+sF3RLclwBYTc1skxD/ctGwMDLNOhLCDYwMm6UexGPa2bKICnkiLw8
ayj391SpzusDQFzkoAOMjCMSOMG/gMKnwMerOQvCKOBphTm6/g6mgUUZG74gPtyf
wp0l1VC2xYYQWRRgWDH3rtJpCqNPatx3jCdjFr7O1/i3VZCuSYq+of8CZuMQ4dOb
D8pHDZx1aXjR91NUwqVoCL3vuObXGgTDA3I9LtMCLCrAR0o6/vhXflgdb/wd3aDv
00AM/E/39h8K0Q1++XNzZ8YasXwL82UJCSu5avmb7CXI/E5gOhzJB2QyBZ/2MC7A
ooq2uT3eGEKbWkCGxfo0Z8H/4bxI9LyM6jydPdf94IpNKlVYJP1tCr+m2tnibAmN
sSS14erJNmMZnWoPWPqeTLI0d5BeoAUDC5wSSrLJJ2sgjHKlYChvZDm0ueDf1cQd
ogz0jluNTAmGvy3PqYLGywa8tzQKpCLbFS/T6ILy9pqhMwfB8QwfRkXCxVwY/qel
INaNkfOyqd7TbR0Ddntcfz6vYgj38fkD9Acso+/IM5hcMOvWGPewM3V4j/YzkHDm
OeGx1F4OxJfUGE5H1knwIEW2dYNfbVJRi4cSf9tYGjIh9PuKK1pXos/T2Pw1yODJ
/4Ftl1oYModCyLUYfGb98ygs18XU2syM9/g/tq/GoY8Lg+xWBrKuxFT7LdgEc70d
HlO0S3LSsDFRCj/Wqi+syY8J4uIV7n+zp2/UKcei1Ke1kWLxnbZzrkLFyWx/W5en
CCoZ+7q/6G7+AD2R4c1IVFKTfD6zTueyGvHxQeXoYrHnWMXoNQBzPw2XsVtl77S1
Uz81AxajaGPx5TxV4szdhXpPu8PoefJaUs/pyso0Gd99wrMlSRMApY2Y2Ch+/HxZ
JDtSuHUVXJKO+hmux/qWBkFqui0y6CoPRLPbgSZIeJvsgp663zcJFMPou4u8kOJr
FEaxNmDXtzRrEKFeWWAkPhjn84KRI98l/mxnSlOYvcL+eVb7ES9hWP234AVI6VFW
YmvKcmpWc8VxIuGuqhz1WasuRSN4niCc3jnvBARsDQ8AcNbHjAiptozp2Ob8GMNb
q32ubt9qOIbNL9D1vtcWr+aO+Qb7Gvnrpgac7GDQ0EDZrKLImwT7k6rpIHZCjNZv
SNnU8Ns8S/YAbKmIbITyqJ5NX3Nx/KfkhTcTfsbJYIcBUPhh7O56mtQhVXji7flj
bXNnMkKotGQlt/j6HsvzFIkP3iW/Qply9p6y4NzXpTho6Tk10V1b8xecDhOgde7b
zczemu5zM8nAiAITIO1LtwonWuwcvfyxZKfor9MaMXUEV7d5a/FFfRm85acEXJw8
gTKW2qc/AkBIpomFKm+m4+gpqRzZSTDgqTixoroouEl9b5I44YczgEqoFGHxMBPw
fguP8kPt6QFI8/qmpxFPDBQkYqTxt8xrhO0jwb2QSmzeJjQxV9of30Q7s1CgfPEj
KxWBcC+8LDEUOedmczWz1DoNk1qUIPnJz2I9h6q4sj1zrdwDriNDsQkfPjZlroiI
QvkrrtaRoMDideDE9ACBqHneij3bsLxQDclTt+CJZOhuaeY1sBmvSbwsfUmEbkkS
DpVI5w93U4Vm2T19NbF9ZZ0FZXq/et2VXk8DXxa+LsP2/dJMerFYYvWH7mZqaCjn
+8ordIuExlpnno5hFP8M3MN2DgL+ADnMfxYn7+RFwF1IAZVnLGulJXF203elNUE/
EFPtfft/iWmVoQLChUWgeJXgU8Z266+Ey5/uasKu1lic6KAcYyUW7CAtbjoqNMLu
rQbrnSnNbUdCmX6ZkksIGyJY1bW6qnSSW1pcf01et0ZHH4sNPeQ3MHkVsjrTQW31
uOVoGv9Frmdt6sw2GDlL3dKCWg+Tw9d+lJhOQLe4LtkcAbK/qXe3iFT1y7EfkVDN
widP47pkdAIyvd57RqcujbZo8UFlqhsHD0d//WVUbS1co2BWBW9Yj+OQd362Z/hL
31dpa8VPiuXqqFbryHbdbebzD9NPr6SpVTYTyelp4W1LJTEHRLL/r/uHKl4Opu9j
AJ+AanO3r58TSMOSJMq8HbVaZZJS89+5vuoMz9CcOgt5i2qrwiDKGfI3LkwZUlDP
4uClStT/8g7xBtCBtzOZ7/ExHeho2PGy6uRlPx9OgkeX8tzUOtAoTLKzqapI4/OI
+Zp9BkN7bzEpQGNUgXMWxG8mbMlvy4Ajy5xtCP4lDbB9cULhdHXBeASsPm8HqXJt
2c6WhVdoFw+hPyCMuKGQCcItWfHKRcebhZe1y2URXOnjyZ2R9xLUjDJfRRYtnCUh
pHjlG1i1AIB/DCKHQEtWryEATJEgXwbNJAdDCbX6RP7T6G1QtbwJCzW4Ytk+ojQm
lqacoLvrmAcYp5JEKiLye2fW5z/mmHYeDL2HASmwblMqIw9oQGlqoogh1eQq7Jwd
mCBbhBD12rr2ceO2LWwop478OsJ1rAW9k/jmXsGCByQGtvE8jg58iMyjARniNvcr
8bE+tiI4yAvWZ4WzOFBNbfyMyrqYmfdOllTttuNYztBHcecVLLo2gnEasBEy9oA/
X4foZGEES5wLutRWcr9/WaP8ae5RRkHlFtTkKmVIg1nV4sYjI88MrjB61LY+1Vp5
ykmTuwX8ORj+YTSjSWseQQu2Y3w8eBDm6sF+qzkUkX6qKUL/1Qo2YKIiSmFmAE8b
+x4MakneJcrQjJQhrcjVgjStbKo5VcekmS6pNced0h9LnRXhgjupwb4wLfFDwdiP
jOGUBqL9zH73e9Ku7Bk0LKptXzz/AKjsy36j7BCDkfuBi6BrqSL8jtwtE0MtKYRS
e9FJ8MxWgPCLIruKGRBLl17QNLDajQDhxUF2/ezK/QJqRHUdHq8Su8b0hKDtALcK
ZUHASXtVoc7x3xG7gsMWO2NDqFhw3Far1PE+jB/UdF9wvIGrOlp+M0S4h//x+gkw
eNCIMCVLpoqiRZP/rw1tt/le0iEPIkHUBBcygcWNxv2RPNGhTOLa8dV864CwyJJy
VI+YYdrHuC/q5CR0r5Pd6d2zfNZdJHPLWolpzlhuYfZMcv5izJJ5scvJG6Ah84VU
q9ey4T8wC10v3vRpvvOnxKLOCqADeLfv8dSnct28iON+knYw/VOg3OhpI2ac/Drk
4QED89kpb3xF1jyRZ2oSP/YETZHmaG9vVrzgpKtTVtQhtX78ViE9Cy8gWnxzKD3a
lH8+2ea3a58p5pl/zYXOiS4VdXBDieTRdtFGuUr6LEmf6ajFQ8bzfkxImbsHiLFB
bkBHIj8YHEWwwobDjC/FD1lObQ4fbD/OZ2u9y0BZ9Mlf7LaaHrDZpydWhY0eYtfl
Jo4pcIvMr+TyP0R/vRIRZGXYYtqdnj/tTNDzISCCamrWHzVCc2RFnXYbXC8G9SsG
gqXrsqlV4l1d1PshwE7BMEKLqv2IGZn3Gr+2ExCl6vIhYqb/SQ1RXL4oHig/+XfB
KTxYCyd8Tw0uBnwRV4IDBh6alpaW3BIFlTuX3H6HZHUnfzoyOR54AB3r3fuJ+Zsy
j25IRcK/qmfD79bohwVfCemeJp14Zup9i6whhAyI4XWQZaHiKZfxjYA10vrAQ7G3
UGzGYIg0pZgmKApT/Ev4on3pnZCGdAiFxlseL+eJvtegr/qn3o7morkMVrB7kgeN
ZZtoZ9SZbCztjtgmqqzpX88qmGXwzRTWZkDaZxKnY8P4w9ZJyfSok1iz9+aKB8aI
Q7KooeRYvir1FQFQn1S03kZuv0E3SoLMZQrx9UTBvyUtbcrSp+BGfwcmtRvBjQ3e
pPpjJHrsHbw+am7RCgzO8Ya2M767odcnE3gMT2XT3Lv9Sit4nx5wEMvRKuRW2T1S
+2Ig0Pl8xetf1JslPhZZZLD09dawSypCeLnzb7MezX0NmFCyPnRItjCfoSMb2yF6
dXYWIUU27Vs+2dpKBtpdHX9kWa9IbhusB+KScyubfyUMPBMBiv5PJq8Nfjpk9Fon
37Gh6co8FkWR1Oc3b2e5JLqWuHq2lyMUhsnJ5z64PrItUSNh0LFGQsWW2B4ffKCz
gdqzrXhFHlXr7Bbqkoy6BcZffP0GyKDr2EScZQM+ym9NgZ4VuN67M+K0t05m8dOI
4ul7I1XT79GgGgoeUJcDbNYLFxoCp6Qqr4wyu07WpEDiEBoil3K75Eim7yGwzEBj
xiLLihsJIVl/jg5X2+3o7jP5JuVbRlbzSzhpMOXL9G5VFvLfXBrhZ+declqBWeX7
HAvOX/FokTW7+cPsKcCR8ubAVSWygHncXTF+Pnqrax0pg7KCsbsp2GsgiGI42ysj
jh4WIgkkg9PkaVOeXUKFVE3kq7SFrMEM/rRlm9aIU1JnpMPYJahDFWrMIq67wukJ
c1o1szMsfVwch0u3Zvr67WMScL2Z7HTklVD270mA4IcDq1iQY+5aWi5iSmyFeYji
UFYL3WKkJvEdM0P0elHlfKSI8tyEpBvAInigt2EMY/yGg4TAn1Ow8B2EqwGnO67l
dlq+gfPcj27xId0i8hbZL9X+jsS8L44muTsaTbRIz1kUDHFtmVkprfJNPaktAqM/
HLvHwZNssrt2CKrgySK+JVmsrP2y76jM6x+cW7nppWbdtNFm+z7pIH4IH69lYdd6
qsEfjj6yyBko6vPuVDyCV7s+37A7YN9oSkuAYJxStBi7Zt9EBK6e/kHiyVSVCJ6l
oNrTpH1g1390KlO2Jk2fL1/ymZawY6JtwhtLA+MYR15FnibCC9z0AfWuGtxTZWKP
ss7sgHflz4hnvXiuEvWrKuP2aMVLxosP1lf7zYSwRzQevadCXxw0eeEb+vb8EVPL
AQxekKwXs5Ml2poN8vX0TI8ToEYhugS/iyEx8+xPIVWP8EYzf3IrMQFhqhzHiye1
gs7BpwbYnehCgXAkPbam0GTtSu2M1FTdCocs/L0mBQ5vzNuGd5QRi714XiZTRtNs
C+AiRp2u/EHW/odUuXOqEMXY/nm9tvqtRKO4hNe1qH9cfj2Xow+dUDqddNeZlYx0
Xukj/h7s4jF7p3M0lOdLZMxB9Lt3kpgh9IHFuKijzYePTmXMsg1Jyp/nEogEX1rT
9jw7jBSn3MPdKdeG3lcA9fSrdqAMDEQBEYUFXHSCKQhq2820VRWd+hJfiEhCHlVM
/e14pceEIqVhtwQJq1UDXL3Rpt5ld9VPuEJcJSsxPnyaleZt9hqVVnkCq4I+vDB2
+sqLv0oZzLsEZQjIIuI5VrJP/kn1CcTK98yCJwkkYoETOrU+3XY7Lw1TIfwhBIBH
7ueyoU4XnuaxmqR8DX1Ee69YiJ8BpVcsdJoGewkB7sw/WtJu516DM2ksV/1RBf1A
mPKUewAkR3hxOT6ii1sHUvvKekhqDi3nuHy8oxF9GwprZoyshCoFWsr7tY8/cdJI
7e2tsCBLCD8Z009k7llgZrWMOUOMLlYIqrwsBGOcfkkM0n4RMqWrK77pSu0svgCm
dN2CIM+ZousW+GdHhq8cUzsCJTrtZtV1uJzyd+YAeLDORKbbhPVGDp3NxU3s2K3j
8DjMCOsHqfu+5CLFflM1TCneBmybZ4c6k2OLlThDEkbf0c7XEWnJWM+iTBkr66Uw
Rm7k7f09TLHeLCiiqMSQGdKg6x2VqxtceSTcSqvsE+yGS7iG8S1rO+qxGvm1qjgB
l5BUAqf0uWROSriHI28aK1dJXY2vdhvUHJuYiqeEYthXz0XA97pJFbGSQmISCFr4
YbYZ2aLZDJENI7LpyPBDsrsY02x5DFdJQmRt7Jo+OPw7NG0iyx1oZGgiKDs+z4vk
noRcYiPkYF2qKzsQx+nrnNojwRLd1nRGQh0DyGJcncP1MACnWCkbJerH2vDzDxWu
OG/fT7YbX9cNCRgjxYBjcV7e+aqSJLJ963CQDSoqRkbzyMcvRhtl7I7yfnLLaPDA
NmZPGLHz/zHnHyYHr1rzeD82/gznD7XP0Jd4h1r0lurzvdS4V4lqBS+k9fTbEP09
AKSo3IFMnStG1qmKAaMzzM8sL9zvIqdeoEtO673+Hci5/XETuuOH0ntUS8oJIS9U
Y6EgfiPstcDfFTA3vst+Cx5s/kiCZZq605ydQlZhLgLx5cA/7dkcPK1sYB2yJaPE
5ru8WaFeC+6Ty5E71mpNFQHEMDuz21jK9nkP7DPt8Tm48ZFrh3K4t1oQXEgG2WrQ
TD8MNTRneQ4dtc7aCpmSr8hXNHhRLG/MTHbiwQjT++NELiI9OLUlQTGBXlYFNfAQ
ocygOTKnL02gU0peSnPL0+FoGpX5/a7U+cCJwMiFvdzNspKK7vszWJ8hxbmMTTYt
f0HmkKYc7+Kf1EIWIEXRsC+QWfBramL6WpmdQZOD1IM7Hr+7SzikDSvFxWIURDbp
oMzsz3LHnlJ54FS/U96ZKBIefxFfAKqYmYWp1bAJh4R4EGtAJ7cA2//lsKBsP7Om
M7We+Hms6TQ7PbwA3Iln8QaM60bPrcqZ+j3bAy96XkK6sApkEJ3mPRquga7+LiKQ
qapbUbktnORztR/Vse0nLrDueGCp6iJKApZ7u78KTr6+fc534rXXxqyRrEgKcdOT
qTLxPE9j3ICL0Q4oMfgeje665vKxB9M77hVGFo0zJ4p352LHQtAG2utuGXKz7yuD
WxvNUrCkQUl0m8ZHsAeKxXXxAf2R9UB/LG2o1LUdK0ZjK6KQawDYozcb+DBJqSF6
lIF6SeARtZIO8Q1oEdbDdC3bEmdobByMj+2WMv1Nr5eEROTQpVaboS4SoOYLbYb1
cCboosC8BFu4WpZSMDCX+mO+35hHOD6cW0mx83RLOYoD4JvickMEaZwq6A6pj2Rs
p/A4LJi/D6YcBPiHl7y6UDSzloM5pzPRjzDEpBzhMaRrzBDJ18k9hABNpeVxfig6
ftsfLOwJj0h5HyapZhEjOwE970qLRbtxhQpHM/OO1CvsPEa7dp+yRTXxSs/2Evpw
Yw2U7+646l5GpWG0u9Undmz3H0hwiRsPd1M+Ey/uekKdlha0Euy2f6s6w4lnepEy
Icc0tOJl0EXc5s/6Pw9pxUolPoJQabM6q1sR27oakYfdADW2qYZRgjuwqob+cMzb
b6iyHrxuvMQ2JBNdEGImlty+giE/urxJm3pPYOax0JUBc0sPaZVxLJYRlDUKWr4A
vN7d9gjoDFZaGttVwmxGuw60CveBrs4UnJ7mv8W6Rfle4n0B+9dgw29KXjaYTJYo
WHZCMh4FvMdeUUAjTJeH7G4sFkl3bXJkue2OTgFJp/aH5Ser/1CBNIxMitUJ4M5h
XJpOpKBSBdoFRIcSw89ZnvIGA1kUl4ECycH37GFqbSISJ29SbLU+Sq1exFxLvrBg
WK5//qFD2tiHgiXhgLM+RyXzULVESOe6RGeng0XtGqsCJAlpnZJc71iorCZZhuaL
6F5ElfVtGFeJC9Wjd7rTPcJVYwZ98lf5Nc/1ezs0fxfC96/xXwtTvBEfxQ2IdqCA
Fzte9jntTyiAUIP9nx+uSD4NTiKo7Sl3OngLnp1eqTog6uFZgYBc7szlr0udsPO1
C4/YW2+nNkdCmHGrZ/o/48dIjEUS97M/htKeZcwxNvBt0f8udAlKGL/QgqmyCq5u
Ur53ItKAtchA6IXQT60M2Y98u6wx9VnzEzAKaNG2NdE8LlHWMDKVA0b69eZYnqoP
B9HyuoqBogIlXwTjWdlwz5ogsQdGDmnh6aCr4Tzf3KDwKVQ5UU+/6ZuPwa41MCL4
Zz9Fbc0Y9hC43xbSI5cRdCzEIv17IN2ACiwGny6bENTaqmD9FPjyH2MCy6On/Kvs
BHAYmXdL/8ws9xIDwogtjkSxoWHUaPeJlUMp6Ts+Cz2VinnKnCObamJojb9KCqYC
QnTw61wM57z68yo+0GNC6ExVvMgo9IQ1pyEs9ew/UCHbcNsx9TvG0UE6WaxwiS1O
kFfekCcHKGXCtU6CqqWy55xEbeLcyDdAgqWShnTM4w3/3ejdp6n9/JXZmQ6LuEQ/
k3a7sIljulte3ioMTb+f2q1ngW/85ZFyV8dE1brc/GXuK3xFH6AyA4qFVE35UsBY
c+6y+DGDMjPKl6cBgbStcwK8Ws2hkzlDy/RJ7JRP65tLleVwa3q6m9kZpc3jFcme
d9cHnjUpiZXK/fYhJ92lz5Z+0QVlXauO+m0XLOi9uCrOSca965bDm8pgwl40Wnko
kJd3rKznqpUOB1tODvfwuUoC1CqZSjryzC/wMqmMGF1964UL93cAsv87lCXlF9fW
c3Fz4MvWJt9Jo/LisjLBoG87dxRxd4LkKYkZrHaYZrV+5X2nhw/QOu24HvuNOdmw
kN/bfY3gsWr9SlAo3GWkeL9R0wlahBvVvTBiMlJlyR2kGVQBCY8w6AbaxVteawJL
nwBobZG2fSP5eBf8sSQZTEjgSp305ln0sy0RMVxr5zjm365gG8KgSemkwH/MLQeK
jzkXV5/sp/ZOGiRKxQpWmaCedMCICSgOIDnbskQIM7Yyn/WPXEn9uzGsOBE4+Jy4
mYnW1TqJ0YTUA6tRUy/M1VDA+lIiBMugiFxx3QqxeXoBqfwzrOttQ6wh5tOEBLC+
zVZwvkAEVZtKIlVQE7zjbfGA/gtmMeXB7+8X87xlRGDDWFagXbWliIIcPlu0rzSb
aCzWC3oW2FZgnMwoUM5whTLhzGuMWyv0QjxSlK7LDnbYm8arcz7AQ5MXcZlQdqUE
BKKeMqbcNxt/Ci0IdirqUvfYnWgiCM/G5XD9yw+rYHtY+HjtDWPbaV04bSRSmqlL
DHPBLS5kmXHkehNggdD2fFerbJ++u9Ikp/x4ofBMSgHxb2VWJTm/0XAcQ7WRy5BM
pX8lr4EcEvkGJC4VgYvIFgz1/y7zYWBpAlXBuFoSBMID3oZAm7M5mPVBaP9ADOQP
JftocJYFg1fa9LpowpiGpx69UKr7IrOuZsS+k5CocJpuvvuFIgnHjur3vIDPR2cL
GnukQ9Uw7f05/t+RnigTqty1wI+em1d93frT88tpKdHwN0dne6QQQiCKRFSGExyF
IzTvOqczRTUmuvOxhe1RjuHVi7M8PwEjC7m6jQpX5k0gbvXS4XZ/QTrSeAEevrSE
6qGbhSEpf/y+KyuIvxJUSCA6sYwvvGBwV4WR7CS+BiRmhXAXug+zWlbQqdCPD27Z
gKk7YtCSbKd84e+S05RXZcQ57pti7tFnrON70eaLxQ3re5fudBQIVv9jm8OybVtp
Wdplxh0xPf+Ph7nxzXbT6627ep1XCzwRWgXpjhy4LygBKoqYPdYH3izCIJ8ISU7Y
eR4uFdVrQomWf4Zts8hiq70qgYr/YjBBqbNvToWBXGP/kwVcqG8yoUn91Umzp461
ka0LX55y9rlhPJKUQ2/iI8EWsPD1b4el3HkE7n4x+KsRWUJzqgit1hqjbxx4gMpc
XjJZ8Xr/uE+JuLlb6jH23Aw96+/fMP063Pcrl2Aa04wCUpwp3PSOHrqMKStebSsM
42vyFmx05gN2GqZD+vO3M228YMd9wVo974LQFWm2zrHxJ/QJWWRrGTUVSe4K6vTc
Vi0s9IJVhATrf18qWF8g0h5Cx6qVUlCE00NQkO8x+wTmfpxUOKuIQr/AJhg45muV
lDgIiHJ8al1vyixn7K0VZjG49bGA4iz99Ev7PKUdnnss1JEFi1elXFaJS6Ej2G5q
SzXZdVIA74hlWjS8H41FXFSVwQ6GbQkZFhXBQRnAXTbZqaom2E4/B2ps64Lno5ZV
wYJZCf4I/5ZXRHUEkC57+klt1ApNKri3fbTJD9Lf8SHvhbigc53nLK54nNyeyLdH
81niMIy9XemHQgParzNwAtf3UbU2NmTF1W9s4HvH9E/+e/DWMTWpm3dJ4gi/Z6cK
f/Nl1dIlfd7BpRCwmY5f+TU1tg1VwlxlH3sNnUGgv/z/qiltFe2pnp6wcZ7m0U/a
YNhszLNzT4yyku+Ynybee1g7OGrc9oNhCAdqdg3UXqumG9mHJcMY7ADlpLNl422L
aeHxTn9k4D1R/m5k9AnCA9UH+f3/OhmeOtsVCgdofFJ+WtzJydAhXB0mDkcpwAnX
0MJyMLALMb76eAZROqVmg9yR6yHb+I9E/czsk+GVr4XEuoLdd3+mTo4/D8G1Bqed
R5KFmySoMdRY6kHqU8V17tNI+akV00asIvHK7Crjc7vuxUIqqHq/rwPHBRW3xrom
rK5a3DdtDA8toFzB2GzC13ziyS6PtVneQSJZ4HwMMx3aM6BuU9z3V1c8TK/8Kd99
NV0ay+6Dwvq3DddsO2jcE+cnHR7hEZ6TUBy28Yp50axs/MENTh+4yK6Oecnl/pnT
WW+aFpVA9O120I3jio43dXixn47V4cI+BlKuX0gLEn6cu49QzyofGW9YHF5jSEOT
6/NyzAdanZInD9DEq+ehQc2TFGhncwvMuxxKKpqAh8NpPHDnVIjjR83seqxDprhc
8jA90514ZcduDTH1vr4UcI/mqHXIQ4YAfbKLMPjs2ix3Y3SiM3m/A7P8tLyGPZpc
iA0rhxQZqXgUW4pdjjXDqPJE2TNlk6M8PlfwDhQeqz1s7V3spBxf9uN/rpR69GUC
p2FdYbfiE4rjYVBLYFBCejXKxL9643RygbLuEo+N0UAjA1ji2L/a5qZaud91/mE0
UzH0NAhlAqIFiISFSHy1f/mRBrY6sfFMeguTamHs776cbaZp9EKorbgKxkm+Z3gw
1W06qAsZHe0PTHVEhW8VNVulTBctAM7PtCMR1EUFtlxq8rAJq3SSPaoo6hUfe6NX
9lErJVlaxMnIa+BtShPLIcdbazgt+hskhNXx74DqPSRuckfKUDGveKrzpIGXOpwS
0/SaZfsX84e8eBnuQDNQtaIq6ZSgo6wA5YddZCce6uKIzva3wCP6KvjQ7YS4kZY9
l54m7Tbxk1H/l3G5rjeRD4on1dDQD8YSx6+TlUTzdS2VTUpvc3tM/3FJmf7AxOFf
GBRrAsD9opTaMOM9Qnj6Mq1A3tRkYlACiIrZh/rGm4hivxC2YwJbicw0O5PIi2cE
MDVOznosvFEqFUzF1nQ+bufSquK9dOz2N3is+0toWguJhTDSHo8hUOuvvbtIztAw
8W7O2ImoUVM+fN49tN/o1Vj22YbBc9E1FOQFgNWd9Qasz7yj0IwEbE9GWSCIMnRL
oXz5MahNscrUzK/n3gLqs4fjlMiVED+ETtoHpyyapiiITlFIb4jDABd7kXeF9Say
w8oxZQhcHbkq4lZuv5IcpAKQqWSV498M792NIJahwaa98TkhzXEnaQNAw9/dEspp
iucTUcFubDhHWQb9UyXYWLEZdfYSQ6pDkxnSDJGrmuKfgyFtJxwk4+k1iO9Y61f1
oEBrnWQBlZdgCmE7OwdIxF0T9eJzN1xzNNJ1fMm+R4ACDq2xtwoZYVVhY3Wj8hMh
WmpMqqhRSXy9MN3WZ+8uh2rK18nULqbPU7Re2gEs4dKiPi5xYLVf09MF90gWOIj4
OgHOIFKqyVOIc3Mz9ipGq3V2aHV1qnNCbUVSpsUQ5mYGMrB4niM+GKUtAVt7xhv2
CdWl9PopShRvxA7dKJ9WrbjE0Kms03tm/xsLK7jVxK/OOJkwXAV5zWXIAXnlgkh/
Nv32t5lasaFhYatbNKnK3zvtACIaPXQXibKFwOm+aeOTA/2Eai8GN1Ktmr2W8aLM
qORUqTk7d4aUuZ7GCfsCN0KvmhM9ZDyFVXxvbwYY3wLqGIxkTbyRvWYOPtPKa3tR
uriNIGgWs/lzMzXBg1S1A3dGmhGbnyRY25zQvSggbDguR6Fe4vZc7gxDU3QZPh1u
7UlZxA+nWQ7Cd1jv7Mh84qBfyG1BqKPKEffKik4Badw962uA8YC151mZwdUIlDbB
XcFvYr3uQ8Zl77GC+wN52NiXEx17i1qMJLObwSsaq3GC2lEt6riygH850onkaMIh
YfXCXt8dt5jWb91lwif8FhXPOC1QtdmJcLv7RfLQJR010VtMpPq4wu3dtfLIkT8b
XWrVRW0P75icf9DQEocfwgGXNAkxmgobHh2lp40rVz69mZX0LrE7fPVHWWgwA5Eo
ybvyviAAbtaDBAB0PFHL1eC1hJORy4QCZCSR/CYQD5fOl/xKc4WVKd9MpMRBjt6V
JmL162hhWXxzzbS5tvQ2g/jRxLWBFkAoQIrCwM61cFnjXsl83gEUHq6QWbCJVaJc
Y4j3ZrUFJCqyYZ5XIjIPPoaDCjNNNwhcMZenv+ccG33b7AL+pEssMWuv6qtiAt9Q
pQH7rFHTJAu3IVxnep8lBZIqtGaTXb5cbzXudpbkp75upl70itwifFDOPC+i08L9
J+ehNx1IFS6hdhl5MyUiw4grgmgaJ5RH8Az5IjNrpPmwZfnY/XvUmalD2EExX+Ra
W/XmzksgIuK9Q+vS7on9auHkNdz/uCSgYoc6P8N1x31vBSGU1DgrpoYV/uFRfquw
Ftr79/ho+MiNNrQgUYPk8cXt+YHWJhtdKRK5g1z0tTq1sVJJOrPPvDXUkopE8Tom
kd2j04OEgAyjPpm5LkZIKeCcPb64PwPvJCPHMKf/0C+bjoC0LDFt3qIF6kuZdmT1
HyKngx5cwXVK97wkC1drrbI4qtKE85pNyoabdKraf9uDSbjRBT18Fdp4387NzKqs
8qMSc82SsBX+0G3jApk3itC/bRaqMeTx3JTMTHMiu9FyQQ0Mp2yueDqlNTRua7JS
ajdhrssMSRpuKvhdHEZRcfN6x1sW8zqkHOH4SG7jB8hdAWO4cDG2s+6db3Sgt+lD
1sQ/j2qS/pV98jm1t46p/OLTsT5cv49uSCBVZz9PhzNuiFLSDYlrKpxWlrYe4fkg
hGkKSrC+6e2GwWzlWnYH6zN2dKaNV4jaAtZuJee/0gnaEfDlsRwLP8pHAOmHK025
ScXivF2cjS9crcgSG10Xopem/l9zvFstetjcnzxUjojNDg1P8LHHDWd3TEDyUHkm
/ZolBle89YKqS009h3ELM7XH4Zeq400LbHHiRnGVuBRXUy94h7yiKqBUxAGWZ+Q1
yMPFYEbofGjP9pYBmMJ574Ev1ETMGcoDDnQKm9/AeYJ3Uf8Xgda3lSRqq/whALmY
OhVMZARMwc3JyCXXT0qY3oMF4S/CH+8Ycfixg06ZVfUoDXEzJ5BmUrAyCk9U7TFG
48JGZ5ROEo7VEfRfI5V/4cNmRqiOjan0i75j3Ry+FhnfgrL+oFVZsaK2/o9XY+vt
5hCIEp21qzSWeaxFGsBtURY621EXs6Qd/zYbfq9/7htRZovae5EGK4eTqqM4eG+t
RlWHVUNwcTcj4WnRIrAedZGpADyOSeMThJUeEcaNxTIkFN7RE9FRutiDvcwhTZW2
RlDxyDi4VnUdPG74SMHA/fmkhD6NNa3ObPXggLilAZbPnldwqg8cOs6Q/NV4vTSB
CkULssrGGBFYse5BDSRh4FC5wkJ9a6/08V8CHlrTLc6N96q6QyoyTWyj1SkSGN7+
8mVzZSiUku7RrOBe6VcSLMTl+CLsKZF8DYAT8Xz6jWwIF8FqcwmkANMWI0C5+axJ
weFbluzvV0nWSrJicnziwhEGRLj+5XpLIVRh2QiBUXCUCZtMJ/V4qArDBschbjIT
VzpNReietcvt+Fo66u6MF1Rv30g92WCgHRtcEM4GciYkbTg0a4jfMiqjoNrY2/dW
a/CbFCb9enR+NAyWvY8qRh8wGvPKdkjMdQMDs7HBcpedTFCLKFeBhC7xpaBKwEvz
i2BzCnwiktjfs+N0+wkABxty47/S1lTajnflu7C0Vz5TjDH2W+Q+t/BNjsfGGlW2
VU4B/hTjoBniIhGhxvS6I7+cq0P4Id3Tz8TpE7uqfBflZlcs3z1Yz+/rgv0g+39k
0ZTFZMJsSOb0vEP3Z1UQn5horhp9DB2Rj9U2dZt35u1NeVoDBW1gLC3Ydh3nbnVb
SsCKRmcOisI2xQutjKKn8oyHkJPQqT82QlAM96Gk1AW8XGJ6lU56vVR8t193sY3a
+FljHelszWnF15X4Zj+YR9lDPBR3u2XyXD+uYtJ9u/GYSk67NKhP+s5wS4TZlOJQ
mH9fN0OKS7tqlT2YWOSHMoj2XsIwgxwsNM8sUokTfYNoi99siiCXAGRfygH3Q8lZ
BT6pCqOih4X47KdORnihoGRljhOw8+X1/ONKfiSUncmk/vuRsmEIQqw+T4fKDbOy
eWbeZshEjObi521BFfLdeyLN7iKd/8wefkl9aPg1uoLwdSug4U3J8SL+YVu9wkTK
mVpFEEvZeIK2OFzXaHyeT9420KuCb/sFugbRKeauDZA7NtAtn1vWiuQLBHDOMS36
6lcNf+lLshPdNbj38C0wr8zgZmtMy/fevgWFDK4cPK8kWBZDFOJm69B7ukheqKVr
4xs8ecQsGjKAwDSK9TnjXJkI0TBxU2FGqRCMJLl/QgQyCiJr++eyZzQDAIFiVHDd
oxEqrO6PL2YtFQE0D0AluLt8tKL9oWZK1A+TeHt/71Bsv4DTFjSKS3KHTidBl/tD
Ed63kY7t1EwYhJde1iOr/2DGQzyE77YwwE119LVhs8vQFsqes8QauZhduRQTwLlN
LQMjP2EriNknsi+7sCaAWz0EvNn9j+a8PmoVHxZKoPhhVFytfi3u7P8vU1SwqjVX
+dJLhYRynATjwiI4CfW7Z8dLt1OL3F+9tugCpwqiQpMMHL8ZxLFoO/JvJV5ersaF
erTbdu/FORgqZk5l578plNRY9qy/VGjqsgi1ux6hz29RQ2TeXiY3ySUgLpEeN80P
/xz1soCz6LQhbsy1L5afVcbFBVOV0LKI144pwSHlygTy+Vns9kCIDTnDBiL/eC80
Q+uDL3oP2zpP9zv+/+yiCY9j39ttQG0L1SUbTIyz0CopCKallfdgyTa+/8Zq6kyE
rD+N/87TpGD7CF7Y+9wyqsBQRWuiGyt+r1IP68ovY8ae2O0321hY4E0LPQU4HdEk
R82P57g5YuyaunxfqK8geCmfkHoOQVNcx20ybrobTkwHiQOgQypyD5aw1mDdB9KY
ap43Z9pb94ZDvVsUN33Aw1BWqZFjehOnAf0h80JAl84MfSZIsZRaBfaAKfVcj3z4
Mi3koYSfPo/JD5HvLw0Ug0mMwIvCdEZLDDVj3XCRKVgfBO8hCIfVdkIv5hi22lyX
HV2uwPxY8leyTg9g9TXy2RuJ3Crd3fIi2SPHUMfO9PeyNT8KidKLwUsn6ccReZu9
4qftCzhMLpxFsKGsCV3OwGJ9GiSzv+epGIldAz9RCFihTW9R6YTWxhU82OKA681V
7IhCZfDMTusmZvFImi1ulA4ZUVhrAVjOBQSCs/eYIiwuVS/ZD6gsPAWQA0ePpE0n
vTA51g9oFt7SMOSxta5XRsd/FGAm8l0jF+GZnIKXhxwduLn16L1DRiSwUZttqqm8
744tCIJYD+LazCNmI1AYF0ZZRwoRuPFyyOMtyN9+gVu525HIhvu01AGdo+eTR0af
ZVjD2SJ9acYLaTBRkgjaE+ufwKDp2tZhrd6opFF5ea3PDs4lRCSEqAgKEEsH4ZV7
h7S9wUi+uRfyySbUZh6ZHgxDOUkFXv80+317J7T8OjVfCqTz8xXYU6Wg+eMj0N+C
buc11tksBScvpjfVqUlUE5135hX24zHZImeBEsefjSQwy8erhFtKbW8CzXWN3yG9
yMU7fKMT6XH5yx9UDko5IXNDldJKIYRfJBCVdD7NzklOd+gjhe9UBl4Page03I4H
MGdtb/ctw95uawg+EoRYmgzy4omvSGygVvAn+B8wjCWe+az+Sj1KtNuCMGWk+qdo
oW2m6voG63+WbX4Nc6Be1HREjbV/SCqQBFGCWh25AMvDpkch8anebHihHwYwtmjC
HzyBOoaPyU8f6HuYIZDA0siB7qsSGlzypk5+Hh+n3bq4jaSU2+n22ucfViEuJb6W
OTMgUlb0fCawfZRVvQngMR/7gvqo4UHXqdnxuD3ZJB+yemfGgeQqsvc7SrVpvLPQ
LBzrsx8jqBHGExOGkT+Epg25+66GK+4Z7kGgN674YMUnovtXDJr5V4UABgamvXHg
txuMJ0swWiaredSRwLsDm4pS0orJGfm8sWRK0OcvCYa/nPFqlJMUfAtWMIgUdbip
dIH7w/XP1vKQjSFkmpjtvPJIbBhV9wgm6RNlfD+ReLW5sfyw+G9t/JeOtS8dfx2Z
JwtZ+MFZOk9aPCbjbYK5ZcM1nZ76r1qruSo3L0pJU9y0m96YuXwKQat7auQVJ+hy
gZCeXEbPOaazoKPyCnoufbH9bXEsJrN3WgUFUU61F1EVu8YXcr5TmU8vJZH1Qo5N
pUhq2jRxt92gm/71hKUKJIGkQFc0Nwqk3ImIv9Fjaqx+81RA7y3MF3Q2L9RKTA5G
yEvydJQe+WWOZm2YNnfXtb2RyX8QED9TYzbCNGs2l0U1REEnR4iim8VKqIGbQsEQ
4Fkwz9WvGdOz6YKBhwh6GOseGt8nBOr17gkY4WU0F7RKdhhIPzG9u9VJJge5430o
2N0NF/F/O22AVKV7uLdvdcIO5xxddKRb+y7y8NX3ykKnVRkc7rLhGNpE/JVprw/w
GJCVkcKDbIdDFh5iMFbEb6JmHAT4Lbr/CKaQQ2l9EejCbNEtqAc+9ng6P2FLXh21
ZtxnYe6wHZWaLAoPQaTzNZUgVuz4m9R3kXA2pz6EDelf7BtHtyLzC+wkuAusZRMw
gao5gqApGl7PM8t3zd7gK5IXa2APvAh5njLAUaw+/cOAbDVoYKM6Fhc8eG5CHelc
ESm0KBZCh8JOSTavNXKT9nhjW7FSXLYXv2iaqymdX7T02XzFRchUDtzpySOrewRl
nuXV5hIGYe1vVrLChZs0z84BNC75sQ64qmW2N5WsuX5sLGNCCywojPssDYzlcvW0
ziHygLERfX3GCY92fV2G6IaZSTnOoiX9int3IXXBGxhBVBmfaHkPbXmi0UEvepYG
24LvyPtyp/cv2uGF5odtpXcR7wstvXl+2a6/u9K5HhIodJUG6aSHpEtbZ8IlBr1b
PHKd1Pg1J2D485I/3BW6rv57cx60exNWlwMcCrEjnhl0Q8LI7U/3EbxHSM86U7a9
yhd7r1vlFNc+3c9YkZ4c8gXOVgvys6Wwevd6VcdDqoV8Dz1txA4I3ZSI2tr+fymI
ZvqzWzh25Kiu/ZgGRGJLQbiAFegAv5KRgUR3tbyh4OAaMgMVRuykwl0DTpoHtiu6
QZbk3me24WX5IiWk/WeVrnIb3HEM/bmr3/WcRnpQi/DrekDdlBT+moG3krH+FUYt
twWnboNtlJO1a3WfZwREibFwgwRZKneZpSsPT0o/yQQKZ3CjUIupS0oshg96FBmN
2wAQQhbic3OCQFL1IiwDSsKirHw/3Q8wbekL8cLqUizCiBeT4WdiG7fvlvZ7RST2
2biZHjoKAbJqHwfpNtuL2zoix2/Z8C6eWxvqt6GMB0vVq9SWzy60gk9LJyedTezi
uFZc4urcYKRsQOWHlv0IRFWyZRGWvdkkZcBL9QGT4blqsk8SkQC1qmKJBmpx2MXC
pOkrhD87U23QmbFACvX44aErXnQTaq4f6kDxyYcngyRih8n3kQ206VUp1QRPfUkD
p3WjmOtl27l+MFILFt4C5RHMk421oZ672AoNupbK+83jbARMFTPk0IoA1ADPZNID
e6En+Lm4bfsQ8Mn9IRffYAiLVhfGunWJzvrRIXZjz5atYhPI7QuhutnAlm6KSKhu
9l7inwFGc/T7thzYCBZY0c0wGSOlBKfbLMxw53gtyW1ZundkIeAS/RqF0/xI8W5y
8vsTB3WguZKlPgHR1xxF27H9RXQTUcW3SPidtugZgOHPVZxLn0GEB/wo4kfn0MZc
0UAtQbGQCTmgQxuzCTWOxAnBQjCmZPbb/90cp/R6/OP69qfO9p0/JgQF8xNPrFwr
qxc7r3cLginsDL22na182VkfBRo5fyIRJebHJeqQX4Gm4Ld5lIK43VvZpP1pmZw9
Ry7eOTmK9fCCpn7sj2/uoq71OStB1Jr6OPUbxGV3VhYf8oRHRf0zVJtBUdf9Pfm9
AavoisOCCRuBxTLthBm6OA4rx/X7dplFiySySsVZdYjJ/NCHRsyjcdac29m3+Qa7
XnGxheX1YdZf/UAUR2+uK+JVG4Q7NFmi2FVqoITMlMs6FsKMAf9pVkpncwYfdBbN
o71m5ew6Nhu2ozr8gjvjYOeDd946V2hl50KEy5mQ9iJWAURMTtjWjaGhTLXjJe89
7dHOgjnRET9sIB2/nKazzhmtNSDZAmwsXVZywaUCug1DiPItZM9GQ6bbpk+aZVy8
Rv5tFlqXNzlUnkJOyHVXHzURFGfpw95yXTpJyR/RhjBB9byH14gVZJWlmKqbWqcZ
d2T+immqH1h5WrtA6hhfk28rJkg6ly/KikOvP+HkgbM1uvfbH5NnhoOSbKz5hO5g
Orn8jlTczKH4ITr6ahpBC0tZhYieMPV+M8yWW4sBXYCVeol0GKDjH+Qybk5EadNs
4LMRfhp5AqvpRr1J995hRRXz7McYQDpYc5q2/ew48o4fndZBjKbJvqzbYNH+kGWd
6Gaa1REfYh2QE3pgqQmnJ6ysw02qgQ/bAWSOCRqMjzienDXA2ti/VVDsW17cwVaO
vHkv5jalChwsAURXpPjw3IxM8OtpsVM4JWKv8k/RiLzmRgWiiS7+dNRSPLelitKl
MfJX2INFUbSJruHfnHhSPnPEWvOqOPq01Wml7+gva77Xew0spJyn8ZYTMwzo4vZC
inp53aAPlZx3qD4bxe3YonLUVGoq2B9Ts+7NsdS4W64oxfRu7PIWxNi8ui2AJSgI
YYLg5herSEQK+YvHnryqDIVrjsIIEWeqS21wdjS7wL2fkuXVrbWCzzhKNGpuAnfu
StEZNSSFYN5gQvHF6xUoBZi8Ddi5FPu9E5qNsBNHElHL7gqMkfZ0/MIOK/vIHFDY
USwpsmFK6Te7tf8JrbOL1bNOcCPX2+rIk8TdYFVY8wEJKXqy2NFPjjxh8zrT9U7n
SoTFwY3eOlNa1SbErj2iD71VWRqB/I6Atm4Llw6BYkVHZb+j4aFRqgqovWEf6jVJ
1/6nLD8/NN2H0saZQchMym/4ACidTFMERElzeDJ+Euzzibl4ihziOkDHKIxnxst/
Uup8eYlKL0l4dY+S+hNDco5Wwh0+3Bs2gGXuoeNn9H2+MgXnOeKXz44BEKVs4QUO
kjccgvhs65ly3rIgfSqT2Jf0VSJVhLoqpVaEuhc6addgvLO6nQ6ALHuO+jXefWpG
FBWVY3Up6DNeTiqv1KmlhesUxRvHFVrvqtudFW2fAin+hNWbYs9aIf/RHreXe/lF
JUowKoZq/onaONcO31xJ8QSGQluGjffLlfuj0tFj74zHCm3VJ3LPL7dK7C6TdrvF
DyOcUDQbLcr37EO6vJHWdPsuwZ/hWu1o/ld0uGq6ulXVXEha7xaUXBcGW/I9+743
jWdIHZMO0DvIg9oRk1n2KIxLQoGiM7mp0KW7tCXwvDf3BCN3SyA+N9iB+aKNZxhW
ubMvB6at9egHwkRzTmiijbMmvUfDeQ1qhbzpaMsM3O4i+27CVJ/hvBV2l2Bv0SQu
hix/RtlJmT3oB6J+3yqSNymceJzn1nQ/QaQ7ad9bkEwBLX6tq9YcvrxtBp7z68GN
FGQKpB8EMnL+V3JbL3UGZ5diMmwHY9sIbkWmXA6TmpGOwb62/9aRODrBye0dbwTb
SymzzJDnD1thdNdzp8XFWDp9UihAKFFoDOgMYI2EFR7jsyV174H56hJIP0TdBQgj
p28zto40x7TU4EtNSkdvAEe7qFP5L1XC9xrrQ60l9kuiSNWTEHtK3tnJM9Tr9msE
8tyH904zFEGpY6aNYxuG1C4i3UYACw4YFlLfhVmXYVYVRpGKjEgne34D18wtRu8d
42lyQFx24YLoTpl7ftx2v5cekcMBahEd3YB9an7P8Av9SIHDGuOMHGe6McrNanw5
k73RAB3gxhckwXHLv+2uhF7V3BY5OA8SwoNCYivgO0Sx6d2Pa2IS8Ix7lWeQMrFp
Wtvblglnfvt2DQ397IMtOwAWj8mue4lFqZ2rW341JGGOhef11dllvCUSKsjDur0/
yqYIB/cUHD22XoWwnzxe0+QrXA+60Yk5DQ4lztXsYcbr7WVplBeD215Oc/e0828h
xhtCftxyRa/sHjFeqIUvx9aLWZRpp5WLdPwDuFAdBwMHzUKLQ1ecG+baR5ytL3kf
tKMD9HcGu/YrM41fmfETpESniu3geW1kkfPPk8zDlz8p0IlJB3xzZyqUPIKgeO/I
H8af+qjArZeYjwFf44Ag2JIP9C0pfFhqYjlHFPsVVZ0a0BOlXNT78rfN4fAiRCh/
/JFM022u9wciHehlu9X4MJSCeYHcALoy2h5YMDc2nsfOQCR3jOrSoDGAHQCQuTG7
djfB+NTiSq9Yak2RbP/tk1Qk9DIzSuil/xlIX18BJEwE4z1ywh4FuRg9uq7Z5MRJ
r1msL59VVMGNFTmYFvTwIYSaPhbMBuMoXbicOFa1LCypvLXt2NEh4Y+7D09/28+e
enlm4c/kAFMJPjoOcq+eIPyO9VeyPBZXHNyDzxM6skxuqC1tSYhwuRJ2CNUcqM8T
Nqi7cwsxZXx7ZyDr+PQ/fEYpC/Qq4dSk83/tFwZNkSA/f72isJ2ZP1fNc7b/hGxa
v+UQQxpRNvdrgegEsB1i2oLstcEOCadpPFH3b6sxt5UNYHa4HPLrM2/MHj4iRLCJ
MZRMj/Bomn1Fw5zQ5Uw7CjUtYwrvlRsvzyjmWfsd5488O783b+MyGCMDfE+jBSQE
NMV+mx1iMK6v7CwPmv9yiIy2nRBUUylZzIsdrGiAYEQHXDko8cZu97Qck4lE/hSA
QCl3dzSvddaerkaihp4XRDD5s+rYCaPXCZF8tQvtHUU+OwVteG9JDQmiml4n2Uz6
2i4OrpVO2y0eAjYznS6Qm1dgpJFWv9y/zJUHp4bLQMCOAuDDtbMwfPtgi4fV5Zon
YIaZEeXWD/JCKRRyoCfadUER0yyInsgjCxt+ek8N1JYl4TiwNYODK9WkUpNiHzS/
qXt6vLP+By1GGycGVtB2pxaUmgJR4ZnV910xBW8dFljgSPlN5qT3QLQdHP1ZG+EI
5nWpZFFLBzNugMcZVZjc5V6tMGBifLMPhPYe3XUAsT4UJE01eVCn9c0TScpio0Zb
eHiSef9JEIBg7TrYRcEu71SF1wI8/rUWEut/vwEopdyijLNFcP/jcUsQ/W10PWw7
e3b39jBa24BuQhuVVlA2qzyJMcGG48xTrB2oJh1vTNH3d823rHAU1s1cQrtN2msI
sHjf8nW7CrlNyHei9wmUv96u2qbcM0T/NgXxWOjHVmxzcctJI93Yhhc2Sg1GYTGZ
TkkKFa24EMKicCNP7ivouJweYrq/9FZHFGK7F1TjheD/dmOHV2IjOFeMcz2FzdHo
tVya9VCJQvHtjruI/CKL4p2wmHvPOBvFd2CQF6/F0xVb6F6OQV4ELkLLk8K1blSf
jIgg8XSxemUMTMZfgOxMqJgtdbpnshixZLPEovcu0KHSjm5uXzNRbZNwIZ2caf+u
c1EmgeJpov35T1u6l7INmOuQhXjUJz4KzGIKTyaOOHvzku3MNvBOZEZZOADo6zLZ
vv6LOwJjcm43rzVfpJmawvQu6y2GaIkF6dT5PDEzDUgzgP7x0IFz7KFKTi+5TwzZ
Jxw7j/XmqPh92VU+U7bsRXkne30bwNH2I5Y2Jbjve2rk4SZN3aTYqMB2L9qUW9CD
ENdm9OqlD3C3pZS5YM5q9B407gQNE8mZl/Lph1TKdXWRc8ohcXqu/WucCS17eDNc
QhPHiy6SHctxS60F6aapDZyxVyY2X1vJ0f//ED0jiuW/mb5/t+LNv+uZ/RvmfwfP
8xigJJTv064IDiQuUU9NoCpbG1MW0uFmsQDpaP97fERJKBYq++J/9xOMak1hxo1W
o6H1KE/nwO+Vh12Wg+SJ3TxjnwirRgyK79xLgpcuJ0z/2mSB852exSxatGX+Rrya
4o/6DvpyLcqmD96KtqYey0fD7MW65JTG7XvgFoXqgUM+IpPzC5JW+dc2IGahE3ha
n5qmpkAJqI3LiCFw1+OYYBKs2s9/axau1AcfOKrHFRmNNONfp6Yw4IZJHhwrlRWx
jNJNI8sMyEfqKWLMg1BBy3VhtNVrOxXDH4WkmqooaKI1iascFrCwQddb20n6908I
w6nsTryWV82GDEEVf9hVjtlBhQUmike5aCE3jXLJpmF0NWrjqI6g5qBVDRsb6X3I
PgpOo7tOaUObQrGArGg4bwq3f0wTsXkil7XUoLk0WmsVDEiIeKDrNjsMX+6KjZJk
g4UDaO27MO6ihqWD3K0MGUE4/4BRBYjFKEi5YHKtbKULv7MD4MReasjIKbROKXm8
KEzAJIUgXXKN8uXUSGJQfAEA3jMoRyIUTcdz0ZZJZsfwp5SAvz3c70orx/LXFE/Q
WVfLOOrN80/H+AAh2/DjblPd3y+xUxVKjp6VdJTaQSLS1MrQIJpPfIDOF3IhXkCM
GK7wwI8fOrMzsrDDpyY+oEAlz0TvVDWxtnaxLswLwgXKqwlmP8tiX0tHmVq3/Khh
eWlWxwRI7InatRR9uy9BgeVyauweCrgahKIYxl9OBo/flpn9aC6fd8qCjMN1cQbj
/8TbXsOd2aWuO+WKgN1feRD0rqBOlMZQy8ww8yngWWieh8YHhJ9vA8TiWK7rTmmC
HoMEx3y5I2klQbiFClOJ40I9xPSfaJljhZGlynyakftZExpy8HJxSJQpHPgnYg+g
lc6xaTOIO6QbyHuJiKo50KuAYw3m1GAhDJ1uktfqsYBcWjIHHbAXu+bTz9twNs9i
eesK/sXOvy1esgVsiTeH6Z7pl1IF/Z/ABAkDZCmI3EOBKuyu9O+DNatgDOD6mPit
Txaf2tGkyyqsLtdKm3zvw8CN9TWiK+N9LesXKFD60bavntga22qUmr7Qw6b+VMqr
psBEQFYFMhSuwGzwnbqrnJb2QTEIMcDyA1q10GNvt58oHXC+amVxys+7JX0Nl3sC
lnHtxGsUCTwU4IiA7p+Lo+ki/rXICy3aGD/W6BFg4vGPNL91JtX9LQCNtMF5wurP
QVvRIN2DX6pNO/JMUz/OhU+4mqr0NNfHRq09SSrkD3b9gKm4Puxx94m6/+eUW0DR
YEK5dVDGY8TPszTkiLUaIJOz6s3UFHeaAJ3idYAM6USBwNZ0PAvXe5YDBPEf2o5D
9/bTOpIGPS5aFbsv91+0V366RVe61AkDLJ6FLM8dN+u5NQmfDK0SsfK8BfMEYy/5
WGp+KyYR9VVyG5MhndeaM41OWUcIaKnqDfw3m7J4dnCQxzLIT3HxL8vl68oYxNwK
eTIE7X82dEMcd7iYnSosiH6pLoIm4qzjKYjxMQAfywvFjyBZxK5Wl5vaJ8GHU+rS
jfBxT7UWCwOOd5eVq4PW2m5uQRHczYC8OdWxdKsC5Wbx8l3j6B8D+GtD+S7umvlg
TWgVJB1EUGsQgqwj9sY0ouzxPGngZ5UYFkI12X7EpyVw710a+1jIhSN7vhOfMlki
toDsqpCHCHojyyQFAsPoyt2LKpNO5dfAa+umLMM8FwFPrQ/KkgHK6wZocfpH9mAX
xasdebIkgLDHsPs6ALU/VdO504XjQaLTmrbx8oItSrI9yKln5hSXzRmJuuO20Fz/
ccd0PqqRI+SEalHd492xcR0MEvOhiV93QLeVmzsR/684ocjRmImK3iMIyfi4uwKu
pWCeZw3cITh3bxMhCkEThZsg95LApw9PoQXTICrlx9vXQXeBIgEhgDaxMSYxgijR
5VgPiTsJBMiYDMVAc/mGIKXpkE935FwxldTBkFbdAmMqaFRTsIIAoEPoUB36W1Rs
LfDnMJwb3JXUb+Dj6p6bFmtWulhI7Y+8ZyGqFMdxaWsd0RcR2P4szdRmGyM+Am8/
5TYV9iLPnywVRYa/grITrAW5fdCRLfh1kTvjT0IE7Q3uWGla/Nx1DC4rk8Qwon2J
YDeeMJIrv6RfEtl822+ypJ1oFQ5dKKiYxQAwTfZkotorQEyik+hYFN7Qj7V7oE5I
i9nlbymdQdaD4gl09l3651d7MX/mVk0C3ZeIFifDoiX0Sk201v8FcE0HHkAZWII9
RjsIFAyPvs6imhfcMVdImvxhHzAMb1CKu4f/JzD/KTq/iatNhNvsFbMwpOPjeMwf
2lg0smdbdfyO+ONjE54SZQpGop+/9L/fv/8NwgLLVwyB3Jmh1hqhc35NX3bxZae3
OhybHdEfkEi3utQ8jkMP8ef2+o2PQBqlXBY9qKEBQu2WWiTGXT+czkcCfSTfPt+G
7BDNKPnNot/VsQvts8tPUTOnQL9ANdV0LVcnMGnLyrYtvBkx782Nw9jBKcKpfKb6
nHsTBVbTpYoGjxxaqStggECPlGmyJnugkMQcJLVfY/dJarODGvdn1pXBBGhYtTCe
DFL3O/x/h0pS2cZT+YAM4tMiQCeS7pigDafWOCEGah40OEvFqc8AtvW6hLhmB+91
4Gdd1t95aYVlCuj2735iDsxITl6dUM09TZsfnIYHuUlgNoIImGC/H2HSOrmgV2UH
K57cqA1JG65TwhEKbQPwBZFiXb/V76D2vPEbnemM2Lp7mB+SNdbU5nxvhLgnWsN0
NjLm6abXhMvic8okVm/Y7x+F+DEjK6Ql9yuXc3bbNYHnR1HiPEKL9EZ6TtahKK6L
gG/KCwhWsC2oJcmTS163/r4mBIN5jpyJRaDSjEpcd/mHYN9VvNv2+XdAOecxkPJG
uh8H1lJCzj3I1IAAFZdcya9Py7sdxme+au29yKxOoojzDbAjxc0PI2jtSO22ejos
1yE4cCqv/smXcNWSSaSKLZ/O6ip1H3hXxx2geUDI5o76Nt2zbZCfeIJGamiBuJNo
tC0rOpBt5RBrUTX8nmybtRkzQvR73Qck7hoESLkce+Bb7HFmRPMqfVMKrHdshfSk
qVg7E8M4mOsIFnZa3P2MvQbieo1726rogZe13VuaNKo6McsAemqirROQMX9InzV+
PL/vq7X4dLntjy6gRxU4rBxenoHUVLjutG38YDTKjsKVwl/8Z/8Z2wq/ryK2cp1+
foSjYTet/K7FOnE5Ltd7KGRxFm+JMIZDredjrgI2Iw/R0pNyI3r7CPr4jIcfn7vc
K6jaiUq1hJr4JPC8/9yoU4RlRwNeONaWj2gbuHh1TN/p1VoFHO6Ayjigea8pzJOF
e53UWOER//4byLyVG0G62BwCvZwhBVlnTSLgDpCvCVXf/brcdQBEZumOY6KXHG/2
ELh/weOzq00oSue1ifud0DY5wAGvXDRNGu11zDs66sp681NODMy11VX5vuUrCuuH
ii3swX8uvGKt0T+UQlDdDkvbcxBUz8lh/AMYRe92UQV2UZByevZUpWscaL4WdZBo
5heBzFagC7jRR5bHUK8hNMM+AzO/zAJ8AXWCdFdQZ2m18OYP2hcj8K4ZamtFNSXU
e6SQXl8TK7TmEN7BwP9dsZUtiwuQ2mnmtmuFJ7XE6yi1rF8rOhaMvKYz+2E/klkF
RxpgvTWsuF5Aa/NxRTXvTGxpHV3g/MbrIO02dbZTwBD1V+30Ik7dr3KL+KuohvSg
mrL6GJwNUzE5ZCHR4pqymKx72MigwJN8lSSsLvruW4hbxe8yih62nAKDLumB3n4w
gt/FKwDiIfJSdTdMKMvYzzc6rV0YhfZ9AQhwyg+hz6eTZTMfZIFTjBQW9ppzY1KK
oAcjVIqTBVpbEKFo6reIg/gszenXzb9g4R3sT+p13f2MKcq2Taum/HBg2gVxUy8/
np4nSdgVWdeIRTdKaT+v7Y1OWmXrpxp2AAF1cIPeTX2lX7GbOa5kKWoOdjs+5apL
cPBrM1hQT3wiaMuPmqcegYUUAtnfSS/MWsf4bYip/C04NGJoXH6mi2en258ER4j3
NtIve9H4AFkY3HzzvJhACdvjw4ILp3WBsjSd8oaOSXMs/avWFRSLnA5mr0METntn
EOTgNFl1h192T0Cl/L+N+3b6vFopu9ohSRDhyWbrSFx6J0eo2ZF+/icqX5ddpwYF
qZNLuv780tWNB5LymnuwZSBQMKD0rNSdhYZ606pB283/FGcqWlWv7k8T41Ev/eJW
6Qr5wiwm8g+83Jvqs3R6cSTg/rzHEZ4uwSdCHBGosTXhMl3D0Ss/OsxVqDN0Y7uN
d5bCLn9zwk3XkeodiYbr4uDETWRWK8XXu3LdUWvxFKBCGqrthoji/VBStor/L6LL
SimLWTvr/yEirsfJZMMaxBMVJ92KsznB7WskeD+DAd7pc0fE3FdwtGiCqCC860kV
DTGlqoQveuOfxDzDQwXbmtFtOWmSjWsxO1sZmXmzRaO5XJ+7bKmy+894rlD3gIvQ
26UNn1xN0AaMxwiRndU09FhoMDeWpmXe8qCjUFDwh9HoYhLNCr7dnEUpRcuM0n7i
J8o0FaJq7q7miud5HHjSXpvjGZqwgBJN62SIXSJoY/kWjS85OTbDzq5dCQ/lVoIk
ZTvGKMfxJiTvcXteXepSw8RxAhaDhaunnUW6jRSt4zRMDQGt3baeqBURo+K55dWa
D2xMGZ/gbRJR+Bvj52GuOVwmErFqm8wsguqUjXoRIUb7utPPGHOiMiDu1eGMF8rf
Yh1Y3Eksgc2PungD1ZnUQzztbleLdP82Y7YEFLT0XszSrEE0DJuY1fRnlWO/8JIy
l4UcMem3r2mG9CdwuNdUrAUbQuoP+/f63aUbhjdmeQ8FYcsig2sCR0IsgbzfHpL9
RyT5/2VhhJJXOeDtNMWbBgnMuVtaysq0/pZkVAtqk01rNqnU1avK7pQUz9JWQ5rF
tpJqwSuXfnXjEI3uCFjpFO/dSBBhfwpGl0aMFeb57c7xwG16HFIpSxYwQ4m6KV8P
7UuMHNNADVpEn7B9Q8ebMmssNY8zz1ebwLzqm6pGoEmKqgYnnoAG6gUZ4eYD6VQz
QXPMCSrpHAqF68IpGp9Qd1NUBAZ5YUD2ej8c3bYDfRcMZTOTaZipJ+Ja97xRlk8g
2rqvAPocl3SBWS1BlwdbYWmFuTCxf+hqunk8m2a+yNKtAkEpMeRUG2n+MKvuK3Ll
oUcz7MVoCQLUF40EOUFSolS/pk1HHGYxa2Lkdmtri/yvweWZuSDlh8I6D0IYhdaB
phFsJaHjcxZlNTMF22bVkQ9GyFw9n03vRnEdtEb7BkHf8LO944n7KWOUNFH0Nt+i
/p6x+qsbxA0PksFZw7kQTkk5p/f4gtEN44y0lNyPm4p8gzB2Q81DZ9CbcKvdo+mW
L7INfuk7oDsIU6OYL8xwIgfi9qA2VU0+cXzxRGO1jaLz9NlIPymdwrN01yLFImsM
12yGhke492mG9XwVnVsUwwib0gkNjdXaPOI0eeGGLafRbXjgy+xFWJzacwX/A/1j
uTa5qz52ZGsEEm2bhdF13BRF9G8N42ThehgTIQDe2pcappESMumfd0+gzLOpQDsq
Wkm9pqLPorLVA50L2wSWenJDNC2NgPpUAwFdYB92U2wblIKRuQre0D0cf7Vt0xkB
lgFg7/uOLNmh11LIs3ZJIoifaUcy71QhJAeBIrmuzpsmVFlE7WBEfK2czOd8lVvx
ynK1FSSvBiJpDvoYRAbpK3xClCOsw411QRQe6GNYUOH2ydv5SKw10TVChJmyX3Ih
neuvWxCjhQie6u2AVm6KI7+aedeFRAZrMcccG1K8fGDG7O/LANWmL2AK84rro9qG
P3mvAwh583NEo+HSKL2IkGg4GG8FtXQc9UPGcS7NI7yVC+eDXOo79cF04PxDq8HR
OGCK03TAhyh9DqVJB4dko1OM1cXlIUo9+I86meDEXDdKvQs9MjbkCYgmPpNdnCp9
jW20WXYw4k/kJlAunv6RDRD1tsDCT9K3huFEOKEsla3LH89N3ykjhXY0TQE/c9W4
KbZefvBVCg/Zth7YCwB3EL0mxSy/a4pe5KR6SsJgBovexyOhrNAGYL+tCBiXJEeV
xj6PSdJ8uBQ4Ho+9bSsIoVAJd5x7L+rKUWRSIoabHfygDGzFKxaLwtX/AlOX4n48
oaZETrAqmw9blSSrK+Xnicjp8pm0NpbI2sDINvrr2iQGsgpTUhnlRaepIcodnhLH
Jh3AWl1GFq56gcejIZe3MzaZjCIxb31X09ERSEXlzu66w8TKIu5UVmQefvbQTy7S
iZeSPnCaJAPZ1JSKA0cS2tx3l0aXfVn4Jvw6OAU+YlopfTxaTtKrKLJX854Mo8Qn
ADz8Uz6S/iW59bVV7TEpGQebjGs68C3Iv6cSXnZa38NVB4o8FYMmHJAdyS70CfyW
B7sGjKNETjGw8z8QBX8xJmfMKt6BXu4Eq1ZKx7sQ/pOakYkyRuTF4ioQLGjsuFSu
9JBB0E/6LyzqeOrZFupepLV4ePQllc+ybdBJDQRiBUJEgsorjgmpTqTbQGZZ5jbT
zdEEXQCyuigzimPkHaioKDL+kLueXzeHvYShKeyvYqtujHk9TQOmXPi6fP4unbuE
pVsm/H38tXtlVS7MBO6wlmVbav/19bSkCfRJUFWJd9p0j8qwmGBP+8cqhbQJoI/f
/J+nUL2rBuHidA+nQxsjW8c2yG+/vaE+YpR80Kpy8EigOK+VZLmUly5q4vBaWCnQ
Ym1e14CyEJb9Cb9QA6jlLtKwVQp2w+m2XmcPqUJo2ZlP6H8vS526mzA+ZYnSPLwJ
jroIkgJrfPIn7ZzZ+i82+VWLTTmmOpz5heLnIMJCsnn8YkdzM2ONaqJB794Kjqx5
MgMDkZKrSnDdxxyP1ROo8alJwhqOJgSTkqc4zh4Mdu1pJE0LwNno6+6tp8JcJh9M
JMJzV3iKDXmeixBSUXAsMNSCmYXoMxGoEInhr9TODlHS8ev/1Z0A46mNyYV7zshW
R9qHL/xJcMN/HNu9O4sdxA8vcft6IdTp5rNvbOYMOclI3FjhNobHcXymaP6PFpNn
njevtywCuFKHhw6DJNNhbfa+1hdkYlkXqby+Mn0/ZirNUuGByAi0jXgwQLiUBSJc
xC0rRfNgDixWyntRnfwH28jT9o9+SASrdBrfq/dcgZZh37QBSNYxGLFDJB0SkEXf
6JaYhtHy9rA9VOmclFVdwEHSGk01sq+1jp5LFBT+2uNuh9J6wUm+/PHwDfU58KYE
PoY1hRQRb/G0ZBAF0e6cblXw1+4tGXFXYzZXjkCd+gPzg41Kf85vbYLN3I37NdiI
yImpITfwXZPG7Hj479EgfQX4eWgbYeAQkUUVBE/v0bz1l4OD8CMTNuTzePG07vcR
FzA6J+n9YQ1yfKy0oy+ns8iEV4LGFY3GjsuackMQwwg1/bzI0Nb7cbm5CknczNtw
1g4WUC4driK9yrVwzQNFZ6RLjeYZ6aCNuW/803R8MVYQVOhH8JOkJpOdTMFwcBpp
mSdEuQkjv2XsJqHiX8+X4BdWdyb81BveD28lXxX5B0hJ50DuWFjrjx23nkMQwkUR
IUPUyNe0dCa7kQ4AnikH/ZI6v6LGo1SCYEhapzEMFBB4yl48dH/bLlRD4372pJHl
AuJyXul7qyAcupSeZrPERNqKuQOYf7nfBVutA5DCUrKTuuTuTjyXZdsUkWgjlvDe
cpYVRurxCJH6Jl82PZO5LVhpHSYkWpl7g7194YZfxxi1Xjn880ASA6unmi+Q0bAq
vFhDg40D0jr+zJvqK8imp+1zjE6KaPdnJdHgCt4exFajl1/RxYwjzezGpm0wfSoH
FyhvdY1RuqJanh2WoAd3ggTGKBR5U5cIccUcuw/yIHZjNWt+9CDzGvL8Ia+RyFHu
p7/3tLSV7JsjAwC9lzYzdA/cOi/nS3qi2U59Jw6TCYCC7YHPC1+lLhdIlO37LeVs
TfJf/IwyrjbzYMeVtnfdOGz3Yz0+H0YleCTwHHILFZ6JtLI3J3qZcYcJQdfW86An
8ZSBsyYPL7/eMOveCMGHHTdim5B6cBdb6v8qc/gT7Z1V/qtGJPpJ/SezLI67S29S
CE0Kc+Uo5BaoTA48UU1zAUjHVNchRL3433g6EgLxtEKHV59AlFkTN5+PpUBsjcgc
kj+Q7sb1MjIeijp/bjqGWCXFTa2Ab1UXx1bW+3FxVhKYS2lddkGsHbPNMnKs3q28
iEuE1E6YVr2qtnNT485Rrb6QxJh0++npgEZ26IzLF5MiTe88O4wfQ1yLs+mh+dxm
U0E34hwwQeKHuLIT4r5yhoilPtdwwSa3OoBYwLaUtbTRW40zNpixJ8mK6dK0aL0Z
Ij1rVogMOX/R+xXTfZerP1HXfJnwhoXHioHjnOPyZw0VouL3BDNX+jFJA+dQcebQ
6KgnKkKdGgfH50butciCs5RB9IXI/WfeyMOTKs3uEFFWT/r02HgTNyMgxnQdfw7E
WS+WHOwsonc7f4z2OlrOygey6q5A57QtuSfJIM/HuKGEsrWMy4Q+AbpR41gRbGOH
QIeXqBf1RF1blBlT44hru9SN1STJRmoptrtkA73XJkQb/kTYgPSMrpv0FFZJ4DZp
dCn+MTbZkgY1AOzoDzIPwIKfHj0wiiTANSepZOM6guRSr1qV8wLQ7zdXOiozmEl3
xMDvgVwlEOxl3jiPsPg9FsWBYndbP/vSZgIUb5LT8HiOYMavQimN42hWLREv6b49
Ea3VBMPBERYY2cZZA4Q16vhrmfWk4w4mnUML1lr8YjTYXe3gTO3YwMQ8YWRtVXj6
UByhUPoHu8CgWy+amyeHV88BiMf8ZKWzvWJtmbgYaDkOf6kIa4x5qEpAmgfbPWzK
aSZbN5OdPcC4StXe3bqBKWbAM5TtRvh9kVtXBpIGooA3nHW0MxPWTWJ4Y0j1amAo
VUj2R6mMoYUkvRuySSwLOW3+kNLNACWrgsXACqP6QDutrsnylVb2eqOfel3Y13VR
EJ02MK7G0uIS9uEM/JN0UjTeIjBpSFD6YVsjVo+pljQfCaaMDg3RPCQo7Av5gQD3
L+ImWpF36hLJtSEHuWF/LvY3jV3ynTwlka1IwiSCj1DoRzEyXYwJeGtjmjmB//MY
IizMilbKOKtsDiNwM11yJ9ZQSU+FsXGcGk2QjYujOIw6b6LW77VfsdphxZm8CZbi
7xsod8O6avjcXW7eXyAzXbtE0/4iE7EfdlNBZi3vXTOzswRnFxKE21UCMEFrjYb+
1WEA7njboso8ZvPwR4VnxhwAJnNySls6pIhy5rbFRxyN2MaSowb5188cq9Ezc7MF
gRH3E87o0G97udiLf29C7ZpEWHqvjLH/65m5x1IiarcSW2LUxbxHPxkbZB5W2WJU
OuTTRrADeoCiujq37DTDw6VdSieeLRiKyAsQg2TdRGxIqwarL5PccSV42CHTR1Ei
Q9gIX6TenP+ex3h4IuTePEtEc+ituIFAQ3JJetur9OfZeB8jx31vxTiImF3XQXWL
ofwYbYfAE0TNCDo7YFpT3HaWJBt+rqFrfYv5avm37ASm4nCbGTJLKrsiWfAI0s6f
OWJeIpwKk0lFPA3r4jN9Y7udNmu2mOfqk+XI0L5mcB3ZRRQ+1cVdzzcT0SJs4Tve
Q9lWq731Uc0EWqKlaz8ZAuShyKPzJoxrmFsreBYkpqD7p50RVyVE7c/AoPt1Pb9Z
Q/nIEGQm3Y7/8U6bgiesIT9SClB+CjXWOqXy73tnGSYXdPy5nex8qLvIHXS0TMWr
UQ7wtY2iLTM9jbmxiEg9v02bwJQSu4N1aLa6SApX+2+7svIw3EwQCmjCsgV0RT1E
bPjeXbL9unACyWIMwfjg5nwwlb1oJ4bfZF8a4l1gSUDmRBhsPhs2YhyAWjAU7dbv
t9Z7uLmFDZqmKJTuWWT6Cklj8yjF5omT1J87Y0zv9weQy4JQ3lnCS16+GEGKC35c
1o76jkdFFc/spg2I7M3wB73hL6vodbm9xOlliyeW6ogRs3Z8W5OO5MEky6jCVGzy
Ja5o5DOuqpU+2jdzpBzbMGtW5Q5rZp1eaVQgK8P27NsD0Ip/gl6uakJeqMM1v9KU
+dVOd8943DeUexIFYaNQmWPeLzRNNt4lwwdm65YjzY/Yd0S4XbN/frUD9e1PLooR
XVadbgw2QkoDmpvjUIhjcx4gJfQ8RYd955snqJTYZOrDiwptVcPTlu2yrgXhTFde
bOHt9GfKGILV09+FXSuzgHU7eA1Bqieu/K7z+f8lHXYUEW2UFl+FVgIBfNMfnWp/
l+fo3j0c4QpngWfu8aAYH+RlBCqGvZ4f0RAM5qKLE8Wm2G+dSrGBlAPF87JYGXVJ
yAJUuAcfc2U+62EtA4oZsyVoRe6NtwWGGb4oLVeXTcaCIhHT/uTDBJpIWA31mmVp
1KyizAhIDhDiJsocxHve8VsHPkgQrkRdnYlcMtZUjmgcwEurg+SEawvV3E3EVvNX
yGl0MfwZ4RwTpSaN/sS1W83dTh1ZrROKq+LbsIvWqtJzXJlG4k0sz5YofoXzgl+Y
Z9wf3RRSpOwI2QICBTWccC7ie3CSNe7iFQK7R3CBWq9PFqdPW/VNbTXsWLsX70Uf
uJxfTdNgaEX8BBj89/awJZ7UYectRHJQB8KTWGs3aWLKhnJlk9wT691M8R/qGtMe
z4uczoVXqoTG1+NOpN84T6ymuRKmIHyyhB77bJ1Msp3Nf5jo82ExL9MgnaNxgjQK
KNZ3gbnbFHz+vIrvTDomqlEbd7dmiw7qTbQaygnMGP2LrTr8/R5z7UetefadH216
knRU9xyOTXYvuJkPOkhQUKZQ/+zJOGeaTczAG5+tSCTFvhApFF4tqg6B09Gs5ni3
3/5a8D4Cdfi9nf2Nz7a/fD7+fiWA5gTu3/JnqjsT2M4+kgmHJYdySwJsqdAPQSA5
ib7nH3miNIfCPTRHYMOEWFKmXA1x1oJ1u9NdTuqDq8ApXkp0iiz2ItcuG3qu3n0E
KAI7/AlayW5LOD5Y4G/pqUs/0V0ETrSM+e5dAe7qTcQikuizMlBrhHrvJdpt09Jw
4Ou8AeB1bLqEjUCfv3tlYhuaMCYz0oJN813Yc27ym+9FmZ8yHzrCYTPrdp2tNdc0
/GyoqLxBgL/MWbJxMINrejti7DtMoWcfXk5TlDjgZTj3JSrIUs+J1gqlo4q6AaH9
FFWlMZxyoP0KOEWuvrFWbm3wd3bIjAGzVWpJ/M7h1YbnF3RNlDRhlRhXiMGpC8xx
kCiBetTk6Fqf/oudrhkgLExJPbBOm1NlsfObeAZUgbSZdiPQ2SVjhvVeaF4r2oDh
a7aq0X+anXRpHhtqvAuVINijQ1fMK6OO8cSrMHALAOf1mihW+IHa2XrgeehAW6Be
tZwZRHBCgVLsivCzkbORoSKmHA2204kGpmckiP7Rym9j+RagOJ104mYZS1lat+am
bDLTIicD5YTkFJhmTa3MwnXMBtbXYp5B6DVOdYFtWsct9FEx1pQww+K+urb1OLGV
2DSajDPDfxnrls8R7qmT3Edw+FkwvWMjtGG3sdEhVa2/+YONNxYQFQL86e+7d8XL
AhBIEb8faZ1MHrBMKDNpn3B6c77IwlH2k30+Zmy9bx/yZijXTxhY4WbIyufS4cK2
DEtjUrR1aZX+hAwR6Z0ax7uOMhiRnxfoUJP5JdeJzBdbglRg8R+xVzleQmrZro1f
MRmK3/3KahYxV2r5RXLMjJTVxcsYL/7x8rAo02F+dIUTNG92fguCkOnsghWnuJtn
6I+RiKvmPgz2aDQa51f5olsFn8FtJ7itbBN+tQsPYc7UiW8wPzY7ROl0RZSQ3l3Y
2HawBSuJChx3O7AuHktB9/v2oHbQCnpUHqhUmhiKaNs28pxoJxvVQRVczZeOFIn5
gx1P/kw8Eh7jRGvWtg2uNe3y6ggCfz99bLHs3NvpjSYfsvy8MyM+R9G4JyaSobz4
uzyfOKYT7r1Vechk2C18X92GISXJIyfK1OSJyaFumuKq8orZK/pZXPk/+tcCvB2L
b7j1xhq2mB2WrZbD2LwV0HgnQtGSnU3qKlG4ZBNG38lSReZiLz3OSh9MgKB4P6Es
3cEfRxN4Da92lDfKVDu09YtrcJ4Fx/6mSdzAn48eeh1CIHgTCAr8A4aKmP7QAX/7
nr4XptT+CZ0yGt0ztunb031F4VfNZ8d/wIv9/htlhZFbFP6o2UeNLRbnuYzKhY8R
Gvu7BUF7zB7l1j7yd8km73bialCDyRdpe/tje7GdPBWttmm7yCWr6s8IsU78lVL0
lgN8Xa0eZFcyyaG2Ifx3svyalXm1j50vuJDKNL8Up8a0VDQcrUCOxjqziG0iOEf7
8w4wIHem2kByEw2WRju9hpoOZbdYR/zfPGg3yeiE+0K8NI75vlqYPgEcaYW2MUtp
hwQE9I1sf7XkqCLUDA30itBTdbdV0csyMtCGkJepu2rr/b9gx0kdS+QA+gnFNXzI
3XwhRW6TqhLQ/ZXjNnXz8M4PT1BCocAwpKaVbKRQVMZxL+csjWwvJEd2NOe0CE2Y
q3cX+WtkZsj1NU+DdkClZAQCrJWo5Hh59xmznj5L8CdajX0UIVrkecb4RkkjfC9R
fTAXqxoQMiLriblk1nObcrGoLO29fCdE1FGAWbdVcvgqGrDx9YcpX1icn442MQ/b
CFPswFHNFOC8m6ynkvzjRAynZuFI4ZljNb7WqCyjgEvXkJN74cxh99KyTkHAUQY/
U1xVlgumBc0rvwsWo3/5JWDcmI65H2/B7xpqTm4eFotOVjx6WknfhO90lD+WYIX7
m2nl5HhC8nhM7AeuO6pkt2jHCV39e0kRay7rS0thgBhHTDEPgKB9JGItW3xsgkAU
BpBqSSpgOPQXj/6BBA8KUdoNRRLVFdcEXfDeDnN5AiPE3rAYLTmJap2yE4mUbCAt
bBdOuti2UL500YTK29JF8ohXjohdfzhnzJ1k7FJ5tYyRrtbriuwHutOsKxYVADUY
rYp/PWRT4BtqSwiSIt7Dpm9WCXixacnxIj1IfaAC6WkESBYZJpytBchbOwvj6Naz
3VN7FYCFQQ9ymoFjJKtTLec5X3Dqctb84KWlpvWMC1JTnBOCc7uHj0L9FujqO9de
2IdCbUiMGm7VkAbUfukdwksl5+Vudmk08da0UWy/tMgX7dZBDjtt+R/x0Ebr/ZiN
EokuQm0IbwLrkWmX2Zxu+ntouaDYD02ku0QBWpsFrTsMl7nD3w2xK9Qk22SJBzWN
mJepR48vVKESux930wzasFaceOLC8MBXcA6w9vsLTlQfPiIecYRONrl9scWe17WE
jpH1wjyeY2Q7Uc5SZVFsUUiIZQdGvV+FQJ0hmLW38qNjEwElK6wHA2cvDkatagDg
E1pEbx0lFyHoAErbg6/OdWtf7R1u+DtfkVfDvo4DfmVRYXiF8y1uQw4CUGFLgQcy
TC3iFRccTFysMDZ1qRWnR6f2cta782WeIsf6QbZmFWirOGelwLBq4RimXtmDBFoM
WZbChvh5tGVlQeP88B2kg+pDEO2TRQyzKxSm6gdc128bFcJP5z+h+NgVqzi5ZfGL
nJ6AohmhQbSKZY900a5mGOHcXAXxv3JMeawgqFzGS7c7QQPgvskNtoziozyNumWd
XtGXPIRJyO3/YqWqfp/vKx8V+hPieuyWMAkM0LZjVO2qSDI+HhXmXz+kxVub9FM1
byU1Yf8JEEGMQ/s+QbkH/0+3yYGOqCBGZqTBya+ViJ17ulmEg/rsnk4aKeCmludE
xJjdPEBM2c3p1kxPfXhFd8/Q3y6GlQHP1qoBKZPXSMt/R6nS1uPQ3EqW/4x8ViLU
/myl4zDMQJOtg7mV0IVvs82sMPgOYHpUhvIdgIBZuM1iXNAnHm153QZbudcl4MiM
EAqvvi9s957LjNPT3sJblHs6j0EMgTjM4fgtE4cr85YMuvb/M54/pAMAQfEnkXKP
+jtxMD8My0j257Qtf5juGjJQMgGn4Hir+uy7PtC0Oi+ZhWAtRh9nB9mS0cDQqBsC
ZlhsmBETWM5SQrbQV1TMBcLBPt5ZaHjSYtOsESMgG34fEf1Qa7yDl0DrmJ5aHJxR
FCrTDdpdKDnbD6f3RZWvxhlHYEBKZ+xSivBXFDeXzpuvz6sike9kDmsf6Szi42uo
Sp1wXNUH+iKlGBxcjKdCaEQb5B6P+afP4v4FHDPC7qQZ+vcS7H139ymEACc/2lN6
leWuVaAlyS8YarFxrJY21WTUqvmpMT+qPdEg5ggl3LD09Fh0uU2c+Qn3vBndulSR
UW880P/OLK53AlQ61yvXyluMrR8XkykRswTVpe9YW6B1cV84el2r0+E4a9WW+Tnp
rHfxqwmfZ5L4NTKpkSt+Lewc/vDRYSgpEhw2qeaPS37BkQyW9jUdd1anK3nq/dXt
ufWF9ITWd0v2jdUUevYPJZt6IS0r9AuTK7uL2T4Iz4abFmegSq6+DTL3X2ob2X5j
HqE9OT2W5TD+YHpchPsCW7bDgqI5+GGqEk8YW0xSYLz1P9NfJY4/cJ6PexkrY/PW
QX/E4hZ5+6QzYQoI35qTy/Oj266a69v5b0Kw+G8Xz0atMb9wcC/8sJeIFwKxEDMb
0BrD3nQGauuDJ22FsWNdpIiuMB9Swv7IwwU4JTlITCs9yOZLn1uZoCDPL7JrocSp
qyqzJv8BOiuZEIn+HWsieMA+XRYNUfipSkQgPxR+LN3H06Op4kjTWVymrY6Iz4r5
EHnPf6DqoPSmqOKeynBqxKGzcdpo9IzuFsjmR3wQ4hfmG38rBAxontwcmZM8Irk7
9dOnIwgYnfR72wlJ8OgT5PtgaaJH7LO/y6xNcuqX2EivATpQSlWVA7/vLQnw9fFf
zlZol4GPykqHOPJRWSEDJcfz39Hl4MjMN/YM17PYZwQXnisvB+gI3QDCj7RS237R
WOn27aAdGl/zQBHkvBiL8Mxy4wlgGrQN0DyA3+xZFRLl+GiABKEb09YVdySGD35a
wLFFqQU9oLGkS0ALv5hyfEhoGS0wFgc4zmWrx07S+PK8Hr1L/kjd8EWFydit9sZj
p5Y2toitkY/RPIaPiclmLPO1ZmdgmgMs61GHBhF+Bmfgskp85PQ0ZfFXHdpq+PmC
ICz6sIrqNiovgCZNj1Wilg8vO1IDuEtsLFCVHmphxeXJpkvCe0593mrRr3Dh8gcA
nleRvBixT4t+n5/RLHTyAlagsTLGBxx1DWj3wNBfzPihEjHfN6TyklsvFBp7MvLZ
1LpDO5MLF4uC3ad9WRJs8+UDWROM1ZqfzMMDis6obWuLDaOVTW6b6UeUIals43T9
wGue9gTAvwxKBwHPNNLpIXY+OcbiREhBtsYwqLZlTw+n3OQWCOIAFsjHJa9m5J/9
TMlGzW46bJ3JdTNmUR+KlBqUKRY5yIddBY9oKlO3bIq7EYS/Rxs8n2dG2wz+Tmhw
yxBJJXVES2oJVArgbZfge8rv6vUiY6pZEn2Aaj/TPXtM1fmge0AktpZHZY/TPrL5
oWbUQXYNg3l5SeN/ee+5258c94e0TWiiUEE9Pj79XltcNxjUK8YeI7ezQe4x9uTk
QDZav/YcYCbnfEpHvo1p48I/ppTqBaCRGs2esmmePulfft/epuF8356j83h1CRQg
nCS09YJg8UEmTK82KEDody8MXzJVLzJfpH/Qq8t2+Kl1Qq8tNf4+IiKjNdMjoljM
AD7fVhZ3BHs1pmEt6ohK/+ZWwkVZ4Ci4JolHyNQiRhHKBuvLVR25nsFVyu8qggpd
kcTZdyvUF3EXJkpq1QfHjGRjJdokZDm1L3RkCAqKWAb4pyGtSlpo0TnOGXd6FziP
AdwQcH63efSofl7PFqmoe0rByLAnpICY+7P976jO7Sz45NGOBJI2P4r2dwglwjCF
WlQCZew1ZzCtRh4+apQGKcgg9BbgWAq8ABdh6F38DoSuehM5uSBQn/yTM3Ac/myM
j7DJGz8cFTyhd9Mz30MigpQBul+68CYAHRjaWj1CMCsnbxMVwvvDHVDE47xhdEms
RLl0Wq71BB52WZ2neDqDFa3IaLDSVfzzE6m5EWqL7S8jIjdQ4SIIMq/RDEKy5vn9
ozRb3fCGXsl9tRaW/PdSkZ1uI1ag7JvYouPmokXhpuu//UyHnK/Gq8+4UCmwSmPa
ZVfKQ8KU8JZ0kfFgYy57TWmdwTBgTMTW18o9H9BFVq5MGCdKLkXEnEhbzsE+EiZz
hAB21PHzAGrDg3KSbZ8iRIFXnZvfEKw4GKGwHFHbRsmAf0yLmkEGW87mP9CKrk71
Jl4XEz9VYStJS1E863dIri4XBLp3l1xU4VbnVe/4EjCC3uGWo0qzvrN7NTxgrCyK
K5TzT2lt8jDpKcejvhNSfl4m+Fe6oEoATd7rMfymgRtsQTUHqw/S7Jr5dda2ZVi4
8Y4hd9OcngF8S87Q2mCm0eOGo2T7YgbeqmFWLlGk1rV7lhCzheNvNa4bewlxQtVh
jaVQCBIZADcWcMGHEH2ELYCkh9y8wJ+twtu5FqREqswM5qUQzkk9cAc3DO54L7Hj
jiPEiCXKoqGqTtdY6iN8eMD0kciNMe1PALXuKc0WKdxZ44gsGVI7CxVl8waz0kbp
7Soe5J+ks3l7Cr5SnYgCphQDjFOn+Jku3KEClSrPwTSkY1A3L7lkEbzS6OVJXMw0
c2R11sSrDIBgkQutlGySBNdeussP6h/B7FVI7STlBFnSPg3Uv471ldpLkpX/bBZj
iMbCRtpv2qN9FVBxETmjaNg2pzn9GoNHWtnZ+jFWXC8NXJdBn28hcCFYWXs+wWIt
mL8ifGVhZjrMSX+y6fTZvvjn+rFYpoKnbGazzwZlal+2eiw4bchbMah+SXAM8pVs
vhCYzONJk4H6fxdtzxByagOxkMUl39EZk1i5WiwbfOtmvZFeiYOj1raYI3bHm5W9
CEhF+zBulp8s55KrFZfSSnaiVKwpIuOv5+bmz3boYTVUsvuPZ9lMv7bjLip05qem
OeFMa8cboNd+ePXGtjKHYF/Q49yt9HiOAaytVqhkd45jnaPP0fYAPHXitPv1sVN4
9cd87AN/9e3z/F9vbHO+bf8klRBv4LoNkWcB2C5pAqSWZ+440aXCPXYTSAqs9sKc
aBXe8m1TU8bzY5SFzRcCSZAm+FOR5mOvB4BCufPWLdML5LwzJKEvcJOlac8vQpRH
yydoQgkPo6qMAA1aS+lY6ZxMmavNshBkXT1kWLp5ZZcxnC+hNnXyZI2uL6o6ysqm
BvgfSDCaM8FG9WEt/25ll3abBA1aa3KSUAUI+sryEmXTLW/rpB+wjvc+u6nDeiI7
9XwghM4dlfT0IAu/JM5P5Aw3W18jj/M6R3ybZM0K5Lvbs59Fpmf75/YK/Qqm8joT
/nUzXnL68GfwEAlPjpN6iQIvAOk80dtwINF3s/KebjkVrBcr14H9cZupcBHOiNC0
4Sss04sHfckQRZ/wm/W/PQx1o526M9WcxCNyUvJOk9PjBOo83X6+7CbDObZbv2Or
uPla/2G0/mrQ949JG6p5A0Wq1fQ1ixZMKh2mhINvF7h++Yc4XluPqQqZvWm6g88B
TjL6Sto869Er/IYXm031kxu/c/9MdnFimHLuWdMyZPoiD6hC5+0RDOIo0MjBibzK
TxYP0S35DKOsgfUTZMsCLh5aMF9CJQpNMnRUMrMz64aJ1LnbBqodmzeEjjy365W/
cOVpQMC/C/bpwDp0I4CSCCk5RW2oanUrQZcHIL/4gPMkCxSrKJ0z3XrGuUVJSiUN
nCXaOU9ITXwUARlKCfbqtZv65IWGECH1b8L/tGkuKNrOyiPkOETm4SpV4PvGQKrs
k/1BnORL2WqrZcah00Bd35K9Bm8xx7B04U4Q+OVKuiyVAsMXiSQkiyES4Icx+52v
SJwt5iYr5VLzD71Sf3MMF7r6Jz/EImKOPmEHI/L3oU48tKaAZ82FHpx5vdH1J12Q
H1qTPcy42AKNG3ov37NuiYvbmYXXb7zcBayX/+vHQAslZUxO9hP+8FadzYxXOL12
p5XCeIxpXQjABgCDexxOmVz9uWPTyw1/FEtswv0HTeP8U2Pn5+oVYirpEE6XTzs4
p0O33P1FUhJJKCV+zH7+cDS6StZnb8JjMdHEf1fbTVV/bpD0jjTG3p1166zDlapE
XaIXNpafx2MuN1CLlvRxxbwDLehjBjqMPT3UUjOgKgkcGli8y+umDAT2m/2MDNG5
UCiA+cBsUEHXPHc7/JqY2P1q9jfCfBNdzFF0HpYpxNU3xZ/t2DY/JC8ExFy7De4u
y9tNjMANuVtLzRAyXN5xRTIAwrPsR3wjbDaDmEc63b0wEk8v/NaJsxPg4cQl7erw
ZuxssIXJ2htanDPFLY91V8wD4ERzVArCI3DrJxKk/uWyFXPtSXeka7qSPVsruNTa
N4jvTrGO+2zY8YmTVV/Q6ZpYbtHj6kybXZH0bnbayDlXwHIzV1rFytHBbPIMMVkv
JCfyU6eK1MVIF7KiXhs+w65aDDkxhA7vWOmVzUPptsjcGA/F0cUMwZQ+2PrngyMC
zcoBpF+WGdXXtuWMx7Spz2EDWjzs2OJY7/3aGQWQcAkvxnq1S9A+BybYeeEErms9
tc3Z8GRkYRYlMHRqMfG8n1/vvMzUomWnVIqT3Nr6Ch+e1ycv+7XLFi++WuaLd/C7
q6MPhqRQ6peAmp0dPdlCtXyJUc2RGT/gyueKvCHJW4QcelLns/yu4LTrJSKM76cJ
OsWJl5huqS1d+BNJviS53hejz/zVmi91kZDNcbfGXpnKTYLplThb+H48K8UmnXM9
H3CCLQ2wAkfT+0bELMVYNdPpTcigh28IHHBnb7mI1ZpC9iWeaDNQImxKCvNLnSB1
aWkaaq09WirQRDJvF7L13HAW5kGSmScbxcstS2tk5738XuyBTO0wp2jaOhBM5qrg
rVhGWdYBk6Zr/NziQQDK15vSzKR2Ufcz0PnQ42LJnJ6n0M56QWGwXIWNqwMW2ZTm
kXPIchFNBe8Gs/edYuvNQb5G29OluwbBByfvhb6yZpF10GvQeuodO2NcsiCyp0Yl
8p6PYhivbf3kW7Gt4Ep5ByzAd2tBhXB2Bhgxr7RDwq5uQtNdXpnQFDrhKGy6Ha++
jREOCP7uqfsV+DFdYwD9BGF8PthhOGo0oQL29R85WhQXmEIplR9HU6Mkjy4PfKBT
Yx4fe+Ek6EP+4w5BcI0wyZojYMmZzzT22mJZAezwdZfR0wXHiclq1kEaN5gbY5cf
bh5Aqplx87VOmFrcpjXvm56bjZ6/LqzSsUi/W5LlPEhB8ip1B0P0LiqJqzdgM9mx
63FT3Uh5ekeixSlqa7QD7Mc5ZhoUXPtFEnSSsqgsoCkirjZ2Id5+oAv4jD6+wsaY
lZGuxQumVR8f3FprUijhO4wnjcrnA7p637MaexIgqvkSaNkBnBD0f21ZyqD8WRTb
P1ltIdsiDxK+XtXtwftoWHGWvvWEgPGvPzMT8qzGncN4gaptKYvsM8KfqA0bnQg/
BxZtIabjhg1JQZCM5e5QhZQ2cX8kmK1esM6zdIzsN+Y1d1TN8JRjf4uTIJuOlBpQ
/yz5rKSIIF+uHmFBiuEANMuZTRozwMNslpTy3O4QZlX0MSZWvMMN8yWs/smeONaV
VqdX22mxjjN6vgGp/IS4AUn1J6LaiUc/9tA3Fb3UVcOvkEXiFg4QSwj8LzFOWf+o
+7IEqDF4sZQhfMX3PfLfxur2s7OPaA0e/a9GW2DW28gYvh458+MUbgdeQ53zcQ3T
Xh/zb8Wgihexddj+DxARsmH19jB8v7dy7B0vv0Yqo5cI5YhJ+HPnvkNyOhE1PfXt
IgLiLYjKrsc9k0/4QY5jVYI7Xpv6HlSsy/395Z8FjNzDhvXPsbYwxx73Uq5bvKIH
p//2rWuLlW9C7x5IXJp09pHBh0MUWc+TSO2LOG73D1/VCkJU2KhGDLoOV8q0ZR0h
p22zhhPupO3wgFvOhm7C/tVQA18JTehmB4aGilCDTHyNu9OjTqt+2xwQhUXI7Uvv
fcW9yajNKiXS04XT9HQUHzAwbCLwx5wEZJ1PDL9rI9BnYWykUtBx+lQ5AuLbb3/j
cO+A/wZbfMvr86g34txJqAo7yRg5g6oQzhiQe2IzUq44C0nuEaVPmR09gXBHuAYC
rUY8fPvswoeTW6jGWYxAOyDd9ufL8XtdyrKtFmDMDMTDKM10dQPexxcTu3UOu7sR
6mixUF1VFWCrTAVlvmnOGZk86L/1tTEdM2uKy6fE1h3YMBQEn1B9yiU8vDftavlf
l2wEEYD7LI+FrtvPIbKrflx8FLRyyb/EJFs20cf+7GDEt12XRwofQI5Py/lJi+H8
GToKnF0/sPb+Peg+CAZWUwkY5Jae5azsB8DmR+CKUZDTZ/dvJHarKMhKnVzcINkv
E0CZ37OcexWdoTm5W9pc1hQQX23q3NQXLrpmPCasVYFo8apNihnbOggqy3mlx1eH
gMAcDYbarq3D4WT6hv96p6/Q+Q3KtXerFp1Mg6SB5j6+Sc243p7TTU3qDLJvksZy
blitcoLp5Nl4KrqpTSN7SAAwD1si/SDZKvaYKQJ1sQdtvhmNKq3Q0T3zCa/8TABg
rn6dSNxGzu+yiuTbmdOddsjK9xmfC9iGp8Hzi/WTcKmDlG9WIKUXVDh+74DdIqtj
6yWdqSXSJucQSjSMB/qG0/NPyDMqEbrMxIe65DSdEGC3i7OU+TeM3b3tetjuyXvN
5LqSPyNwIKzempDeDm0dIcevkRhysDBRw1xN4wbsRmX468wcRTeAHpTSH1EfaO4k
1du6aILzgQulB0onrA8HbipkDYqrwqfiGDcuPx//QZPu9nCT4jkNwY1nEONfgHx/
7dnif5+Qcxd5k/enW0AwDQX4hH6Gc3oVv4N8gAPIetth2B93m8JQN7YpjWrYZ++J
Znd3DPKVvLi69OINPo+yaEcfkIyoVb4zXVwNBQpqtl0ZWtUAQTvYmI1FUHut910s
OdQbv/2RE/8ZEA7nH73z54xAFswReyQyHmcKUq4hjtnCan+36Zoxml+G/98Qzrvz
UK/MC027rkGCvMICwlhwvz4gqjzK1stgOWf4pdhhqEu10MmGGkofLxMcsJgFs1PB
8Po7KmuiqxYEixcg8XCJ0PV3IfewFn5G1u+g3Y2DarPYsuQJtuxpyJCoJfpKf95p
5K44oqR+YALivgZBM7VGE/VSagOcb7CgS5mdlKtpdDfU96xoL1NDVkW+cjLBfqR8
/WPZzCUHGNEQGtHM5BG1FMh0J443wOgxko2MwR+cZUOxFDUpL7cUtmPUTnujJP6+
CQ5CzQhD3FaHD4PyYh/lpvgmwB9ASHKq1LkugftIXTxcJKFbz62JNUgcBpX9lN9/
JEZRBspTKLN18jmfBJG2OZYZXFTsyQZPk40cR7QkbhUG7mucaKpsUL5BzbP1kwFA
tJ6hwClBusCXnNWx140P0QW+J2IfVNkTBvRya9BEhlYhwfz8kkRWAs1I6SUr1OgE
v8tiRy12gSMI3vONoYH2oQe9V6KbxVkQstxVuYg8YyGdHH6+C/nIAHI0QHdsMLOb
NFTa1zjhPgizPXAnnuq1/fS6t8zixAxpGldYWyEOf/F3cFDJGOYSyqFlkkyD8YLd
StcxV7dmLK6XskhlS5NYMjGkM5BQQzRoCmn22fhDiT3LbTOYZ0xbtfObHWKbgQqK
oktIvDgMKBk6zx63jl3h8c6zh0VrVyBQrlXcwbZBtlVVcKrjXKzoUYE7Xj8LkVna
/CK+cCHFxwpkw2hZI7WeAOsI7njBZUc1zKypf4GL91Z3NGJxoJs5nbdSCcA2uwye
R77Ig3B5xtz71A6WLhQBdCaT1q1UN2g3zQ0ZoVk4LbLYfVKtlFYWxUJKIMjwJgnV
C+SN8S8VSJ4ejRuNcdMPz5y1dRtASG4hkMeRlsu9eRxqwSzbhj8iA81aiCd/cY+w
8i1jxGVyzuIzpJcQrWE0Y3DcbYcRHakjMzBZRfXE6erVfd3XHTjYFjWoZlNTSWPV
+tul3OSQlszXZkoc9xnRyx82AfuhdotlVqkPRvDxUWT+Ft6ULwQLWJSu91biTFhU
tWamLXa1fXnyxmsR/5rQhqnI3f2gbJoJgceHmkykvWQKZPgLFJHIUrTbyG3BcD3a
KRe+Kf730niJeTEbDOV5T2tzRe+DJX5MfZGf1nThKzcvVvizC4ZoSpO6iV4kFMBk
vP+UCLlniOy8WBLVeUrbQXVZBBjk4M/82JixPnoQR+60dmqbW3llti3DssgitZOX
e/a77qmtRNgjcsoyX4p5J6fStjRIMUH0EfFb96xyN2WxQ3Tmq+Dg74gjky81IdDB
TQoFDzro+WyrpiF2iIUM8oKbqVdk4l2wPXKtLwpMz6d00kAMlbx4lijExvOD3qK4
fYF3PQDDqcGx2SO9oGclwj7lyULqvAK2BrkfRPTxmuTExgcw1Ok/X1eDbq2G7zWC
IqUBnaHOxb9Ij2Qjk+W+DMfABY+sTJ/EFDEbsLPifQZETue76U3hgDFDJhMW4ysR
pZRlX3m/oZWtAh5n8cp+O82UjT9HUjen095qfk8CWvwyvB8qQu5/YylJVm+vi26Y
HxVvmVwW0t8hgdkVoubCLWxcdsPixw0zrV9rFcdxsZic9usOmjaTE4E7X7QJUIKB
iAegyV0GdRaSqVhQz6DDTACjl9hvIJjsje9Mcpz65+NVt0Z98Cx2mdS7++eeb0ml
wWjh1aGG1ecQpomYOk3iV6A91JrKVTrml1vt3LNySt5FE8kXJyof129PO2pAC5hM
XLPOP72plQ5kTp5o9v9lrBk3PCYqg1ysSfLWnnKwzUUHIpsZtWjfG7rJXFO/xkqY
O+AjOo3l/pa+oZrs+oWPnV6AGZTE+UhkDLFfYyWcUn2urh7aJgwz63rVzbRQ+MFL
MtmrlOueiO5EJ5PDpITTXHuU3mMUweyAg1zoCCtKAvRtVa1qqoiCZ+/Y53OTTmx0
Rthtlos4AMwO04iyovMaSiFOvzSOa0KlgfsMzwLxoxf2x78KhqvV7avYgbWLeJsg
/FwL8rNZh+l0Y/Z7p6VQ2fzyaLkSlEcyTeXI5r2lJnuoECzZgAP74VQ1UcuQfkoZ
B21vZYvqN50dCeNswBccBAekO7agG89rxHXbTxptyyOLAq98w9uc1xrszi0xGCaX
MPvSEsoOBGiZ2dx+a7F9FH8SZvpzwn6tSRgihjQy72GGuL2Jgteekc6Y6PKIMX7a
JEyWIIRz8w784EFv1Oqzo7RKBkpM0GBe3XJzcckPUIeWC3fvu8xYyW65LO4vH1AE
WIouWer0cFpKhPewvV3POaaf8LBiD55Y16AqlbNoPUFct/u7L5ajw3YgZ10Br+H4
kKVE98Ux1znAEY6Ne4PvEc7i6Nkw0S79HcKIRpkjrIxOS71JSQnyOy+vKj/z0JON
h0iG3CtPEotwMStCyLQ3mFZa8BF7QGOl1+up59Xlj0dZWssEc4HGsd/7h8w66E/W
IO04ularweq4fikc+NEYiAorktLqu9F0PpicQ8sGYa0emihKOzH+5EfX4XMFf8+w
6lMVbHRvvNYfd3JJkryF7jcZOQNyX6s5Y8VvE/+4utH+AYo0/aQtFPQUSGUWP1FK
5R4pyqt+OYx0s8ptViHfqk9R1vRDXQe8vvEYqGB1xoct+ZcCzE+8yZb1P7EPQOB2
r6/H12fMXCrXUQQujqa0k0nO3WPEZkIHz8rcchbWuOigrPttTCRBOxUj/SXHerZc
AERJOoe/wGZxtU1vJgy2iTsPTCeIGmWMiLLvXk+EQaeRLVYElpRSrSiJycsDg7VA
a49uPzhC2SAe9ELpFM7Y6healiBAYxvywTi1Vo4DupzejBXYI6U5e4gQs1663J68
cSMrWGWMKcqMBEV+HN3+tx43cF1TShGV4QyGnTpDUMsIL3jIan/2zq7hxClS+68T
LZsVICYSvbxuZKM4Lyt+nUWvsrl8FePC4u2sRnevDeqr3vX8i1AkeWlJhTQU2jo/
kMDHljgkJba19gZ/uOwkU+zBFxme6qbaEmlIfLtAZF2uRNtKg2jNqa1MHrw9PNBO
ph7dUNcUSIy5eF4RAY+BKBUWR22EaU3q1e4SIA+CoCNpXtJakFDH+DPB/8Atw7RR
dnTHz2sH50tb/BUwaR3IgEaQF+IN+YxfCK7wIbDkKZrxZ8PEem5uI2O6S4GmeN1E
BZy+0Jn4Snx08Iyf8M7MRvOBG8vVbD4QXec0UlyR1teHbU1UjGeI5KvKnbozqklO
lbmt1Fmx3ogrMU8QQVafCYiHAsFJroTmjaEfOSterap1gmWghT4vrQbN57Nvg9aF
i+5OHbj8Z+l/EazT3eks3K2J8dUcO7U6UwP7szfoPbNR7KJuE5b7DWwagkUgqVTl
w2rOlkF2dakWLFz+B1Zt5Llyh5RRCQ4lAcNXNSaFFU4K4D0gNHIz5SNV+Vpbaa3S
ffwrumghDp+5VDPHEwU483LHFs8colDvIxQ2+dwECiPzs5hb/5cs/Ci5gdNYVR4J
Qp1VTUF/fzb1IlQuIe4wfnnA+kAxuqBGobOSxY42jZOtxfuiU0rHJEtFEi+8ZM0V
xQAI36yNujOOs4R6o0ADldAZwisfxu/rCJFQaSpmFKppehsaqjWlR+8tZbaFHlqh
PEDriKRyFy0q4UgmqVCQjsDo5vRasAeTyVmDKSQFax+80SINU4CZqczS5xCKWU8N
xXeC33W5S1EWE7FgQq8Kj935jMVwMlN5FdK6mtNM8dX/+0vFP82342Ez5O9fxEWX
kmql49Fjkb8ihNTMUL1hvG0y2s73I9aXsRxLaHcURL1M43bmPcuZ+RkBg+mMNUjQ
zbtGosal4hl9sYHjHgk3cEpv1FwDczETEcNPyFFqVdT6q8ahYkC7Z7VW4pCc63Xd
6OOHOlqiT+//KRZISWoM9JmJhMt6tlDwV71H8CVAJzvT/PzvV8APSIXCf97mBdBZ
xrBuWAhZL3lke1ZBBR2ChYFvKAoCjP9vbx5VZ7555KiI6/n8ztwJdGJ/PPH9mcTt
rPp6m3NXBOEVx1HToLIUwYXHwU3e53M6RqWNnU5P4G/O0BYKF0hqcx/F0x8D/Loe
2xxq3chucyftsiJ67+Jd1YhVP5pZaJqBI27Elp57ZyAeJHeL8M6jpZT2lYo1FWgc
l2tQoUeXLQT25DJuiIPn3Yn7mA64lKCD9v38WtvJ4JpiPVHG9Tv5LmDTd4JD77Rh
ziJkLySaKEe6L/VHPgyIR1KiIU9l1xIXUv1jOJd2xLD7F+6HwR+Nc22xRcSKr2oE
YQQVqHr2S4gZmN9X0sBZPIyJm/KNPo/wHZVmnPERdhurJoMI8niTNhIR6lB3T6Ok
qI6eTjOeFs4JUCngQoR3MeVWl8Y3d9XihsDO6BWR8YEZvzMIfdmhAz1+yDhh5pk9
ew2tIUvhpMvRIApiqpD4JWTOTOFbe7PCJ4KeQXwvcQJQIyGBXI8wYOHoAWTYagtr
R414PrSNGk3cTYldmHnBmDCTe+9lll4y2oTVyKLXe3Px/JgfXheP6THSHSTPVi/S
w+/+VTFfuWhXKuJ3grPdXGwq/lqzzlhXzrzMiWu87YTEaz1cw6gXL+8IJ/s1u+1q
wXvWPmHsu1+4TxHN3lbqYdMQh48aD5eaQmBqthB0U9s8pMOpM7Shl+/zVzUypgia
oI/5JcsCACRHH++r+48IuGu2ZJ+/Ic6PYxZQIoLRggu/t6k1d/3qFEnjlc4Pw4hB
lOHw3GRXn/JM4HpSILAcuGn37NCo4ysmeQfRGRzyXNJGsVSHgpApW6Ay2Eu8ja2p
c0TgoZYDyD0V8qXaqgZf9m823SZj1toERB6GVdthPEQs1A9llfPkGD4REYJETvZi
+QEHe1Ohl478CILKv4qmLoEOAjC5S9h0HcKqgIrc8uEYp4snNykjCqZgmHylDkUL
JHs8gSk+/NKdCEWWz0W/ucVMzLLzPQoUzOiLhL3J+px1t4GyIGfCfTbS/XDbnRRV
BllPgRICt8n+jXaFyKGkCdVxMt0/VexkOiuaF/Kq+NB0pY2gg+UApLyQ2S6X+9LT
SVoknO6Hn8S9ArMsXZhWlAxqQI252cNySQlaawVfPqRwCSCYbQKiZm8th1U/LzxN
SxUmH5fdvR9goy+F3m9gPw0OuE7aOC73oKsWRgVz1MfKdlXdDXe71kAtKm4WBNbx
Yq4NIRllGV4u4cemggece6uqDlLmgvRnJx6Fr2czJQ/oSwUPqHlHn6TWJT2bkRRI
ltWMFkpaOKGDCAxqvNb+Hncw7i1iXIXC1kXik7qNuUzlHWEXOACWN3+JhN+QWzDu
LN/52Wn2k8Bu66vVWKp/3iGUL/tLKRbmLfuWpaHq6sgEYknYB6tmoY5ebr2mcwP6
VH+cUSk8DdJVlzIt0xwyTs+ccTewPcBXAvjvX0wJagzAXiWleowZuSZiHHnMs2A9
nfgmpSBv1mxS6Pa2rb2zLFzfVr6KmFBUaOHMWiR3R7TgNfZPQcgh2b+Jn/qMQhNi
5DWw5Pxf+tsd2XBGfajaNYx7E9PQbrzNtnMHBkvueUjxPljLGIe8Aa0p+BdKZhkw
vfbKWQNc3veSEyyF2xvq4w65+c2VZMw333IBQqt+iRrkZZA9hUemRVURvHiV5lSh
opUvlRqdC4awBzqYCVrNbSls1MyiST9mPgMwAWgc62b15wy8ajXEPrtvjXY3N+I3
GAfEmeSlhwT1CEaTM1YPzGFtb+bPCJkCNTFgSmi2jwkHMh0Fz6hthTunCis4Nzlv
MZ5Q3T+aGi4iPSWQWsV4ggQoo5/y5Ic5wjhwiw19jU+Wy7ZuGumCZbai4WN5t+ZJ
ysFgWaKvTq1eenl7GQ33L7eAjrl+E0/shC241wC1WkGA7MMRz6XFaunJvhvenCZH
B1ReO/Go6g25gWpUorTVjZH7l3IgwF+YCH+1l3KTzx9uN76HaWaCfJB8ebJgZdA+
EbUfaGTZsSuAr9sUoklunjtmH7HCkDZ9Tpm3Z9gwNs435YtQshmi3PzLweCObkPv
olXoM5o87csnWA8mrwQynVPka+j7/6JyKlbL2LnNfk4l57U8UkhL0gBELT4nc3ht
CrvvVHgp1Ub+oya7DB2eplLLDvK5FLanrMGV5QUnvIJpj80E1MZRUSWytQ5ZBNAb
gqr2djL4UQxx1cce6zEqzifFryHyAxggNeSAf0MKEYG6ldz0WH/Dp+3mfdgVAl8B
ZgxvooIjrZHTsMFEOeLH43SQhQnkCYAsPcXVglpr9RDhjmc0pYza2QzR0rL4J0QT
GPT0qwzUvj9fVlrYnfHAmUq6kPcz6Q1NL2jw5W9EHztW7vvwhyC7Th9oSl2q4RYT
Kg1SyUhE11W+UbS5jgx6YvJshNEiERHvJHLlqAahrZbRiErQaao7zPu849og+hgX
Z74h8nYU2LahRaTpSa7IWl9FpXNi+N5XoyIciNW3EQjDnfiNIQ00O9A36W3L6ZHf
NhTE/Mz1r/MWNoACwqfUZ999NKOFSCXqiliG76xpZeWkisoaVV6MJvv9p7hHgUK0
lT4Pes0wMKWiReDZI1Q98WADEj/2ann78RPcc5tkHj41PHTp4qJrwhPaMvzVuJ/h
1rLy6bkrvUFyImQNCrqHKOyH1D83yl1CY2UIhnv5wz8zPm3FdZJmvkgTFyKXgNXz
/jB5KXBwDZAvByLUHl5q8XvO7vH5fcum4x/RPwTyUmQ5xT9JRU3FKZo30pvpiZKU
ELclNUCp5645AxZPRnYSaWIUEOj07V4wBKO7UoBin0IHipJ6hTbFU5hAYokRAB94
hYKtxRrUlxOh27Sv16Atg6BEruFnW+Yg8rekyy3LDEnhwF+FA9tTxhttagVrB+KR
9vQ0vkh2D3zvMwN2ytUA1uqJwWnGJaEq7IkeO5F6OBnsB0HJ3TDXocJMnbZngf7J
6IRpXLAEICZf6razdae18OKomhjKat7TH5eGW/HmaNDd7lO6LLdtj5QlZ2D2RIH7
QchIkya3NFxQiPXr5NXFFPjWiXm/D060HZK8IOFJiDw0a0jRjGHGQ80R0N54AuLF
N0u0FY5toYUFRBRHIGOHDT11NfaIKz1sntHyARKZBZeXGEQjbiiZyoxcHk+WvMSp
9oBBBfrCZY8BQFiIU18AzIZh5jUIhdIVZ+o5J11IWiQacqNmpHuPH8Mj5cH1fm4d
JG/If0o4qDHYm51/AoD246P7bph4F/wdpDkh6mg8ti4+AA4rqrJLh+PXto9qWfZi
gFimO5xNEvBWdEUBuvtH9caQrLvpiEObxh3UDjsY7aiRUHxAlenyGYOofjAs1OdM
Kwf3QjL1gfOzqJgD6nTvn8wGNjHEa0acrQWEpCZtuzshpY/OUY1PfZt68O5jw7Db
HNmptMWSDez1urxdmtwyiIda0Ylucf4aKdQ5ha93WeZa8YtHtrByWzjscVNqz8OA
oWYI4Hd2gFlthUJc3tmQu1Ty/QzhjOObOqUSYarWf2likeowHvHEprfo7W9HyM1/
bI5DVcq0R3KdYQQpwHdqPwTDZJKQxfLsN9xyFaknP+N48hTfzi+mw5788jatVkmD
Ur3EpFUwTO1ifVGr9qekMlbuniF1ZpjeGmd2nErgl4BQRsX8aPgTq23131/yidKn
QnrK8+/xTP3fqDP/BhdD0G5U5WIz25uRNdXxJx7rjx7AaM21etmeqvBx+GWV+c1X
DUQScwVFTFoMUWXwGZPpkDsDjIJ4AZtM+lNX5xxUzhM5LnS26X9i9dywopj6HTSL
eYqE9yILp2zGSBJ4aExP5IfLBmwq+DJ2o/7gpk2tRf0Qt1lfHEC4nKXku2WATo2L
hge4L7WY49tQhvFIS2uDNnUXC/dM1nhu1rvpt6FOo8ZX+GpLQlwkmpLSl9Bmd+2x
lZTWLWXdEuEF0FGoIeM+mrO/TNyO/NO3i83J4PomrLppX7YbY6BT5DHT4SaORXUu
jYxssYWucjI6whIepsD8q40572ZvB+lgYKjl+DBEvx4eOdJNgvaeXhNFjGsP7KZF
AtaKogzxXNIgAn1HcKozqXiIvNa6dlVtItWcHZALsUq+o7pQCsNMBRZzPtz9ZaXM
pFUd19zK1PNQE1UC3RQn6GJm1q232tWHmVZpQKXAiFonGfko4jdtH2MWTztwQ5BT
QMhvIBf1ooBvf5sBAYl9LrNMMYWYoEemrtsT+4S+Ucvj7WKRL+3A2P9Zrazg/Maz
Ngql2v9c8yXlrpBKWgFQxwmAnctGk1txes4nA27yAIsklaq38lgNhOwS1TodJFzO
dSCSOkF7pYeoShOFVzWlszyFr9Cs1/MheKEQAqeQUOeEhIxJsoHBgsUoaf3AhUAn
TBnF2blQBU7TgCf8lBvJSE7ZfQFdhXm16J2rxveM1vv3El21tBTXJqFojdHYDJZg
+uJYRz68v92TV7BNyn1YUrMMVhuRevyGoFcubq1VGxEVFCvAL1xT7vmc7u88SKQd
I94Sn+svmB1NyyK+K6kscyPvzcPNUcn5wVRuJ2VpD37xhXB/CmFcyzyxq76sGJSD
epwgB2K1kGa8K4gok3QJOq0aJazyPFiVwaF/hhoVo7cvSXakFL5GLJkHUrospxoy
mNZQ6dynZzkntuCWSe1jv43nsaJriaucL/ea8zPekbTfYa70Q5lGp/ql3Ke9SRYp
4lem2xcOl/5M7uX8N6GYCHwt5AU7Flc2n77iaEPmr1/aznz6Oda50Ykb3hYtPMQ8
fnfsT5u6nJvG7JVTb6G3SIjdoFDLGar1fxSbgZlx1BQ77eozsYhV3nb7wyK1mg7W
WjXmgAH28c5PUkr0GBRcnuRdYuxr5ZtTfl8myXuw5I8qVjX53iY8wvOqEE6QSjk/
8XQbHF3YWBFO2KCMx6cWN/gsHDPIilI1hgNekvD8LXP2VckBLJT1kIyHPsCzEk+b
Dxu4I21ki4zOmedfoDTP5IWSq6A3DMRBZUd9FsEf1Fly1flYyL2FRw2m2mE5NlRv
KU2zlfhrzccgUqA/i++CBFTJnbNAuVE+hsREZfL8RCCfGtfZfqrdkleGvJQYwVGw
8L2SkFzF68SAP69pe90ixUOGLhVbKQuH8l+oJYlsonDUU81nrw38I3Mc5voJ7KpH
4609nshGA3wITlbjqMg2/vnvCCogV+moOnGTMPWlKIfo6Yc7nC/g3oZe6T9nyQlf
BFfpdBnajrR/xYp+jya1WFHDVU3EcZ8rxU70WDM6RXLqFb4hmQPh0y7lYmcy16kY
cCizqa2HEzLemWjDoPcnMFFsoYvqyFM4ZLwoTk24jwUECuEYDCrPjqW+WsbM9pvm
Rsyo0DTFC9CqnKlbCs7ykUdRyKjouarAjoxC8UXn0pVTblOz4/d5GiO8XG91hyqR
vJkU847hMUPu4GFqsIXcLM7TwgTm35eXW2YADg8yZosJliq7Pb4baO5fFlgG9Y9e
t/7BNjpSH2RWpdqVLA1PSTjn9uWvqWrGE4jH7q0fe56ovE3IZ/1IimFWsXS0fJpT
T1/3EqEmzYdSwd6piM60eO4Ag/Y1CwvwRx7J6e5A2XpmwMd0u10OBNqG988Ak8IA
d4Lq6U3FXhBC6ewQLxp2kO00K+YkK76TolXNFKhTmQKmq4ql8iP2lSVt6cY1dqs6
1X8998oyOFpK6h5JDTr8N2UxWrzRHePJ7YBvUUSI5/zM05imyJc2w7B0nyBshbZT
2wFdtCWAFw9B4scc7OX7hqsz4yOBkEFiZY1Tj0gYaltN3AoBX70za99obOwxvPGa
RuBEevkzS5GvAxUKiNXAiL4Mguu7xgaFcbNjdmvvKLTDSa4npXtrnWI/cpVwMSFN
9+VN+eIv4aly1NGHplZFEkZr+90MGCg/bfTxgNJdK7aV3FRAvMAIgKwVDg6nMAOS
9n/ZrI+JvTfF2D/HIwsPqH6pprFWk7RQo5Iaw4/+A5eE/IW8uHEd1cVc7Oh+r8ff
idD9tzx5I7jZl2UNs8EJfi2YMK5BUfUU72vf2jWNFX6lF+W5iiGPDHNWeFlcClLC
s2w5/XDHggOBgqvclKXG55399VP6nDn7Xc3HBkeAXvaJlvCA9b0jMRnsCmI9iXUv
c2YSumYs3Zj2xQxo22Sj73ygQqeY/JcdlUasP0PTn4hJENdjKdyIIHpWDrPhi+0G
JhysRtXzzjeaSE4HtIj5VYqgef0xYr0A2dSjQ8Mr64wUOTqLkkIpIiSRUB+CxtZD
vcP9nYsGJWZt3hF18YDyAfrAeA6ThnxDedk1I6u2qE0x4l3NE7ZLHoyBV8n59HM0
TOP1aeOhR2ObMCcbpqDNddOeWchGLDKboTnr0EGT22pYhL72ujjkUqKcBHhd7Zb6
H1xj4okrGBjo8Fn7jBouYmXVrAEtA/TF7MfbSeT2JF0zaVv1lLQPuBXU1qsXqIIN
5q1GN76ENmWS/VeCO67Wd7ClUPvCliZKmYOk0Cl4bS9AaMkwieLGfh0cFZHcEG/F
tmuDAA2VZWgCLvQWeIoWHj9nk7inTfFyW9+YxG4+e8qY5afs32pux6NBvteDvTxJ
NJ3SljSjgxLwnCtqgk6pXtCjGmNKZSyX0KcfGzIYc1NQyj1k+4sl0PnJ5aLdyLC2
T0PDuoxQz3UH+fOgB+DfhqwYCt+ZvUIlXBARA0PN4fmHWhE6AEO3kEYKPTuoxedf
GnmhoWkW0wYl+as/Xz46MhvKerpNiGMdNsC1JSRfmNt9maliavWubRb8p0N4Lqy6
PW8Sj82ZiSinjQdl7RUnj8OsfS0GtcjMUjy4Wnk0cZZEc+cAcGm2wOqliMp++TXS
zRC91MJbBDcqUW8nEVGZNfHjWCWcPSVUackmryZ7nJF5c11CV032OkYltbK8Udlf
gXFjAKguk7pwh1YHg/flFgXeEYrZsvJz8Eyelg62Q6YMLBGpdKRuZKHx5FvjKGT5
11ErUjWZ+CVi+uFiJsA1Z2Dq5HyfJVqVjutfhV+HUwFcQXU6O2JDLxXIZhPmHT1q
BeVjN8eAkHBnw1XQrIx0FEFZMtztjN4aDIaVzhVu7zOp5FKUoz85pCigTdfP23d/
vKGfTvBmnPEua6xcIueMBZftIQvaTg22tY/76cASx/EPHIc3r291dOB24ZsmKNJN
qTlSRWnt4Gg1a9K5tsou9OPpX8KD17Ix1Vsv6u9dOV1T8Pk9D6gG2al+65SZ0isj
Q9PM0qnSFb6yZGQEtBLGHkPBQS+uahrEkoRgopmBznQYFojfBYlKuHArF3SN+bs4
uJtFY1QqbW22qQDV/2nvQPitUB4s2M9vjCgZCyCV1NEcLKimG2AuSv2zR9ilswzQ
DCtc9JJoH1YxjCugTrQ1XMnos2FYPWXiBz/BFjy/jiTkVPP36FYf+VobNk04I9hh
SQtWUFeGGhxbFoyD2KDkAjhHgfuQSst7LOCyg1H77WXdlCSA16yKlz/AFirxrRI3
o5xP38XS/WI2dWYl8yf1z9x4N/WUEL3wCSti4GF+xUpE7A84FTlerfs5AdsMwKvf
DZQ8MrJwILcaUI4AatAIDCS/1OAR+4gSuVUPUL0X4EgFA2wPU8YKCZqXJgIqnmBw
QfDoVLBs2k63RIVhFhGC2zF2VR9wYR2xYnerScPYunIk5kGdPVbItGjFxJXVjfH4
GuT+Pgt/xRXqP8Zpj0fimJrjgIxJFpAwoXiBj3AlGlya+Kushjp4UTGw8ruW1Abp
OICxcjLeb2oV4aJXX21WI0BsDaevq5iTT729LSWDflmXggUSqj7evJTsP5O5DSu5
asNTaKq3Xd+2siJdQfhxubOcq6SRPSswnib7Er0V6XhhAbSth1S2BAyNidyEiwX0
uXuBZK+8c49KS8yvjNNDwxY3e0C+kMe9kXWTI9TVqdhsvS4bYXxU6m5H7OjDsYN8
1J5dG2fEFJuDybEpqrCSoKhyX/X7FS6wdHgLRdmhGuEQ44ZbvdCtSanYRBA3pE0Y
6/rFJ6vY5ry9WFXeFChtwjX5HZtyAVTQeLt6imbzsmZLTc7haEdO2Q3AOxUUJbfu
T6DGuuGCyGPhPZrOZfvhWCkxqFUnkArT/Lxwzt04ggAjgwvrA6Tr921kuMzaY8BY
eErZXlHBw1XrSCp0MZ708Pl5qJfO9aXZfgkqIOy2oLtEJgyi2WO4lV5F6ip0dK34
vJIs5zd/UgzPDQb2WKx2CgRRgyMHQ4lQ3EcXLwp2hEPxUPHbl3kk4TAiWwjbmIZ2
9iVt9JOTHhx0S/nBmxPJOR1raiqVEm54qh1FmznNgjkEbTNWfF4bQaxBxZTQiyTO
SGF5gLMmHK835CS77mT3ypdMXBHcHvMetCQHdncCSZsCKKBsQEFY5o0t8m6Sj2SI
AmKeXrUfVtkj7iCkxeVTNWEjKQE6pTrwHXTc5F0/6v8ehwBEaJcCTDTIIOdjLzOA
Fd+KgL4PH6SZHZFgEdewheRyY/QUA18LHP0dFEK9l/b55Q2A/nARfMxfJQdpMG8W
hXgdJuaGG5PwIAu9DRohkENYTj9ut9F19rgWYsFtmNQ9baa6kDynKuaCOHQsjKZe
Q+p4WHF8ygoPhUp9IOVNKl4qZ2bC4nwWY9DEJ8hpJD5+MzhgSFygZlypZmMiJlKd
1sQlvLbiP/61x+v+6R9J3PctbvPXMlS0cveB4uwVopOR7r63besnIIWhED1UUNbE
P3qFup7A0xI6v54m95CsV7a/rFQZMjmxJl10wCi1jfTkDT3aUHVwsL3kKd7WxcOZ
jui6Mb67p8WvUtV5lPCvQZd0wnNQpEadVYofcxvd5LxKGf0fIC3AynEyPCWBFONZ
oswWYyfkO6+ApPFHCZAQu08AcCkaVm2gvcHlAPVR9/7/hyzhvT7LrTBfGI5FWFl/
qEwosUcozJ9xaPEuJrKKBn8u9OLFCfxusJUyIYRrhjT9gCBcSEuBrGSEXvbud+G1
7ji2c5S8xPZVKVqZyP1oF+cdgiQe/2XOg3PFwKgoAYWImKPJrM/izXv6aKurQlRC
SeYEgAkR/fNUUfB7WhMOmAP/T4ZilkUTGqfJaB8yVCxFFuBSC9MyzshvyliIvDIe
pB1P5wTOurddJ3Gd2PAvZdBB2eUawJ0xxZ6dVrQ9CwULQ+kuJwTtXZk8w9VxyP91
NOSl4wvtJK3sjMljJtnY6l2apNVaRR76DNb0iHVL+DLkvb6riIneubxcguEDTZlZ
UzaiWNNt+fE4Orid5IhVzQ8HHCOmmsIqLKa86nR7eRV4Zko2hABbGj+cZ5F/1fC4
x45QSdlgwK5QGbt6Snz40ryyEe78PqQauEx36SigBUdh80Q6b3QJum9lgcge3lzh
D/XViHWQugGSTCo7wfzn9aI1q+P8+yLxTrnPoSyxRX6IsiZO39T14xpOEAFlxnIV
R5pTw/M76Plqp4O/mXyJ44iv8eeRpo3KM6v9zTarZTdTBTTqWHHZmahQaMrhRM+4
eG9Pq4kQrd3U63nCVT5m+DQiB7YPJXE3qokiMGzID1yYbTNrGh3J9icm6kVOUpOB
WBYspeERBRVJ0q0+UxTTvACn2nRC9Tz6g2Lkfwv8/Lp4pzgGD7YvM9sYRIJZ+2wX
t7pocmOCqOYoHG8PaMxDChCGioQ2Gwin6Ph41jBXbh6LuYYj25oEnvob/Eci0MTg
Tx6FvqI+Lm+bkiFVXFzpbhHu6paUgJSg799QdIOl37Iugzf2Bd+9g3nzGar1T6/f
5iynGKO+ldhWZRTsM9sraM+PAofsIhrHdBCmXSRyH7FgmMwpcpjH///gKi/n6QPn
DFfBqUr0cvtx7f99rOA/hNf6gXsDfQGH6aV7mzGVPx9hckxkI56XuNS3fFWIsrHy
6JnEzkBMLnZTRtCFHpM+VYwT77f3lXGn0VlQZq9Q6c6IV8aCRUhtB8XwD7huP0d3
vaNWxD/TPpkI1ERngqiDvJOZIy3Gg5YTYichh7nF+SuHMFDiya2f1g0TeWGkZvkH
SU2tJgJcsHFD/RVIzTcWNJzOsaOr+cWHJIMpT1AkRrCtOj/zWaQmF5l+2Kj0tyCC
aann08cz6kk4OP8PfHpHKU2yka+4Q3Ua4RP7aTpqRmVYGWpCwwlLm7HrXePQZ9Cq
2tFQddvWKg/yjZrcAiWBcp69goP4ENKZZEmtLN62zadNCP25GuG1x+DOsO46ReG9
02aewsx75T/jOCj4AQdrSnK73HE2NmXIx/TKZsyurCfRt9mdJpLkbA9Jyu2vrSxH
EdVw4EaEbmnyfBY8wqGlXaLDIN+Do5ib2+Zl0bSoJ3LFSGCwca4BuCqW08zQBGRa
sAq/vf9gtqk/5k+eEXo4Yy1guqdqA+BHQxtkE3lE5mPiqvvDd1g0brCM3z/mtepX
aKAuKwTjIl+99E3i4I90vTU9rvXrM4Uvpa714lzPIgRDKvmrrEJS1XaLq/rhMWKE
3Kf+x2fs3FF4ucKbKMWPbGSTo4MDLkSWC3o33gDPDxSnuyfr1YtEk2uk6C2l5TaX
nbPV6An0eKnF33RFFRxVkJ86Tgt56rbmoZ+VHFxByvRVojztKNX7QHQ7t0/u9K14
b+LV0EWs35m6ZW+bQ6Q34EfLbZAFNPtrBufxa7/ulp7yHBM2abJBMIloRYFiLp+f
g37PRmGVHBcmV1igF0viS1zDW3cOEkEd/sog3Ze8DkgxkJQl4iV8ow459sihcvd9
p/0nkKDWSkBPy4SOKklM8XXOPOuyedveTG+BzrxXzfoKly3pd9TsQrufb5Z0OVX4
J6M86k2TigkmyNScFumdgGrNxh6r507h++BFBUF1JqCAYxZxpoqQIPArd87ZU9vL
EetlzGjIpBY2qj+UI/AXqL2M/05C5MP5lPEesn58UYbcuQB4cyIVOrKDVr9KCJfy
0QioMy9PVp7XCrX1VoNqIioREBkeT7UTRS5H3jXTU5HJKaLCAuzcdxuLnORgqF6+
iDitr1yH4FdVa+/Fu6vWeblWCBrxwGPNF56eJW6c/hyHiuyax3TS07Nmlj9GHq0m
avlanyJdMnvqJ7DaXYUOzyUS9MATjOgQNTd+D7gn36OmtfRUas0AFoEb4ZGudmMz
RXYfEYwZvGz81BVRSHnT06iJ2kfwvPFZi3Pmt9KM7CAOkGMyLL6nPhgaNNCR+B6F
XB0+x1mmQAFAF2T4reZTnqOHp4MUE3i5IEJN/5UZkffxR4faMsG7ADADtxVyIlA+
801RkHXMzr2pt2DfPOXNga52lT0cWrqoo7J+WUJnzQ+6zr8I7a6FNx3aYuqd7Wjj
TCytqUv/pi1YV/s6yOeSR4fFHOj1d/7dt13spN1l8r/lSCG2uFpsU/1JDGvj8ZuN
0EpYQ9NDfnJXHM85fy43djSibO0x/XfqnKhRg7RzJh4akuEfI8PY9j1+MaT7iuZW
TuvltwRCj1NnzlUs3DpKLlOC1Y4Glf/as8B0Z74hYmMosc2HPWJWMIJ/OoSqZxAo
wXfLCXOKpJ/5uYCGdMKlz20kX8s0ryqxYbQ3lvgQ9QNR5LMe9YELTTzvamiCAMmR
Cql0oFNp/KpW6n3PLrS63J9KngcaEUCKdvHWNdrI2a74F2UU9uSjumVVkke0FQGX
b6/tdHrRCpCZ0i4FARLieo3x4GI/KNlkJaLfAWWRaxTMzbnfUn/K2SuqQBHP5eQr
U6Phv21pooortaAHdvFoIUTMgzMOwPkhsyh0siKWplZOSSKJd2tJoLd+dBeoz3D/
VQw2IwAIrauy99St/9QMRNM9oVO9zdxGPjTIxDAtgEgdMSGBb6kkxXOE9XbSgz0E
yB6qy7pR9G2Osv9EXenUxjceFkPU1OsNft1TAlctNAtuyEuAx1Lqqe+JXHG/5Eff
QizbSouPZ75lYlu3OB7e8hUcCNEsuJV9VQrAwk5fZl9lO5bLAs2iIajwKu7PFNFH
mFhrumfE6T9cPRTq4qsoxuCKSuW5VTJMBkNOfefSds22NfrMNcDbvdgrrwudoki8
RGq2zsLaZCDVgc8DtQigNFyHpxkqmS7reBMA4OIOkTDC5xTish6hjtvzfB4jZQGl
E4YD7IEdDBY/eXIyA98nfhWb430wPiwdSTAhlF0p4TCuB7Sd/u7TaoQaKOqQFEZn
APACPGZ2Y/HJoY3tP3WVNgVFPSIAHLWnD8HkV3RfYsD5G0GdYOKw++3mdfAl2uLz
HU7IAsTAYIn+mmV0qcdHw4q3RQOWv6R+S9breDSm4JUnRlsezAzDRCCYxMxJhJvr
P5KxKAbil4TM4PIujdl8NJEs0Ry9eDs2nN5NFv7A+sEOQFj8qhSaSjhXH4FvVRU5
L5vEJ9TpfoEOS/sp47B4EiTKAsHTU3ois5OQf0Qk2NnzxrgKvCB2Twr7ryRa/kWa
SwPs6AQG1Xj1/3a4kgj4PcuHHimyLKZaExbWmPLGoeWd7x6F2pk7EY9mBo+cwZGA
oHaKstZxcT893EeKcoCpCPHZUEw/3n+4Fw2vgJ7rpC1sjN0/jPS0eNNNZsDi2DsG
KMv2UpDCwa0Dqq8M51QJXUSxhfaodkr7l0Etpm5yQkLjGQY8QtNlAf1ZhO+ycyj+
cbIt7piR7TSs3qv2xdMYYEK91/Lq8L5/3bY5UzA+309GuvdrHbhF2+BjtC9hixww
PoITdlzKbF3qH6+5/sPr8gSk20Qip6oji55KfbdtNwtHDnVgROb5KBZ7R46MENNE
rZCJkZkWoVoEAuG0skQbMQb4IAbpC9kqpJ1s/MdvmRhM0URB+M1VJBnmMa7uQfCb
XP8BIEX+xPjZR7nEQM3o6CyWCbXl5+iCLhj5mPofZ8STFnSnLFrSITT8eet1YTKC
nstKb1TJCllltz6vXSoVcuvbU3zxX9SirmNqUm9Y6dK0iaV4PSVq9lGrg0myIwBA
aBdlYYhxmIWK+dlLUgiQgzCAnr5TEvyXf2VWB/MgGUIRF0OZHTv5rp0qOuUyu4Uh
nssMxbnMhd3KkF8IO94yxflBLj/3YCI07lkCcl7NrB+9utcKWH8rn6KfBiunW5Ap
IBHf0Dn+C77YF++fJHZgLKcotXzrqWEquj2M+jbONt+jZcT5UcGkTLncylSxRGN/
Ch2Lzg/kb8gbT1AnJ/z2MKO+SAROgSn6ZjSXEIru8I+Jw9cYEocaTy6ynxZByd+q
Iy+wPSfTg33iTxvny/gEIW4Rak2MMBMuT3ykeTx6wGRRUJaRIMHg2akJUMayphW2
FSHkIGrXNy1oNpcbf30/i1nXkzhYzFIjRQJ0wf+HkBrvp76Rr72RUZRszwwtXn21
7evqgHOO7lesV1dYk2sKQtcC4AGABKaHIcfh/6DSoROT8ID6WRAnIAFaJrTyQ2W0
SStAHzc2OI7mgaIRK4NNG9W+T1swXCCKAcx5rd2NZogeZ+9oEWm9Os4yZSE/Sb/+
VOw/qE2McseovKxOZWZXqjaZx/ezyLSgAg7deaXJfh+oqG+kEhBlY64zlkYNRIAs
jf2iUE8DW4SXKayZrwV5x8IZVp3ZUOxYqGIBujd/zwnD++usTpKpETd/9Q4ERDZK
b3MDJp2a6mWnEe8irKed0rvw6Xx3dUYnaxjn+F80ByeNtyhyK0k+at0IoMBmIJg5
ZcDJ645GUKWVF1WOJ35ZOOzpjEt3+jrixORHi+Si9S+s/FUIZl7K5u7Bk3s6Al94
vLknFs+spxRenHRSG3g06yUznHi5IS7Fx/nJUoklBJgQWppOduirQMEdhy5f7TPx
G1t1uKlUg2lT4UX8uEpTtwxDciEZQCxz0/wjXZO8nYDCBejnf7THGmiDCvQdCdKo
xuvy/D2cGF3Ddc6EXXMjJ1wmIYJkTqj4L93Q6pcTu147fJs+ve3dDSIH7VAlV1Ab
gFxZrQVJVks7v+6zYmoingOBKClzT5XjArCotUnnTQBC029ChQpqoEPqWqT9yJkN
EXf18N2PY6yJ/841n3FTd4nz9zexv31t9ICM2CjNuz+GB32MxdQZrxDCUYXJxdPl
mNxDzPYIeV9DwwUHeL+NdPhgepchCsOKXunnxbaGozDX7hX+4gvqCWFz+MOPHCiZ
v0n9/2amoWEaWfbMQE4kAvCeoka/ULBdl2Ok3kulLQFaE8ujJVqPoBj6ELR5H23V
UVeIoV8GxRyr6PH2XxqZP/sRRThZ+zNq1y7d4wLbpZHAJdCRy/4hDclAKrW7BS+h
bRwKxq6LxWCzjzPbSZu3EBhQTHHWqVx3O+gJBG8rmB7HjwrQ5KeqU/ZwH/7/C4PU
BDQ3OmmI2c4qty7Oe26xnIbvkjmSOgmrEosvhcH9f9f3DU09oa0cwGB9DvKDezwt
+9HDupqkWQkM8O6pTrjCoHSgueYsXHAR8BoZRRKIVbNfP9Sn2RmQ+Tp4ztxkeU6B
z6FtfZmy92FnyPUVJUFDVQSg8eljH1qXIwX1wuWSM3rK2X79kh66ELkM5j7JcF3t
nJSTtQLqFX4wz1zhDWL1nStyBE2eqJ4R81NmhCXMdF5vGyk7DOSpJ9h43wveGb7a
6O6A/hCdr/yexj3ilBpsGXIcYEEr3W0XnjtpKXc1CmjKPzV729TD3Jtuh7cTBp1h
vgjDxrXIgoc4n6OR8dJ6vBrt+UvPxG1gHwgtO6Sca2MKSW5Uc8ZY4NtKZszxqBgs
bTfA9rk0Ni+GZZx23az4SOQ8yTdq7pYFvIkyh2yZ+Cn2LxVQNhXT3pTkfBSYW07H
k7UFWPC2i40mUlU5kWJe7zBHZ89v9WZhdmoWvGkAQ18yiYJMQQI6qmcZqQqxKHB5
35ueHQd3rnNNh00RgoEmhRg42YalUi11F8m2ksqAVh0XfKj3L+6QbaeDNQoJxqUb
NJTiZTGEl8pKHOTLKnCpYQePlHo/vPAFnINMJPOonpbPbZiOVclh2xDQUDCLxIyd
aoaa1uoNDZF5BJOPcT72nV5pL2EKjmk2M2qFWUjZu1w9kNgfEawDktn51MNdLbFO
yF9NLZ/VRpeEE1LjRgz7T6iMFKECWU52ZSMOgn+MrQpRxeRl7noF9mJFlYcgUS0f
MolahnCE3DxSfHNj22TcuYFEbwWHvCInxU+ZoHy2eMI3GEafEtST1v1Z2gml8kQ/
DcyYk9n3vZLd8GltqGnJ0icGFnL+Lr0d9aoSGT3jpB+H7n8CFJ9TG3TXGkno+Oti
ysF1JkxB/Wx0f8NyaXsN5ez8VlcWExoZXBu7SpXPVlPDEHHuuLuY/edXDcma1Tgt
SJQIBA+W6Yoc5s41DdTTVzO4f1aIu8qyqkrgaFrM0r7MrMsR6CGCkEm4PiExVcP8
YVsYh6HD+gXgGryUFsM+TYNRhME0dTURZOgj4As2xP07tw7qguNpuyOt6ZCwEzUX
ya5LStPw5ECQYb7t4wnuLKwnVvDrWsjJMU1r73XQsccwOAulU/gAmS0CfXXKS1sF
hRuKRuRlXL7lYbqQ73BGRITQ+cZBzfkp9YGWIgwwSiruSst2xY23p6tIVWhX46Zz
bIXS/3sd688hzXQH4nghbqGsZIpJOkWLp7d7rskbuX/sk8DH6anJF0tmvACV1MAN
2CFf/MtTIMt9rgUZfvlzVPdAwU8ifQ58bUm767zXqVfw093/UnvfVX8mjk1i2Out
5tpXHc3xChogWRZJ7zAoJGABb88fQnHuwc7epK/IGvWX05KVwbR74mYJ/pN3lTjQ
e2OKL0LuGEhFe3r/DtC7AUH5PhwWsFeIVxrwQyhd1RR8CnPGbr6zhqVmzTEVsI91
YMSqfoP3ixuRBjuvHDnTiox0jN4YaaAKGxGcT8znvYtz7hmSksiUinDdMdt2txmy
FzeNwbIkAqDGlxqvDQW8Fii3D0iLfjYstL7vq7OD/YmxG2qJGmcpSFJA3+0rae5t
82aMPdq0Rnuow/dAZrFBtrWyPzK0Sixf+RB1Zhy1fCytWne15/y3kl5gFtzIUuE0
lCWEGIGE5MUf8cOg2CAyrX1EjWfTDILrJLDoAJx7k4hj2XnbxQuZs8/voGbqnN04
J7pPmdYL1nkApqRFQ3mjfms/P4kf0uACOuhXnkoaHMR7g7HRvRYUzneLls6Cjn5f
7Ml31UUNpSERrETwt7anQGCPDCijH+uj+itNS0Y8pZhGYl2D/SCINaUI70Ul1wSt
MN8ORQD2/lZh8q0QzCLEmoc+8eTUkHa36/AQzS8ujjHu2Ig1Q4BZfK0XMmcjquBh
9se49moxhaaKMxzeY1SA6ltSqWHDFcJ2LM674kP8N3mzmOxLk+2GzGjeiBFZ1xd1
hngkyB7ibv5C5yxpQpEaVuNx1fQcNyJU0Y4wJ0AY334Iwwgc61ARZbZWAyIHQdaz
3pK1wD6VrKJDR7psp6h1wp6eVuJ4iQFuZzGRSLygl92AyZ7P03ag8B/cyFrWTvFA
Mp4v+SHWgQAZbhZW37G/UiiP2yN20LniJNZcC7NQPVxPNKbrasPMnYvshtmDjhIO
r8/2pYajRPU00IoNifIGoVpltKBk+vQ6x6KBTZcPzjSVh82MoPnA3pheB8j5dyqU
2c4rFH5u6T3cnKk+23wncoZiPctePzGaEzxu7karEEorWBJ3JIwdOm2wt+OWKaoe
Me80GTEFCm6emJRhgYtequP6N+HkoSIXSRv/atLTMtvYUNx5ALEPK194aN22esc1
WYOiNh2bnK6imLqaGtg0f83J5wyc5/fujJT5gGxLB1NcSWiWiC8eVfnJAsXQGm5I
TM+WKDG0wZsB5hTGF58e40DEZMLTuxPFwaKZOYHPCZzaUcoGKfCJzEWcjtfClsrT
kfxl2JkwHfwF27rPCvWA8FBcfGMxix/2KvYrURfwb//mP/c56iT2oEJPkeYT+1eK
5zpKnZWmO41FlbZ7UTYC9au7xoDcQjzEXFmcueFF9dFvBH2u3bvxirCqw2ocsTMA
VFOjoPIcgz1YjP++oeidodi+mMiNCXUK1uwRiHaxEt3eTS46i3HEcCVecLfocs2E
Kh6OJFBPj4+BwkHD1wsvckEcfGv5TQlXQlPcokLb+ScY5fBhzag+Y0caVvZX2PWM
yR54Xta7iJ9p0bthMLv+nox3srJCypYrT5gYehDrMbUV4RFwufFGPBQcXUFQp1LC
9zRS6W5YIzEaPOb16KF8s3dNVLpgwzJXGTgK5+vx0P9Gp60AYjxckglveegdw3vF
lfJeUFefYGK5qlWvgRT06CCXo3JcGeWx954hOEWEC/BWd/EaGqhkBY+3XH+ey7SD
xqHD8hKN2kz3VAP3m2YqCKonFVMQbErEZcqVnZ0p57mfg0eQzhk53znxfiu7FcCZ
5hiGi7nDPFobYlAMtDVIAtXVKVV7M+Xe/Vz4JRN7xogQb7XAw+4grW9MhDXK0khO
+fhUfnydpNLqMAZLC5X0Yt0Rtn8K3wl5B1SyxTXDT1qAPuasWEKdALA+j71Fpca8
+AJkULI1dk19ebeUGjvaf0F19rDB2FTlLZvz0+/6RngyX9Psb3UaN76ZUeLrStiy
/ALJQj92odvBeqfERQVMX4vfAr7u83mUhjbsQarCiW14r5992qwum3RKYPAKehKR
P7aimWqCG/9Kqnsu+oAAh2MX7Fq1Z08mYW/AEeCzj/52J/EI2Iwc0Tqd3UAgI5Bj
pBOA+TkoYhjsyWPmEN2lAUxRntGkUU+XRXroLjD6S9Vs5G8a6bUisnbP9H2OXt8j
JypxKQyt9Z5bKrsptPGkKFBorXjCm/cYeUC+k+ICDNMwS9Sh06svL2CqDh3ChgzK
H9XDEy2j1KbtM4Bvhzpw5gTZkO2G2O18E02uCxcK1q0ep/B8CrC4+WHB6ZHK2T1V
5SL4e+15LlNd3BLvnCEMOnDkFsJU1JD2QhWDcmfenfdk9WngDFJYj9E6gKUExznx
gKoCLUisqIQuD/MCTW4r4AwzPUFZnUKjmf0vCXdoByYB0VW+ySV0WCLiTCfu7YJ+
ENO/C+18AbA3dqqukKmBDERdAP/BQpdD2wbKrYVLxzJ6H9W8d+HnYI9ZlaI6kY3w
BkPS889oPtAmeCEhbBqPnHwiZ+JWvF60t3eDYHXfyH3vkQLGLhSsfML2j9npV/0d
6kDYAiyuFwNzixqq5Z1tUmTUBFi1d3IWvaE4XMPsOrxSNkjKwUV8ABm0eOQF0JPb
S9a3voLtRSrZNWTkWrmzHZMLgkU6y0Nsor08Ok3QEK9QmFhSnFZe8n0vYDkD/dEF
zBQN/8AayFXHr2HXgcBKAVgVIdkaYDP2zDwaghg1CYYogMGDtkettv+kMXveKI4Z
7hqQjyFQN9dz/mLaAeX6my8yjpX8Z0PfGxBsOiMK4rOwH8rFm4tCofywUI6H9tg4
Ef0w2BhswRgOuW1itBpG1F83Bw6j9+MPejtqNHXTZyDdYK65JfNhAFrGns+N7SeT
hM0X52Y9iqu3rUHYbUJpBE54IVM/dcFtBf+AZpHD5I39w67RbL/NdDo7TnDLLZwD
9tiln5vY4NGorl+C7v18/q7Xx5Zhro7j7rJeRefpv0BPgCkF30VnR+jjbUsqmM3r
MScJBESpgqtM8831peA6efWS+l2XsXPmWTvzkyCVFgQFw10HagGdpVGERWKq8gC/
wxsvwgzh8N9cYtw8ECTnzsXrTBohKtQulPBk+4cAT4q5QWXQMTyf0GZ98WjH/e7c
qL27ak8LXaxeqG/lllbV7aCThQTHOrSpue5lfZ8FwibX3QowLy9keQcgrgpVnp4Q
Lyc8qsAqSBsbEETkhF3wL+klo/4xrmiJcqy71DN1cZ5oqIzmEv98rExB/RXU07Kx
dg2YvzXFTd6MmSybSYKz9100sqlNDWCJYSri+pfYoTl25FIwC9NioYYG+3GXD8es
TTbuWVOK8DyLHx6RJzle/cXxxT+sLrGtEBHErgxqI2JcEFUv/KWKPTpXSf84mLSj
jso5buGF6LKT/iAZvcdNJ8HZQ3MP0lTrnJU1CdFa2F4YW+/VPzBF3G+wUathCQ1x
vMDgU4309aohWTqfO6NS4zALmW05yS7NHVNM2RQj3UITTP1NbRt2Jq2O+luB+oOp
AyfqlK4KbEe+k4qI+Tm1M1iUP7p/kkNY64rQsBKFZb9N3TC/+xVUv2oRVeXNeqOr
+Vs3XH8m4+1UpK3V74nRu0w3UVgMPi9YdCVtaR3UX3HahmG76SLSw9LaRxnVM6NR
mcpGjkG2adYfmgT4skKFrBF8nFyqhSiXqMrH+f+2pIOa+z6GkOoiYtsI0X4DyOh1
O72AjaFkBD5Mz01UZhnEqdBKoXPldTYCU0+bk8cGf5Np2/zC+wFrooc86xKhbsze
v2xbXyB9G2MGWANaavOojuC2NToxXWmHfyybeMeRRgB3td6iOC9tKyrJjtiX/hf+
euIGNarVy5f94rtXAmvjOfa082+523R+SZsdEcf4WR5bxAb2U6JovtIeJLuwhThI
eo1Jo8TBXXfbRUwi6LpYy5unvDOVbUhovH2dLWXwYSFbTh4irDZddwPXs4JFNTsy
TLqZuRktPg8oWCWsUObNiSTyqJdGvG6HEx1Bl2B1OmPiGF1aYDrQRFJfSWmkoMoM
vcAbdatumqra1JFHmUKkhtqnTz7PUnDQwN5AlRpk2XGDWag8jo4RN+jtFUTXUZCB
wT5hUqG0Bb8bNoXz4rDkNVYGcD7UcYcCwnxR4CuBz2dRtDRbeTdRS4gOSeTJiw13
DJi+BSv5Qowwe6HEmyifp/QGcAspf1WdmqeL7rbhG6zZSAQdUqSdrjviGtlpjT1H
+Wl/mtUukT4s3+KiBgXZn71Z81uvJUwT6x7cXskjgiBmrQO1OLY/o5HA/KnPfQt5
kT+FnMDQ5eIGVvXrDvcI2pQX5zeZqR3cY6BxnhttuHYxn+ztQVya4d1PPzTm74O7
ZpHYCeTLQXVPDf1pQYdc4LMFa5p6c+Cu72/0zHordmtjR4fLS8F7I0lZBMuqqcG/
odMpNT3tTnBsAqZdKJHSXHYGs82fqNkt4Q80YnxwDf8rGLOnryiptW/oDPWP8pR3
kC74v85ICdfTBc3J3bpHNKrNpm7TfoSYaJJOsVRs+MdvcciPbBb0wOcQTrK79SPR
Xc8LmJUuarN07crE2vnDkew4Ceek9kNUf1+ZPSDTqTnrn42L6g0uzQTWgAwRnM++
V5/8XDayzC3AlXKLGNaW4k/Y1s2BszCxqBaQrb5gSgaz9gshgB4hJmlqLINXINCA
fYSxWhIJqibX1Ik3wSTQK27ZYRxF1D1AkBo7dkKohBzadch3fIF5DUCo01gU/xG6
/L93QjeBSXEEKBwWobVlc0Hmr4A0aq++wD1S5GqRuweJeBOda9q7yfO6jDK0lE7r
cOw8NJGWkaTus0wdfIPBbl9EgTtOnGt21GIqr/ne/ySsfbfp369lXkZ7uHaotmLh
CXU19SUoOA/Sc8fmOS7aLcAKoIAO3360Zu8LcCfhVzX3lLPoB8I+uUBL2Sc8BnVK
Llkjqr1nBuVhvg7f1kcn6aNkFaUcsSIuTzzUWBPBQbPCHD9fI1CnMjZRaX39EtHZ
K713PEnnxnYskmyewFb7/gCmn2w9W7PRRXyMz0+ENbxyO5c4hsIdPMrSeii6yYEF
9QbYZqhr13wvAaLswAsLaiGw3RNHFjG7qB5ZmRUlH8HcTb2EiqyFi/mZfaYeWQ1w
aMUJaaAqvnu7zY0pGoGaOJ9xXZVHF8xHaIikqjkk7hHtTVpWuOcrCJpOfoz4thoT
GjRxQDlEZXBl+6j8PhGw1cUfIEG1XcYhQxBACJOcfG7UnWFrNuAReE9NS7oga3ha
Oeejq9/pXiRMYovkEbb0tLiE5grHS4WfP0kNJYZw/JQA22ZcCDYUyb5A1AzJ4gn2
iXRMkYw09bDlX4KnJ38RJMl1cfDOVJmY4M9jG318mODdENuwa7ueV8XU6W8/YI1z
EqlG44vGAX+Q4x/ggAxQghdDdjmurVCyEqmcSsCntoof1rLbR2bnoMPv9vXZjKKB
JI5f2P3WyNkQHYlmq7HbLAaHqPHiPuDyM1Fr8/5rNZW7LA9B29+J80BBUyHhFIvZ
P+ikKBQUYw8C4M4JZeDaBoIarXoJ9vB8CHxK8uIDWgYNU/89hIUJQegTRgcOn60n
3ZaiSfq+5OWS4ZY1dUEFMS5P+SM9AKEPZH1C3AJPj9dtxFh6m2Plb78kEvdLyu66
Uiv3X7d0j4wBS/VlaqN81020b7mY20Kgdyk3AXTcNeXwb3YmsquGUcV9qCiY57bg
uIB7NIX4yu2KWE9P0q1o+HjH/kGHJSHmA6O/pBzqvFcvbz6wTdxksi7nIbQOnG82
Vu3BfawS3FE3a7ItNKQdYAFAg5ct0MIsW128jiZLpycPOXpgdrQpKKfr3AE3IayE
HcRL5juQcKb0AM6Kh3BPC8Pxz4La1yuy1JYxDhcTqFva7BuDlHLv+Wj0ui40V/CY
NPAwyTiGDIAHpxzVoRO3K03UvhxXuyCQLCoBb7D77xgweUW37Rcw5uNHcCVE2Q0H
GmE6ajN11aBnwPFzjhu3LC0ug/xprq36K4t+vLH74yjpwSN5VqmFnYtPlYkSSEIw
13c6mLGJDlbMeLJJ2/Jbst83AAe/A1I8mAcNVODxKx7eMDgUqlASFLPxIBHqZ0n5
m1QlLFbFQeMzJLQxB+ag/DyNqoHyE2WESSqANFPAxK8sDzeZere6NSFK9tmjNcny
Ms4X2PagdfAKIXqBNoDx7Pc4S6Ik/dK/CYFEuUQlHfiZyPhb2gudbRTuZuLQ0+5K
8eeyLWsgQqkmChcXfN7ZQtfwHL+cVpWsrF4CWqI4mIU1PJvguN+rr4e/KRux8NpM
ZjtealxpSCb3vgluyS5XpHQtDWdMNrRicItRWJjmrXCY4OycJPNNTNjt9phnfUBK
+E6PVs+1Ypt+6DRXnPEyYXpiTxdXBJtSyV6Xk2oza13cPTKwDsVj+n+XgAgFbFAI
4ILeV3JgoNy/MlwLOjfmBP+vi2kR41u9FT0ckI0Stemg1TwuWw6hV76ht27I8i+Y
PiyBN4098awKm1jf6wzrRS9zwKPz5j0AK4D5x1C6/943dx9aUAALihRWSBUi1PZG
0k6U/Ek20GQUete0MbJIeqQu4RcOhwOFNoIL4D0WrXT2ktJzuuoE9N1oO5dbN6Mm
tf7STQf60xVif0LvV9v1/Y5qAX/7aEQ+m2Kety5PyKfNmAYYMBqlXTp+zOTkOCVj
IbpJc6++SxS4aNWlMSrbfAxfSnYEtPCDXFqVGuyR292geF+NQsbnX7894c6DuptZ
FYmrOYnFh9rRYaVZ7KpjqrZsPtTh0+XpZ7Vf+sdumeStmy3w3dhCSVtriA9jK1BY
v9Z8rI01M+Wl6isBimQsExxPYJFVVBp0tY6xCqav33lpNTLYW/qltXtL3xEeAnKQ
slHtGISJIhqcpLCqld8qR9GvfkenC7CVrLTc6+9Qj9pdFb7LztnfYI/FlgDsozrC
ZBDmMjz324AsQZsGJ166yR63EtvPLSO8tW1etRzaSWWeZ8FB0Of/w5cxXBBev1DT
XPq/5E10iugsBR71zgKtOAmQb3IPbIQze6whpGsLAQzC6uSr8PSdA2EQvrWdEjOA
5NbuWiXGDT3akVxRrfz7Jxh/4SpscqZzW+syFefIPvu2G5386+jF4EjLKOsCXLGT
av00iYZ8zVcjiC4X8M4w6CUW0yovBTTehpX85UR2Vf+BF+CXOxmIvih0JR23P63h
KqI4geYw0IzbTGIwzICFOPoK5gn2FEsIUGZuCCncueCuWQaezFqE1oGDoU7m4fUX
G7IxS3HQSPAtsdmHCirtAXLuXY6usnLbgXKGux+shDP2Y2df77CkJtXeInqdcJlG
bI+X0xGXlax43lPWWF8bHxn+n6Q1a7SJ3SYyEhlXLrG7WCqCWFrRiHGlOSJg66YB
0lgIALZENIBxjJdHcEfvOwdJO8yyG2zCma0z73heDB5w0Moub/WYxbsBl4BG6/Yw
adkwyR0gRWa8/a5dwsaglKy7XwDCn59v9oZSHHUcovU8we6LAk4rvQ5sTqGQhkWB
SPw5VQNujxOd+PjoPe3KskgbNG7eWU7tGpZ9To4CalNOBbiCuJ20i/H+0B0e8NYb
Tp3qmOztwJuB+0garSdV/A13BSCGafzmSfuQXY2itEgIjAncRdjzmnS0CrOjeM9p
iMFVPMn4qWoTRxJvryROtVVKtDdGk56hkFWJnTn/V6Q1MTrNJ9XmW6sXZug9KjvO
64VEp1qTAiMPyV07xEFSSRvltXOVlxsFQlKSsSLN91QlytQZgvbG//k+CdrqreoJ
X551gzDwqcWIa+HdeE8cPevbTEXQgV3+DZoBLZBUMXjejWeEnY+4wYMa8/e2Uqgq
cGxg3+bssP5UBVzgWbTzm0w2267yncTFprhxd3tqxYIV4YUOhY4o7rmKmMxrV5l0
jeWbrJ5pe5I75BspogZH5PAGcJHnTrk03AUA3sf0Ely1iq6vAZIMd4G52ASPnFbB
pqqO7B5BBQ5+zEWuSG6rPjbf+SSRFJ5tX1nVeTHT6suUfrV2vLSOx7YzKdd5/yT6
Z4gJDyb0tbIAD8SZRN/D/3u/UdJNRHX2nV+tjUgRU53u3GPL+s6vdFwspfquFxXU
cb4abgnAgzjgfD6SE3zCVmWCsRliBT0pRjj5SzAeVBYQfQwL1Y3EbAIuZfXN4E13
9oqls4cdq+U+loEyGvw6gAR3pZAPTDR/onE1ftilBhEUwSuBlEkuD9pn/hUgvAFd
tZe96wPs9jnton28AMCJIMbiWnn3pwCCxU5TptJQ2tRTM2gQ4gorRtGnf7zoIDkD
PqfNWDMAc2YzetwfrwwD1Zh0PKhmxIFZuKtWIEIVf1+G/ErDhc0/bUNg/9LTypYW
FYnnHAmaiMYw/Tnql+fCCI8h0LfyHQYpo9oGwVuFFOhOEDoAWTR8Z3QCH/06bvhZ
yv69Y1BDPy5F4sM2PQWgAmFRvgpjoSmD1s11WfQ0GXDHpJ3plrmMsJYxf8M5LMt1
8OPL+HZFY5/ZmZgPJMaNbCWfk1vRnATfvjHHR02gJDcj+ISWikxkrtFtaq+fJHcM
BXcIHwrS948XqM5IkT1iV4IrOzoLZv0o6sOxX8aSeZfTxVwpJnqOJwPZaM5Zi3v2
cvnpQlYbiPTCnQWJ+368zQqmnMpKSIoscioKxn8VhNAb7dEawomI2ARup0xxjEVZ
cymw3odeApA8M/Pvro9F7yBfT5dEYM/GRD57W4MU035ni9DP7TbU8g+oDXkCS34e
+2YFbkSjI/CHjmAWF+RGFllh5D8V3mcAyN1RNN93fNkILlvWG96xFP82TQa3AgKR
IluRK29m2t/kiIMVwqeNwvm91KZdE5vE/g+G1bvufOC8N+sX9kOjLIEFu6kQIvnO
9kJ1DvnDF9bGONGacAp7kdsRzDfXWEYKHWuocb05U378+eMvVbRk604FduC4OU8d
fco49YXsg6tl582jHyJrunP1t2Nf5Jv6Hh+RiWJryGvi+/Ye8NwaJgdOVHmefbP7
j1UkqlBmPlHzfvSEMjHHrTJztHrdSevuHqijYvJ+c5a7nUNtxxPisFXUBllPxsIr
RLlpsNqddiqfRGhszgki62xH2chv9Vediiun0dRZVuPKpmgY6EToMDL85UIWSAXo
Qqm3Zypd7FGPFFEYHxqARXeb4Ysa368O3VIY3fVUZlP50yqFBD2JsY5W0+0jW7Xs
nRAdpw4Ca/r15yQHn2tFsoXCdB6OOfOiuZkdk9ZtHrj1Cic16c7DTBA0nwyRX9fb
e4FuJbcF6sr/k5Lym13PGFF02k9J2m7mqJQdLc+nIx/OuoKMHgxyjZSQwKutwPp/
CLwvmwrXcP7t/0tIIxN2H/R7WlO2T0Qfwshyj8Ca4REKtMfi+aiskXwGsI09pI+G
KVuYE0P2TmsQNo4zVW2jBtzf7zzVuC3q2S5dZ0vF2juyBnMXGklIoCOwpcEB6TlP
L+IJI8eECdwAJx48YIxI0Z/RDHNO2drhjdGBMBqkfjBngDx0FWV6gfDZ2P3A/2sq
EaFTEyY1dOAj1Q25UR7QEjULpgHw47IP2KRwIM/IFDjTFaECsKAsYyDIi7lbxOgU
qBMY21uaSugGzUgnsMU4gcXhJmztdYI3RrjpSBD6f1Zvy2W6BTZqjftMO+3PeSog
ZQi7Sx3etKCggsvMP68WYl75xVXDBcmNF1G161aHR7B7JOzPXpuymVxFAwjSBFyx
nfvZUf8OrikPQYNVmfY/2bbiwQmogow88z80Si8y81o4VOVDOEm3tMIbVJE7QdBc
pYfWRMC/KDAlQiNdQZtXKkT0KN2nGLPpiGKP8iXSKucAuUl1UXq/T0Ihk+rZNEEA
GU3sj2XdSSLKUhlstf9NoKT8aL/eKM0rf2DiXyn+89mxc0YWRRS9Hy8f3Kmjzr0v
3jVt+7QZH0kt7L5hJyd/hBFt8kNLXLDk7r8Vv8AFRDGIrtOsjT7tlNTO6kp/Kafy
97GBVSwvPwuY3w02F2O99BStb3JGV7/6ZjZpbWvxP5DM74H32bjV4A124hj9D0Qt
Xnj0xqUW26SoLXhRmtrYpJrMUV1bJBJOj8LioOjo+zjWryjKKmSWhpfoLAWfO+pj
wkWuoKJavOBmjKs3G8IjNDHqupQVZbsptPSuKL6tscmztNaLx/nixsIyvz/MDH8X
+GZkSxUgVZofOQ6GNr+BIZ9qMBSXsvtoyLMn6/fknN7HIhVAp+DQlERMEIV8y5Xr
JiKAJwu9TRnY8IpYTrG7N3RJXbxDAIuY21L0TLe5mhOK6tBZVQdGG6P1H9A4zMoW
j4Zsjlu9PTK5ByGQCUlcKwJxiT9p7XavtXkw+AqBbyUAK691f0OMm8CyJxODaNCU
1yCupEiZFUgE+vb30F5X6iujQPkjX9P6s1Ra0NO7WUUAdWdUFcaYZR2+aUqDKjFm
rIs+kd4qvKfTgc39zLKJsZ7jhJc1PbRmeGaF01Hq2LHDMwTBuBa9xap8iub92EMV
Zu1UPPvPCkzy0yT94cl2/FpxmOEAiuZNDfJYmAI2z7pY7+Q8zJALIYzFAjDa7MWO
9Rqul7QSwVnAnrAWg14ywUnIYcT2/8hCYz6OQlllNjQl4NecV8gIadYsKuXSGh2r
Qx6HL645k4nv74mI/GVre6QqhVeAZVrOVhe2mz0810hjamV9rUaF8zN3VxKtvaPq
EBbiaBe8p3P0IVm9c9HLE9QnAAJop4h4GGJMMW5cDcL+BX6XTCT6Ja07bTPbcD1E
/ZHBvx1F6IAnohMhW7vB/aXiihArD51joz9kxxRQrAgrmtaLJii+LQ+Nih9y4sI5
RO79ZX6VUbVD8Np3OQ/AXnofPJAkfuu7B/mZ2RsG9p55qbbyAK7S3+vgs+xaC0B5
mAVwkKnUG9uZ0yY6mZGD5JDz3F+jwPAlHl8RIP78AUZ/pjfclTKK3tA7O8zffM/J
OisHsLgCczybkRtnvcMKSXOj2gjxAlGnouTvmxEI/9DmKjf2L52dcyiIo+EGLkGX
4h9MSOIZzV1OtbyKqbUunESbEBCa3ljTvDqKPkhAPXzpCLMrtQ99l42nORju84j3
BaqU+Rv0YuAHZ76dWjA+Wn9ah1XO2GNcmv5pg3uhe7CSReurHDuOeqcosQPG/c6+
OXHDGePyJDK0wSD4dbHdyHkoDQuoE1/+k86pHnMNv+9bCLF+51u3Qv4FIBPshXaS
bdQueIvV4So73P1U3okOEsP+y9fLEIjS35461iLz9gNahx0K6VGs3+gDO2MmoyI0
ZxPyeeCrrjUe8DC6RKWvONB+nxH8NBHi+e0WpgaRUWbLnSnKMmSNQQtJaWZ7TKNY
/hb5xDBZ5jo8Yo/KNcXovMfdn113RfrUfyS4M749jjhgSlN8bAEqY68ng1VdrzcY
tpW7hHn+16Bp7nFxlK54uB9hIb5cHvSfJCn6bnQX/OVn6zecy8EMy9cxKZJRcU8I
Rez5qntloia0gP1LerFouZRvzzlWCyPV9VGzqrPdBn/sm4yTJkVrYpPh8CgBeCPm
fO5dAZ6WvlWShrvOQMBQP+tEmrsBbjTZ1fcogOyCfFO5iauEMEEbe5BMu6fcB6b6
5E81+KTEzsDw3b3DlrgJxcvsQrgW0ir4HuE57VHUw6OURQjyJ61ulyIJfhPVdru5
cxcNDVLXoOuVBdVJg/5IQGRi3FxGoOna0GzOhquANYW5C0WPClHyL1vIUwT2zXXw
VzA85FHk9NzfZwljRMiM+DnLmiBhBxU5lT1T6w5g7AVyGcMziD1sqgmpaBuhJEsS
eOQ1qP2Y7PKhXgqTKmTC+PYy/9Wk0FHFFKE0sJHgkQrcHgDvDJkz+IhQmGKyWuCZ
fk7pSf7gbo1nl9qo28n5bAmnIJHV0lCHn0j6Tb0S2p5f2Vw8JgRz9928Ziga1bG7
Z/e//a1s/qLQwSsdEEoMohw/DSk1Fd4iAwg3Y7R8v68vwSIX6YWlhKTHn3x90PiD
K9RIew4l9UW9j+CiG31jjqd4Bam1ShvRqiAhRzYxX4Xsd5RrT5aQM/x1+3sNxHGT
VePjPAAQCiDRFEg2P0wbHFW9fRVIxfYwvimCR6u7X9eGIaYOThSVqqwNLZumQ381
51lKw+yBQfLl4XHATBbqxBX3uHBL02zaCeHaO7MxdpkQA8qtG3LlXmR11R8q1Emv
hzHOro7WZYKh+GMy0/dbtL8VBT7/5L84ieT4vkmvw2+BJSS1VSEl2Zb+HG5feDpl
h1gUUF+Wg6njAo815RptwAFr1qngobVzU32XceE1+JWp0Nif8d9JxbyFp0XBykaK
JmxVBhlf38QlijP9lr1v61tlODIySqFuHuQuCeZ+Neuk8oN/PhwEPHJrSiGvzzBC
VluwY7Ns7tENPu/EPoLlK0jId1vXJ5rW18qYmPOWAgfFu57yfMvcvkQJUiA6xcTQ
EodhWJne9lkJ1Im4qJU+G3nvKEm4owWr2QqlRCwnPboKoHLwGvaurAZ+fG490LsI
Odx7SZ/kzZNOypJksmiTnhBlKNwODoJfXgiJXq3D26f2aOFjT+risxm00GcKqDRb
93PyHq0RzQcioEAQ0KvFOG/bx4UrbkpBKy7S15WOFPTUP25ZjbBe6igSfPtsFiUW
+TZpNPNa01AiL9nZl819KdVMRy9p6wylWHbpjLz80gQ4qWxYh13tbbRHFu+wEOaN
EWKmNI+/+41fZsub8n8ehSWN4cSVjPceX3ERlvZ7voS1w1K44Wfb6w303Dkm9qgv
PI35h0xYItsbHudw5wUAu9mleMz7ssrEDmBW0R+WWheQXS4GBQEYNd9C9TLrXoju
AFX6Ba69xGtZfWloD3ijCQPLVZLmy6HCOHAPV22T7Um90dhJuFCwPtrtuSnPX5yI
ojEBzeMt0LOXOuCP3g3wv5fVd6Zr++pd4/hhTX58k4b4g3QSod/I0zA3uL4MLo+a
NZycE91qOdcqVqTSZqncF0c46iaUO66uJtFgfnQ377Xs/1+3ehnDEYkqLviQkJ/9
XV0wsMECqT+tErLea0fxQpaJRj1PpbSUxXrQyR+KQMCFn4O5za6P0TuJ5ozgmSdL
DZywUpy9bvUSK9BomSZYfcx7Y3A5/Y17rcU67rhlWolLL0UAaF3rKtAmXykNcibc
27smC5WpUVeTkaN2Fi75You2FETnxsUC5Kpo/xGZPhHgNJ1y8AnCiH5j9fQr5npQ
HUM/wP9fewuULO7oh7IVEdr172rdMgpoDVZdSomy5H/Lv3el0jwvw3Tzg0kjf88z
Og4zTBy/Qm5pkx9zwoQjnK5cvpJqgSnF763DBSyh3Cl3frXmN7SvcuURtktkcOLK
gP1rRbZJIpuRrm/QESJJmDAUvyvqbOTmAqAcobEHNn8CnY7smxnn/fHPrCFqGUR1
iNoAr7tfFS3BLfRWaAI1yyvUW9hc7s8DTZ9Z5ImUv9yPlWsN/Y6Yjx3PXj7OHx2D
9aewb78/IovLgCA0NqpTHVSkOyvtXIMAoUdWRTk7k/qiexq0aYNNcV/2+Pn9dIFt
ty+VuzT+sq+TF5FoC2ztyP/an2eNRkWdrw+qVOmBy4JVp9+NsrZoRbMSwdFxxL7i
ppEqE/YERdnlpwoP7gQARQNT96o8oQiCeig2efQ1RVCzkfhSBKRROmOPgWeseeJz
D95CTt9bLgb7RItDqwBy4ggicYenPNm872UHDzGxUFkb4IQUdtO4KMb7H2IfmpkP
nygJeAzJrBNzjagKNT5t9ZA5plwRRqC+LLirPDx2EMcHzqop1CDSNvu3OZ8RdTrP
NtKqeClqDxrg9cEX2nucR/Z7Ap5qTuquQ27b3Bqf2e+PjoUb4fnMey30T2ylantr
87w9Bm7/xmoiU1IwR3oXOjIW1chhaOi3zt8dVHNewqLCUyXP1UsJszQO89RP047P
cuxkEIFO0raB7VsmOqO7JEIxLfUzp03cXCo1fN9qorXXZDwho9EVOFYIxXjp0W0H
pJLVFng2J1EWJe9o4NeUlQ0gRH9EU6a8NuMDvA7EEnSDtgAMu19TL6VlBcfLbZu/
R9DgZe8OosopG6IQhZn5+tq+Z/dobf3vL4M1Bu78J1VZFhwulVSkoPRTnTJ3Bull
v4xSWQcIiUSoiNOZzRUZ6UIO+3JiXusVX0PICW1AukU0d2YDuU81D/GESDDPvSBe
jNQpzcp16S34GXblcDV/VarTkC8J3czPcwbxqPLdyRAKIGPXrHGzfZvQtIJBfb6W
xq+MUs4YL3iWUsikHZn8I+jzi+arHInUK3btLF0vanL0SJ+4taAxK/cxrmJGa36P
F/Y8VHps2uzl0L0d/QqL91ZbHDcpdUkAKm25DWkfrIGi4Bi/ioW7yCff2ZDg7W/R
VZQWxHrziIdf/AuSJGYznLWHwHPrq3tOXflMMKirXlKdzM6+lFyVcMk3vehCwao5
39NxTNkkPM6waMda7KIPATmaZb2MbUykn+dQ01mGG2Aw+xRfmSoXNM7LcYuUOWC4
we6N01OeLho7JnuZdtpLPzHTAIAArVuX9DfDADsa/Z3ktsxBqSV8Ji3rIZijguwt
QhTWvBkT0VEm+djNDwhr2iwCzRF+RAFawnU2HbOJX79E1KO9v5qrcjf4WATtYUWj
2wIVbXxm27Bnmf+h6WZFRYTMxUZib182S4LwoH1lMLpmNtbLUUoBzpzzIfqsKRWK
0AOUZhqdiGIzut3lHd9ktsYtjzwFOIc6GkDcWfmyJvXcVN0k9KZ+vDWyGRVYKVpf
Ypkm3OBRswWzht8K2fvyToz0Au7inaOhNHZkytG1Ea18hQAKphkawaXByEzNnp1T
Blrv9CO23AlKIMHJatpDrZXl5dzL4ZT0aQ126wk9MtRGCA5SNNtvmW/7LJ96sXHw
LkL1yaIeGtqltuOdrvLAsOX7y3yhNp3x30tziChLZ17FrkYtLaRjMFCRahg4Wdov
QfGiRdEOjt6V+BRgaF4WkDlZXE1q914fhYTv1HKx8fQOengEN5ciqzOStJv0t2j8
GiFFdz+AfDHbv0d+0sJJmanX2gWuGY8HGNnbAiSrJZ70Ab8bUwEHoNpBn3nk4YKy
39z386BIyqq0LefxB5s6W/ZShM0CiLJLdFetYttGPd4rrp1i/+KOXvHVcKInAICY
A3QN47YLY4TYAPxi7DLs/DUAhU9zBq5i0nb6Q0P6y1DKSAtAs82/UdPR8llYRR/U
LZOO45GBTNp+ymUgRBeF7L0tOoTgchBgk5be/n+gFNcim221oZkenfxnC7Po2ut+
gOe1atvQivoVw9s44+pzbWLrApHOYeeDcS++IkRp0hwVG5vnSvJ+H3r5I5LbmXMz
FedTh5v5mkxILfJS4usEuYtoUTAUGqHKTW2XnItpS7TJZarh5O34J8DvLfE6g/xf
lDmvFahWK3oBMFx5G/k90wKhP9bZ4ZjawMk5uAwshEemZSn79zFolF1swsMwVpdK
NNEYi/+aEaH7Cd3fuZ7xRpwLcrT0dpr+FSnNiAUL0EtvlitjT6dIKGH/vO8cjWCD
0lwkvoht43BvvS4cg5Arol8S2P/Kc04uZT3JxcmTQOwFLpy9OugbNaYi2w7NcGen
zPg3uCa9EStECFe9ODdNrDx9NXO4ANWOLXeCN80JmK1Vurp40G9Ypi/c0wTpO8bo
Fe0NvsSsmDnDtA2qVcCi5Iryg+jz16nhd+AuriTX3M3ZQRLTLGn35e7bgLwCRFlF
NKdlnKSRRGM6SQZJyqqrcvJ7DVMYNopONMDphY0HyOzMF90qSLuNy7rDXGjIAvN+
vX88LsS6aVlC2gxVWFeOGqs1rQd68oqWiJNrkCb/oKgWUfcuuRBzI7Dj0dLJr5xc
CyAIIHbDoIIPzVEvuTbukryah3suLINkrz+3rDFm4AAG/46Z/C3B9DKTv3/QO6xg
gz4CyB3k+IuLq8mY4+AX1nKSbdNrABzjk7G96/5h0DUeR3L0BndFJeZVNS7QXDOJ
oTL7QtNc1jgah09IMSVTJbfYhcGiOwA+scdPdWFjErCPqOygtgcJKWTYRivqx4nL
N51UDvT5JStA4aJ+dMTAD9+CvnMoUd7hPrYrn6521sy9Z1xqRajT6WKDFNgBPpD/
IH8wTOicyLvEeEzsilb4ZApF03QKb1bhI4tAqKEk47ss54Uy4YERfRAh4VVmktQJ
S3vHZ69ypOJ6fLpIQhKWZNBds1gKsPKkxA7z7hA2jX87MTd2bou5Ur2k/EA125AS
n/LHI+7CkVYQklwyklsSKJkg2TXZow9Cehs4rqgQpTz2Ps/+wsRmMcgnLbih/kDI
bble+BHNsbjjLx7cT+6fmdxEyAxYUxQ4usBVx8n965GIWXk4N8DA1G4HYCX0AOL/
dYhMbBYrXv1W5+PyVvjFP1C5URbk0Y/iBA/zHxfoT3XzDn8iO+CXxTHnle/HlYoA
Dg4W4Z4jZ9vm+LGtDn89hB45X8QjQTlN7uXXB6Q7K0nysbVOBPZeziToMAvyDtQV
md2GiQi4ZXQQaeQt2W7HOq8KTNM/Mzg3zGsdWlmLdQb2vTimB2LSvxKhO8zvnrYF
UIIkzud+lSrjLsFVlxf1zYN1PTeAfJUsvVbICoIIkInpJWiEDiJB6SfcxJC65P0/
jwf9M7s6cRlACbM1nAvPV372c+w4M2zQUlJJ1jWEqXYt+CZOdVKuHAOb3Rq6u+7y
ATcT1yXrzm/WUh1QV0zAPxxL1/wp3ZJYHMhjaMpU5CGXO+fx7mOL1XOsg2BLLHaN
IZYwv9PdwMEB505zdWJuSUYX11UECbnYBrSr/D2nzqvN/yPb/e2cN+9YG+XtNUj3
DeCWJb88s2IkZ5iP5QYx5YM4mq3qDr3QWzdl2uLnIZ4MCo8xyJjqdkJGQLsyhS+D
5WFE4HgeSJAC8mVqtSuXaJAyGWoUIwgmVvdYL370Q+v+lWqkx6DWr9i0hbIueqmW
qkB9/58XKSxD2tXOV0wQMBNCMBSU2QEb+g+7vuwi7XEkc1ZvtHy1i+Fe/X4XFKrm
LPkAiScpf1A1KncYM2W9wvNjT8AsMWvNfuSnAvbYFwS32uJJidYtUCLYoqMMleDU
tFK42uU418MOFpHGqTFXVx8AurZPIlV0NErnc5kNFPdpBlWQGxPRSHTEBYQs8NCz
5ICSLHf76KAHgaYh4h9/1tIpuaWe39O9sBn+HNen2qJBDsRFIJVN9I+vrP+0CWjK
g8BjeBmp2Ye+OQA7x0y8H5IJ2IWjqrgGu6IJexIlBlD6jgMAflxEcwN8ZyMEYsDQ
OVzTCTmS3YhjTtkZCjHxfB6HclxKt7HvTZBy6u/P5WUmtMCV+bRMUiTAh115Eopg
axhfeaxOgoz5esyvQV38lAulQcZAg2ljLkFvhiyJTcRSe3hXZ1ifTtRdi9p8fakV
XeVzet+JE7pHRBElwbeh1WNPLH6uJuLoAThA8XVXAAnaS2E9tj6rHedR3SDfrae+
upaEzfcEZtXiwJmee72swfCsuEH23mbqcuNpknLRdESqZPoscGMU1DVoDrNGGn3r
uxIrYZxnzecKLKL6CIoVhlQOeeUSwMnqNn6WMGB1MCFP0rMt9hkGHAypox3JJhsM
60CF878HXlJR+pfgKlAnzK5rXPo9Iu41cLzkKP07duE35AyhihTjenmRM0vhDOdC
0PsFLT0rSgyPizMJQtPtHzv1o2fshAquJxGzAgjaapLut7iMuCdP1PKFe0FlspRA
RJn4uODB9AdrQmD+2oLm4XTlXNtMppgo9fH4GqFO6f42dpXtGiuQZPliDg2sHOYP
m+oa8F0gxRHqZ2Jgebb3EBFN4xDRYSbWiqOSEbMsLsYHfiMRZJaA1D7d38z7YIgI
0K6MXi7MaMrE9fdPHjI1LBA3UnSmFTmVXdtqLq0w2knIF3kZAt+6KrKeUgzB81z2
VG2Kl1WleL/twvxP8zPyr3WdIin8o6AhhoeH8pLslECqcZ5ffY/aRODlACAwAKoe
6w6HnJ0oemCwn6fybc/WEUOt761yFKQbqzxJyDlGDvdewY0gF0PoqUw3W79boNQH
zTnwdwwVI3YfY4SZLe8PhZA2Zhd6XzeQCBRRbuWnrQ4g3otGEjoLGvfe9cfH5kwI
H95QnXtK54cWy3y7WYhBXBcMXjZfbz8uBAb5KCh0WOUplCCwJiup1JEgpoyMsLRv
mfKxPwOCxHi9uWJdEaUfb4A8oh65wmFLirL9lI5dqTbyn3dTDyN61TnCibNJE2VE
Yky4TUfvGL0QLEtFmDWu/+3qLwKljvhQCpbYEEFEiZVriV4hQJWcFc5HZnzsEgGw
azDb0g03jUqPBQO4LKpCAETo8sVD5pxXoAJMoKe8QEcxnXuTQY2wQyt7fQ5eFMg5
WF0VQ4l2JccRMhEE4oOSh8lbUWFGs8dNLX4+za8H7xKYjhRWNgnKAL0R5ncLMWks
cWQ+R3E+6IHt3PwrLtoMNJsRZLLwgdPD71wAR7MglVNQsBNDme3F2xIfGp4F64/e
PLwvcqiHWh9/EWLJrm6zWCxaMo2yGESqN4uKz6UAfgiktX/0Wb53bRLNqJFPWg0T
4+NuhtHLpq6WqPG6PfyD+USohYXngaaWTW4a0yCJZSleHZVV8MFXOlcer8jfcTJh
pbWUgiTPTJjuaUe1+HupBkoWrhb2xo5a6E2ErVA/VMRnNIgEeej4dlJ0ZM5s4C33
GkpolVI08ymL/qPVbmnBykj054FEp4uZNt2MwV241dqcuwvPqfWhGCBDkw9JuuWZ
bgHvg1n8QP9V0nwPZ1BPyhxsJfblxzLl2TgZkKXLAsQLdZTtOYBbewWyhrO4y1P8
pW4hXSEImULH8oaKAgCrf9dAK0U9RlUl4u7xW82uIOrmU83Q16e3ujRMtG7oJA7X
PwNZpCgGO0d1mPa3MQ3NvrC/tCn3EwqI41HTCrjd7AwNjxnWR402R3/76h6qTW4z
JUnNbGFc6Fopo8z6wjAUg5XAzeBimQO6Lll5AUZiP2X/zhANmc3Wmr1cVHp1TQa7
5o5Z6KRQIvI3UwAXqW+dWPsDcDGTYTbFiGc89ncoOOuAuamfCVBoIq/05vIXaWuL
2U98lxb8B+TIibCpoZimdx1ClGAfynbezfkdLbALL179/Vd6DiyqtABjWENK6+b2
8ihawDseqzNoNvdFNjOY5Lry1uxzVeG1Jks9wBvNkMFFtnky/F4WJR6sQw1joEFC
mcpb2WQFB6Ae4WogWvxwaQXw15DoMtDrqAIOlpWR6GwEmFq1IseXZTCxZjF2DQbN
eRgDleWLfn0mjMXVPUcamKEdG/ig1sF5QyEvy2LmDVSa8vWgbEYhBslemZjuvhvQ
xyZOw2jTiExTJUIlbibprTo9CgLU/9BUs97Zmr0yeI5dGPpMXnr5qUaCw1Vg/85X
dZgB/CD7Yj/W9L4I9NvKSvyek2w3fBUHIJeJkS8Mzux6eBwY9qBSCPyIiXBlqZp7
9URbiUBDZCbxmmYxzZjuMYGuiyvRWFxziQ6RN1WUPFrx+7hzmXwYh2tGTzmofIGc
k0mXQYjuh6zy19JsL3mP2QFNK2Q7A/6wfbqEb0HHSZRRYSIhHDBQypNpvYrX5Qb4
yzS1yKcqDyGDT6xyO/w0X7/jEpcqtVbZhLK8YP7rFUE+4wzOtIDZGNUlvHRxdFhQ
CjtdJjsV6GyQd5pVZG9Qfi9lCEKdpI+ca2dqtZV2Mm/pdz/nevEP89tA34M+ATvL
j2EYnYrobiWcJMYF0Wr6xXLqMpLl0VXcjefctUJsga4bnWM0ZBU83vL9pOjOOw0/
2IGn5uGO2sjFHiHIh3UCZXOpqudY9WT+iCvSy25W6O+qFMjTBtDxYgMr/RcYP1X9
V2FEy0VZOJRo/nyGNnQw+WYuDR39n824NwFFXqxucvM3Ol7GaFApL7wBO9+CSdNq
nc+/XvPmgQTo6Uj7JfUI9xC5BfLrvgQ4OwgBe8oEu0jpk04A6ksm5H6NXW7V+fvA
/Wlp/gNfwNzuQ63/YE0uG6ejiN8MtixaVmJjpi6bc3+6AzXhkYX+Z52W8ibdTbfI
cGDSivEK4p8/ZGguRzaN64UUQ10R4+FFHnwU3rKXBgrLwfl7x/IxCm1GDIRzpug0
6kQ3LNY9ifimDW82XtLAs8PIrJ4qz8IrRlihz+Set5zL4DdcFqQYzdyqk0c9EW0q
DvbhndXbDZz4/A/6bTWnwb4bLuYLjSrP56hVqkGg1y4msTqsSTxKGMURSa7U6TBo
x0dMw/BlpjqBBfYzLBoinYO2Z+7i8pVdJdpLbs129Krqpu7pnPspZAdcNtoPE3qZ
jGk1xlgKLkbkzbULpgazt4CZKvPLhQ6cTbzEAfZnONRk5tTfJMR9umKFFPlPQXdP
V5FMfT3CJR9NopU7nBEFYKrQmo8ErWepfXbJerizfDh2ULcJuwpi+ykKNgTb6Q3o
fiKBbL6h2cpqslNeNcw726GVsx8CVeN/mpHYsimnd9dTF9jJT9QiVxvC92QgU10n
wtdHGoAU3wOcI1jTJ8zS2dwtjOzzLK3U+zdHIeFidW0J/SULvvdloI2dqUm4uKnB
ih3/at0UkxuaUbuWltX/3RXXd1twvRMvsAXzmOnbtVyjiRpomfZsHufCs1aCc3PE
jmT/oxhnO6CPWFerC2s5ujrGKv++ZP4vP7CDk6S+corfPHCJ46YZLkfh30czYpyU
rgazt3gLDbNfV+9CYM7o5MUyilFF0cxbE5+1XFw396UHKo96NVsxE88IC5nSvo2q
wg0tPVZEzRA7skXmrh/VQZVfrcqrEERleAvAyNDhpK6fVjziCHTfph19e+8fEWnc
jZtBfjYjfvB3sWRmZ94uEU0J/ENPu5D6l4Z+ogMsQ4UJfHpLddypbokM02ZPvryS
9jNRpNvd3TanoR9bSLY77Mps0HQ6N8q7zt2RSot26ZnXMSC2IDGYnTRzrkT+z64y
9DD+/LIkSTtghSyVhLdkKgsp8aE/SnJ36/eSouEwVeSBC8eL0NQ03AU0fqbtfCJr
vh5HkwvLRhodfnNWV+nlzaVFa/GbxryUPBWTav7g/2BY0M2PUVJSjHhK/YWdcRSx
g6BaG6g0v/DfWV6vjbqZFgbWgH7fHyORdMX/j6ePVYryDnVpGAVJ72Tgj9ZKt+Hr
WTCDiKXOU7vTull/fsJjcC4lWkl3wtOGzUpIpHbWMhDJZgc3jggt7ZfoMvEMQK81
O79Vrn5WhAW90gqQyKNAwTLrAxWeerW9z2XnASs+cS1iwNJ/5j4D4hGTz4XRVLrZ
dXKFGL7wNCLFLKRYj/FFgDt4uU+2w78Dn/NFb2ksaaG0dSy89Oghdd4KBNyeY50Q
djeMwCBvgDJBjEXMld74PC61qj8xkXPkc7HhgpqcibGj3rkkFWi8iuSkdyHAO5bz
xfFHsq0BKxrf8KatonpEFdH4PLt1SatTorPUcNT1S7gOpBdFj7UTUih0zJT7LWcY
lVUnkIBaS9vmJL7lrLdBAEmSBdwdx4U3xjCWtucRJP4dTeCsDRwkzI7Mp+fIdm9y
f2XKsV/oejO9bY2KLQkfda+59Aga90YmbzMhcMpG8/O8YkXCZumVnDvxZBOBhG31
SsFieqNLpQvpFLUCxaYJdcGCoy+htHTF65t/NS2hFVDG/m8UrDvTv44spA8Q1+BB
q6sew/ZVlnfGB2roLmXMdW93EmsGLJyeAXYYAfVGeWAHYmCRtKICVWJdIngbYAYI
EpP7i8khgTB+EAkTgCbEaQ+y+OAOsN2oADN+kuFBy/5o4wUYs2dLnWg4NPG9BS0D
G+ahqSKsVlJVkX1yWlAc69WJxJC8OTgVpsWPBHWyIWz9SWrIPT9EjZFEJbOtpl1W
CMFCki0O2ywVLWswV5yS7fZGpT4OSPPfCq35esgiainIyHZFnjpQAdQX+rO7dVV7
8rFKCF+X/UMuA8R6NR47KokQWEkl5As8hNK/E+fM5bFstsHA6kE9M/s7lmh22kUe
G+tzyQMjh/fM+WPDYf6twTzqCFEzzhmqiG4cgomq/2ERKNWnlFnPSqLo6ukltFv6
GAuZt0kAX5aKbz9zfW2YooExUyoX4qlXwXehBR5ZBDaNJhgvOhQfSrSjzG3zDARQ
yT6MWjrA1lPcSa/Or52VATsp8W4/4BBL/wSQzHKjhnsVVKUK4FRFaWKbZ8SyO0dG
UEBvZkyD0ZftAcOg5V0oU+fW0kI7fpnaCewQVg+pHhD4GPSiDXUbGitKJENJRRMA
eZ76nqN4Y6GZX3FzjYPwyQPpncziZv61FJdrwJWwSc25xqaGVvo1QncPwZWfggd5
CHC8uhdaqfnTt5U4YKRKwiiExr9EbaKjuy+kvOJ8aHeWaaE9CsmEupu/ufhJ/p8D
Sv9gligr8kzNLRTm1KK40cUoCxouk+qw8asg/eDvq4Vrx1tUS5jLusLlud/uixve
FApDlmRUKH9xTe8L46MRWutpG3jHqwOx9DPBoCIrtWpMIXmtzUNSWCPDCyA2Jimj
MnWahnXJNAP9SozFlVszPrPd8pXJxCmqkJgLEf88ZTSDIMM5a6EEAUVrSB+MND/Z
VGEZA5FGWNS4jGDaiBVt71qFKvp42hzwtQRvPAmNN2q+sSVCthtiajRr5m96UkK2
k20JCkJmmFzb9bCBxkPgjgDzqOM0ryl3Wfj4UNH4g1o927BuYAq0QmnwsskK9gc6
He3IEQF8JgvWjCdkeV6Uycclhx/twzsWnsf2krqwbJwi/7miFGccSV+kZQ4lRpyH
rS1SST910QHDKnB0f7dsINMMhB2vLC2zfxCcJLj0/uatvOaNBLTKSxaMhQh5MOqd
+na7dVEokZg1LIRoYrzcfQpnelFiLRUPPogD92sIdqb63JK5Bkv+GCVWWZMMeXEy
ab2HBeX26ES21BpomuKi2VVg1GzxELu+pSZjcpFqwlm2HUgQKXg3gBQNnNwupD8M
I2FW4aJZQsigMWGDB0UdiHJZrKoyVAbWepesQBEPUJ/DLmVZZoVf70Z88WAryqtq
9scfnooxZL5WeLRZBm8/FxFhfXm9Kd46b7nnM1g1XsGsrq4DzfUhv4IypTKfX8C/
Hp4SLEJao5oKVlpIQkIWdObNWgh5cXAgChbnpnmzbe5+rJ2yenqOtSc4OhK2pkTK
oLeiaZIKmd0UFwjZjkRELLRHaU7m1AOEHcF+2tS+jCpugmVyqrLyh7xQG34hRZRD
DzoQgOj0Hz0O7Ud7ezeOEgzlNRhHcSvMkA4SzQa/sClpWOarwGBlz+L3QFUBBUUX
kY7SKsozYRqDqJ+vW73oY5KtSmNwV0VPdORkDEs6zvQPLjn12KRUfBfGXP1vc2Gi
/IoE7yc+zknjcDA6JaibGuSANR4HkgliP4K6ZLcGQ8vx74IcwkEu87NoU6hAZQJK
/Kenx3IQkZrwt8RVZCYDXA3qRKG+JrjQqmP1xAx6tevvHgctqksSPureUBMxTlmu
HoONbcxE5ywNe0IMi0Za0+MNJoXhnFTycqhlve9NGLAbcjs34Oz5p3i8wTXQIWfp
z7nyaeEJKgayPXIFNubo+8dbD6Pdl8L7Hqm2UJAv+cpVCweby34T6DXAulEir/+S
E6l7KMjVRWYuDizdaOwyYCJiOMOzm8+IGAlNixpZkr+ddSUXdjbMuyC02nqcRDa5
EtGRwq+LiwKLbJD2qlpDXc/ur3UztMTr/OLCLZCPvUafb4Di7e2XgUQnM/XuPGIF
TzY6uM55kvUHOGGUplDnVeSNyWlFwR3sokfaTt39Nh+l8q4VAzxxyawfdIQiV0QO
2bh3cHn5d/qKfJUECwWgMgXJCjbPJD9MapOU/a92okbEBl/AilLgGYVlaaxVNaQI
PFu66O5BwpTA8Z1quh/l01490oR+urQcdXz2VX9mVRj5SilpeXuNz3JJ8/NruToe
+zXO/SDotKK6LTmpVFs0su7satv2RM0YV8gfMJKeI5dUKS2mOedbe6V1fNdMRETp
yPqRpFueznEzXuCj6JiX7WLmNRKxCH83z7yL22PVYAbGOynEmP8T+oPNhrA9QaSl
EcGh4g0oHNYZH1hOaG+gzV7UfmtrZzRW4QCqfaSjMMeuOcE1w6GCAWrV2t/U84pZ
jGSEXjcRtv+eUrR7jYX5NnYkcWihyWPl6edG/ul9+PHMdiit52XsO1Q3KiKuEHXX
ebB8RnS9vWIMGY6Q5m2xPL6f8lfG6bBJcZ1WP+PpUyVA2t18aNfk/UQ9eUn8ISLo
Q9OOrsBENvKt3SVpzMqBzE0gA6wo9+a9n43n860ln7AISTa/uyeigkpLv+qXh0ny
CiIWnds4ce23TWWwwwTKt9QckO8NptIPya+XJJPAac0WorhHA/fwJtfCgGe0F+xH
dQF3IenfHtaxeWmZm7kX+uHlEHV7tdcjoPF5zieKjIGsleoAl2NrsO1LIH3RGNJj
GpZ49VmZ/5VdTFyjCQ8UI5x6BQJwCgmR6w6o6uyjjqG/3rePQr9GrtwuivkGldCv
cwHldNNTfYiXRNi3pbQWFQOmeWyRm9FXO5e0R4kV0x+a/ENwTGutD72AmAD8bwHV
UffPkvvff4AYjJLcc9HZAUreUwAvovoVeqyL+yetc8J4IvdL81+FWalcuHiZoDvd
MMKbJYNjrgtd9zpI9DwMQDWYb/n7EXXR04qfucaP9GQ/NU7Vf7Mkfaua22G5iD29
Z/bqn1CoW7RjsFI/5LskDYr/3lgXlHknXyjo2QwrPCitd5RZy3sVxRjcoj+enxiV
iaxYUBPG17d8p8//gJNnlSE4NiMW385CWaV18fLy8nIVcY1h3kzrcC0Cw7N66qci
fnxrJvHyV4Z/IOB9CZUTVoxHy75FLDCKuz8FwTSB2d0ns3T9/YedAGDa9u2avpOc
jflVVTG9BczTpT/nURRpEVvru+YotwFZvddnln7ZVhNu/tZ0tBHh5e7fCNED1pQl
BWj71OiE8V5Y8bVtfLQxde+3Avykv2VOvOyf0pVgi9EQPWoqk0uP4Cr+yyEZTOEK
lymGe1vG4XCwMwyzJnKQZo4NyLVJAQhLHyQD3Daq1fYcDmT3KXhR/CwZBj9YzePx
EREuSlDnEjMr7K5jP0yywgCjx6B0S30sn6tX0wAKTjxuMz9pxVrCnEv0Q/hDYgEL
e/XpRxQ+AEs7nXMLLI3GO+aatv1Y1nB/wdcIgX0sDUy4DfgT/33rzrZaP3lvYc6C
V6vc1bBTUtq+9NwlAuv3lgMwGpSI5iewhL7tfcQz2pkmtKXJqMuFaNjtKoh0X7Vt
NW7MukYUHaqkAJeZZ+czSOMTp0GaVU+XjKzphedfr0+D5lg1xPWEgHSHNP+DdpEc
3OcUF3ChW0560UcQkSuT1MDw0AfwI+JWx6A0yJjXPs94Px55NmmN3toApd8ztDan
2EXmJdUilLMBBzWfItZZGzOVPd70zudC2pS0QC5EegkMk7U6NFJue/SI466KH1yg
x5yn2diQPBT/vfXibcxxZmbUDiiTwOyqFwv6N9L2MM81ZgnxKYw3b05Dhj4FQCe4
ZSNrBE+WR1nj7Dyk3lTry13p+En7rxwcpVBBftg2gMh3jptGShOInUQHVtIFjPEX
/R7GwGCXaSUshe7bEz/AsmmHGVIoV4tg9yOTNIDTxpPg7B0o1ttarh/G2wibTwz+
WeofQ6UuAhC2/mpf0j4A3L11ITFpmi7kce8NmNW7LZAEArq/JiLUGrSoR0nypbnK
s4DnMUBYLu7LSbqKbQovroh64kOfWqxCMmNOQIFjhsDvoBHNLr78nNsWoVKGf+4S
ysYsF5cfnS0G9MXkC0dYFmVoUHfAlLj4kGAHxolDEDpKvKt0tPwkvzb3JXcmvsx1
JSc3r6OyVgSFOuDKTIShMF/KTe70ULlxt4aciIMOuIH3Y8K6nsvNakFLVD+eKs+Z
IV1A2ojCKVLVTZ9xbrNXMH9MAylIleRWrf5t3fn0HkC5sVMSecIU9OvhgGtZ9WJ8
TIkHZBpqPu5MuoL/PJzX4ffy8AnK3dcNI7jORwE859uwSjQP4NyW7sApYSLXb4iX
Va3j0lCUALyvljafE3IL1fDsj/bH6qhg71vXd8rY/FivwvxveMf/kew2TyfwBxtu
Sv3+B3oYXgCw0pv6wVoi7/okXDLnx2Ps/FO8vehD2ePu1NC7wih7EobHqrtxVLLF
N+9FDQAix9cBTaQE2kHvNzOf6opHevs9yBi6lC5RvjnUkqjcsEJRgCkovOmN3qI5
jnPcKgDIabTQvJaqolkbuEurZa3dldBRDdkrkb8K1ZsrRvuTyOJYk5586fYF30cg
9F4TS1Rw3gQZh/9WNyOU5NjIl+faU0rZNduOZciVJG7xdwMvrUURdEGWWqRZFA6T
syQubc0bIYeD3++vqpteivJxqDi7ISusvsUAPQ68OHya0Fx1BeANwCzh5M5AXPEJ
Rb50E2n+aL7gsB+KB5W0hoWU3uHh4pCYZR7ZS+qKRwTaSBhW/dSQRdord4diJmXc
RVgI3WDdNjfJbHiyMoeifQeYkG+/11a7kOxtszi2LrJLsza0xYPFMcYAf/XSNtBK
b5pV0EGoKtNOYYOnV8wxBu0a2xCjiPEedglgNLiQ06YefYqi5ozpaaXTbPHhMEMR
8mhP2Wqda5UV805/8wGOVXbwd94hcv3wIbznE9SqjlmaGDBWI1N+jaz52HFpsxEb
iGkW6LO8uY0WgeUMd4DMfv1ZmJJYcy9n5IeWmj+6uaL9CqaXCpinBV5mNt30fJXL
SpNCP+wkufS83eeRv2oi3wNSg8cnSncISTSdjBXD6rN1zNBsCjotAZYIcDJBnncL
rW/qwbuKsUW2lDN1MpYR/9tvJZXNf2YokeHAckYvBX6AV9bDsN+7G9qnez4CFMid
O2+TX9jEQqQjvxp7AYhGTfeDCZudoPVKET3BkboKjV4wlJqhnTClJ804RBth5OmW
JxBfIUctL8PqeAZg8TikBauqKMZCrOqds3DJmSEDGPtwfw3EhCEo7dzDbcCptnlh
KOx9NKESPOK/Y5wt+58Sz6+PhH02cOYhtfrbFs5z1iezVnwOKnRfYYSHNwcLgQkz
/AlwgzCJYTxKu/6ehumPSfFCSLXqyzwkI4Aqsa4temgA+oIO/Uz8xdlAzTlRk0m3
8a3P4D3bFhZy/7xDXe7qkuOY9zd8sBsxF2WOBWjdOwOhVfiiS73SASXSPoi8jKqG
aV6SZrT2yGQSZqhDXirdhxCS/feD1eQpBZ5wuKX8q/fbTy/S2MxHg7/7CJBQXdAV
cnNka4fCh1Zz1q64dkClzP0v3aOmL65Lb/p6UgNI5wYRWSZCTEvAZ7X/wiB7D6vT
jHqkfqwL/T724uDucVT8DQBznwzuu5O6Pg1sKG7IlvJY1mf7YLEGU6FFZW/XXyI6
i9OAOBPJF7paPxruMoQeUv3IDMxoc59/JsROUuOJroFh6BV2gJrfqS0QKuP/jsTd
QkJzvvn4gVSCJIBXzuYYpVd1Zo6JD05LtiiKOdO5/whCcwdxVyaOb15A8QyL+6k6
OhLE2N+Inuyx3HCI6TbNqWePNCBnIxR6f/JluoKoPFkVAEjDWPCde//UoPRzbWSp
RGngW9yTgrM0sGFb4SmzuyWqReE90fG955AXe+E0LlPrHwPtmvCrswvt+8OGU6mN
5sNwEA9h2volVQTRkuWcCJ/M4RG9C9d/c7QrZ4XLNVf6o9YF6ph0ckifSUAAl2Pm
YypARsk2PH+gibB3OSnH3EG32BR8tN5cU/DoKDbsby2fY14RagSa0EFfVQAXguVp
XZ3Vle1jQxWcuy5OEhRkzv8y3l1PcWfmBs917CVlfSK25TAOX9UgOotcccdpgjF6
1gEltbBl6SJN9lj6p6T/Z/CXJfYN6SWRtpGBSOJBwrZVoujRpo2By9Y6TIoN8o2U
YnXwPFYiG2D4rAUAI6ypt9P3Zi9O+GUAwTw1GC2hvGa5PnQTuWvT0mwpTYFaokTM
J3LXfj86Y5eRk6hYcKsJGa4BNjhA+0UO5le+47QyKJKqrSNx1mJb6CxjTJJEYdGv
ZHRyyHNntlwlLqnnSI9XTh9WVxR0gVeP8CVcQPfH2BzXsx07PkIHurQ3xdRIBA2R
mwPxPitvq81rbBVVwAP0GFWbrAtOgFqVcAMiUw8PToTJaZklLhCcfLoYCH97O3gu
NEkXlO9hNKHn/lgfOPIKHU+Wa/WZTqcgSucCX6Lar+WKdNr55ZkR0iA9mDh0NlBi
mRBaPtWvkEHz34NscEwg2SxzvCXv0lZLKE+pAV/0Sim/XDMuPEll8YmgvUwjIPbF
pn/1EZGDygXDAmr/vTLAr1DDSkzCzJwaxYQSmnn0XMrUjdQtoN9HasWmufWzcEby
1oaqQp4lsb9nLHTqrd+KrRnoEWElLeuf+llJk+Dr8xva5CBuABGTXfDurA3q4GHs
oSIr7w3Yvaec684RdgW4E29TjXIdFgo3+i7TebqYhauW2rc9KloZFMZymjK+PTAm
Ni/mkL1jDAUN8NaRc/pMASrojlQHNaPqur/KZ+C8qntdcbRLtqA3aYangMYB1YGO
Uv5IzK5hiy+9pJ1RuWTyJ6ARjWq4EBa1URupe024BidUzZJERVrZ1vjPTVopEGCj
FYzfibNpatihQ6yPNWEDEQDJ7Di7ZLBzENLbSTpUBcrOoYwFfGvKkTkqnSBc/v7O
GHlFL1AO/F0o9o2i7/jFTJROaxGG1ae4+4OpEcWm+0VhLJ28S58RpZWjhYkgWnMO
ZjE0zkedwRpHkfMHoKsmUG8JAP4uoVaWXsGEnxipYWD9gVRlRkKGVpqUR/zFtGte
ASedI8l68sNKUWAI1LR/AOdnyPRIFHtl4fgzSHUltWqrwvDDVp/9K+jvDG4WcJmS
mr+PKFdStmlJiKLTwSLCkRl3hLpNeyInmzHkhjMkE9G/0l3o7J3pnpr7mXmrZ5gB
0gpZHx36SedUtlzuGzMCLdP5s35c7QCbSF9pCLQ6SVmqDct7gR9SsDH6aiA/sH5O
5I/9Jwx/G8DrijpLtLiZ4u7e7R8U2a9W1xyVQqAlaXjPaCn0cfWjNwHRdZgEUCqV
FMN+25WPbZR1OUELCkn6I1C6fEbQH8spBdXhS1FsUMhv0KZS3+PLPTazFfRfSd+j
rjDw8pcxOtzQJH123K7OqpO4aPj97Mr2Y9x/8fihOSYubQtT5wNIgdfrE4D0ET8L
SsunRPAnWdjOxFIa5ppPj6wZyJoyf63GtaKK9LDJ0SaoHDUKPBeDkCY9/NNlHizt
mO93nyBcqBw/S1gd1tNp2S9maKzUie42P4+eXO8sRRu2hr0BxRhdQkTswZnha2qn
rozjRlWQYvSh8FAgO0xOHnRUjj4CvbLUTMfMB/xhDewzkpzd1KSr6SW+dlz9smKN
CBRZXidm+FnnfaLziV7kD1HHIF/unPTmNFtJw7+1I1GIW5t9DmFsyiQ7eN8zJr28
CoALpLhQBQ4b/MEqiBKV2Sjk096Bz8H2MrmVIQjtHr7MClVRumlLW8KmvHw7gjnK
ZVp446XOSqNlXgFyP7pgEkYb6ecLyWLP6/PVgYYrLJC8y3p4Lsy1ymkzaMs3F0Jm
mPp0+KaNI7JEGMknh7CAdC651tz+OFyrAXplGKtnyoaoGf7xZudHKGZ2V0sLvPpn
Wr3ygXS/puJ1VDi9iwl7OfiRxMDBdLevBbQgKUp4w64A9nzUOB0GvJ0Teah1EhDb
sjzP3kP3a87uQaTRnsPM7RF/IkqmBVZoCLV67ktBqvI4QpQ0Fpe9aD+qrb5YdylX
4FbjylBOQ1cDQuRcgfkUNjHfgxdBDtFgyz2E+NUWQ4UjP4qRjW6aym1JsxD+IHt6
FkkYHKElgH9j20m37zHJ94f/rqCaQy+qLeqGHUae2MmAbkSpFfge8fufXZW28Dl2
MvP25AW2neCQJQB5uea+0OQkYr3qEIoik8/LNmBjt5VGj4YyeLzUnG+awDTt8ohk
PR6eoJDtlDZ84nEWe0fT57HM9jX285U+LL/WphHNW+qKzYAzUp8+wV7C//+EM56+
ILfLWxRuOn/nwV/KtmZ26agR5gselw2yUq0GH9mJj+3JqSLkHSIAAw7qRHwKfAHG
3MD9aDscZhq6d1XpVCsN6H7eoLbWzmPhBsQQcBkaXcFJgBacIxLHNuu3nhecvYcB
vBP0yqZ28sFjX+aHgIw66CjFzwhNwaT6ARNMQ2fwCfrN+XbfJu7ys8Qp+Gz4ISKG
FykPSrjoQvSn3e3f2Z6VLxxJGyXn6BSUyPpg/w+HPo/tqwfk8MDJ5GaJvVeZK8e8
jh5WQmcGX0NYaE/HayvWvCwwvJdMC+vN+bfSinW47yWznAy4kTVF+hfHD84NkyZT
HeinGmTu8wLXhlpJBRexzNjZFELVe/wmfHByJHOxZTq62YDUJA6I454qVxAH8aux
xB7sOwhb0rBgjW6itSmKsONBTDdsamYwDak9oEk6SAD74fEeC9DIAxOUxhIzBoeI
CD8onb3F8SdvG2QxJ6bw9qX9btfYK7ZnjwrYZRrPNG3LRmyYRFBUPkJuM+ElRPxW
yfxHPpa5RY5wcc5R+mxjHt06qz8oUmpWSjSCC3vu/29gtC61fdu9gRq1WEpaPCkX
QK43oSQhWO/4dZMBtJzUhx7Osmbb5ADNS1/e56BhyFoBkB/j6e1zhMTlIfmyaOm9
KFNPCSGtkLjJdCk1oiuuZMUNVrKP+wM0LhlfIeU0FtNJuajqcMPEn4H8pgz10SdH
+V1GuhuTyDTg71iETlh2UGLXCMuuaQaj/1LowPOZ2+U+EsrqZILCTy4PhYx9nF8R
Mbptwne9LmQDXJRS0lY9DT01Hnh6pACAHQkEpXlOKym3x6YYWVFDRr5C8d54Kvyv
sgX8gX4RThLwrV6h2LsuG0nTqXPTRYY8B+dfnIKNIjsVnPbtoFKG26Zc37x1e47G
LIeNj+nKQX+aFKABDDEdP36jXMnBEnd8tVOREulmu8ZXQ/V4fmKwv+p0Xjz7E+T0
778fN050EeZIQyKHcfebi8CpmfruwVmjAIYCzexvpmNZ6U2wKkK5YBsdux1zDx2c
sn0fZUcSaS35cYXipklgN5AxzTmSP44//MEWFVDbOLCAUPuS3QzHx08v088UEkGW
WLYcfQXYkYrehpfrSB1s52siA87+roiJkjq6zrdm5JR94vgl0IT+14zfFVmfeqqM
oqRBNipgg2RwrO/SrKLf9E5yjBn1OvupYSNaLBNkVNNeDiWj0vPqvE+rm37U6LeU
TO8yoR44wFbzPbbp1QV5KMU6bAZq3iK7oeXbBbboAMqWx/ZvGk+62cY/JrwPHw/S
y3pp8AQi7/s9F6auNHYMZzgsNZixoH7GqWCNF0S5sHYmnskICTxW3N2vxUV90+ob
p47f2TyIFzFYiLd4OphAAdpZ1kUA4zIZG1N8IbqPm2Xm0o86Yxwj8QDEP5gMOVgA
mV0e6bPTQ8sDZZt3dE1s3muIrupLUNGBz6PKSVGjrdAvJ1t8Z0TH1tgoic03G5HF
d2uLGeLX64H8h++0HlC7nQPuiql/kYbSWgenGjGgg+qqZuXSiOmpdkwr7AwrPQ7t
aRXIrCPaTOq+rHLiN73rKWKhmJKJFUlx31DUbW3ZexL4TciCPG3RGjmPjfjiqaEj
w1kNa7CFX/39XX3NIGsoANDVE8Tpe9VdND8JRArYwXkDX91Ku0VawTeSk6NG3Gai
AE+eKC20eTJ6Oc1+QGtsD95WikVoMG8HSqYwNrPO6o6phrfuX0LRIVq5TuWdI8Jv
hPcuF15h6vZBhhr3cqy7VWa+voGR2sGmqLYDpipdPFIW/oTDxEyvt/MdDCRQDoBh
Za5uw9KXfmUkgBXzBdYAtxzFQhEtxH39x6sfYSKkLLMj+mWRdJRwwdW2L/3PMHlZ
o7WHsXhT8mRH24kHRXJbRGeEoTd6xg918Z23qWin04NseRG8dOva1zKKsAFzbhQX
FIKCTxiHMRLhvSelJvvbFDjNksHR9uofAdv4arF0ZVFbghT4y8SxjqyrCRu8dKvO
LRT55PcILYxJYWokSaWSGlJYCfLCwLjEoNLKeK47h0M0ToaztFa8G8IjlU+g7KXu
icO5O8YqnLoFHF4KKrEjZKXMe5obHIPs+IBIu4oQ/cn+KE5aAVEPUhognF6WsAq6
bVDuM/1gJW39lRQdXTPq+E9xVjPBYuPDjprtboPia7wFeH+AWXbAdEuk2XBUiWY5
Bm3XZJMVdsUVEAl1ORIwH8hCzZNA7IGLHpGLrv4vVUthRTG5mHCB/c5riawOTWt1
d65FhUBj4uk60xJt26Z0YNYxo6OuQbYfrj+DaWC7uxRjON2OlpFm7Wxw2nzbM027
ZlwJOvcL/eO1qt9uHr49Ap7uytFmtjQ/ou5KQDuoRJ8hP0FwqwQPGtXmFK+wtzNU
hvzAnFXeavw5AH9z0U5QL2o4E5pCwMHj7bbFF1kr+v8Y1gS2YNDgFy6IZhRRdByz
fYcI4lQfBJLKRytuOZJBJDgJQyiMncY8utmRvYqHNrdBlO4pw+yC1H379Z2vp8Nc
VsUouX7MSn8ZVsY5SU6pJGjXhin39XO+pZ1WWnvAjrDrLqVwODN0y08MIHQJvZZy
4V491fsor8I453v7GV0fXNgvt9fAnfeuAo6PKy44jWlU1gg4b4uFvFY7Vy+z6gDm
3BBXjOi0MOF02HvQjEabpTPNl03ugiPoqE5D3k8yNky8fpRAGXcCKN0YMfA4xCLM
v4z9GJRG2es9ZBdtOs35E/4SdZ+RHn3AkzQ2L77RUjtO9FbPMswPULajtQDGzR1O
iJRZYGYKPfEmV0RdXpaTk2F0AJNJ1y4xHblYE7wI/dRXOYU37NPSjMNHP/PP6ct0
bmAAY31mSzejAmyE6Qk/58WON8877YPdV6CkRdIt3SpexE9Fja7R+sxHEzGkAXC6
f+hcp3+MGkcD8g+nJpkIVgDq2vxDBVFqqN2+5y5DgIpgsMyceOZ9dwm5wEexM+a8
AY8nyqj51l04yi1pjwsAEbkmt+6iN1nN3Tnutt0X45wKNRMFKfW48p0lhMXL5oZ0
k0NP0hpQ6S4f+YrBoCwPrueKY3RPDwNatRwWW/AmpzX5h92UEZZk7Zx0BG4Q2bce
WFxs6kneyxgJNmxU0UH7U7Y7e9cqb5aDt6Ya4OTjP+NAhXdjqfFUGcu3HIHix+Yg
bQIyKJYbWL6e1qHAOUCF4IWvNFkE0PmRiObqpzAMQXLebB5HKYLMrDaam/bWgQME
0rncKd+50hDP82cqpDEqqR1WtITgcH1oY11If2UQaJEEkVMgj1AmZ5+c13DiUODS
vxVdX+uKp0BZBNeZExx9wV7I0qumE8mRkLeYEjfLeWayQC5Q2ezgd1+iJEC/ENuM
vCUrecryMD/vgGIWi4AuywUXnXWgMksPqkDt2XTZM4hsenqN4PB7kg0EHWtIdq5L
ivrWSTF/raX83HfHZP2bzkLurbFFxLyGYBK/wWeU3i1WWrb32mOh1vETPHbp8RZv
BKr2j6A5sLFjHGnor8srk4FdEHS2qRV4AqI0GMGLEU02XZLZy64u5p+DFqW1DqLd
g15blPZl05gITl/xQSKL71HU9ZgctXuYVRrBa8ihU31yMGqQhwQiXqaCY5HjcaDA
YezdAn0ivUYObAxESXnyGHePUl/0RuoJp3GnaJVbsU+U8DRqGg6Ug0wQ0RnzcmbP
tTgTD+5eqsD4IpvaFkMIZ1CcuPAXw4F048/6YAtPqtioHtIzGajqQkRlCh5Gd3lb
ytdh7c9QfC4a9UHipOInaZ5v44izf17SiWHu+sBWKqye6NItiSCrgDoUEKDeUTR/
8v7XRgpA0mBvRbvGyPiGfC1/PhYj6zmxTpRbh5Vxt0IxlzvexwAIpjyycS7mxl47
qJHatBuojPZJMqnTL28q+sW0ntK/dWLOM7dGLfDw8tifwMPax7jhccxQTG+Ke97F
WOMLgnHlUdSgcZ5x2jY9rpWmDB1nZh6/PwE+MPBNi+G6kHVWB2QyimahRhGXuaTK
71BN7IewYHhxsDxbeP0Y61F/OfWE2O3asqxsjOnd5dMfnCZ1OBWrK/g0U8iuDCtX
Sqi9IqcA2S19r/T42lSErBPTd7nlLjJjV8lTzrARBLLnq+BQVhm8fg3RfklTfyj2
tK/nLUFCPhWKtQrFUOomb60Tn2DYlIO3RT4ugcJjUW0Mav++KPj/weucealFy8Jw
y9LTl0sTIIp8VxJFxOcjxOj5GkRvy5wL44NufDZfcHBwCRs3aCUQ06bIxXIsjTkI
AlSnDeFirKwKoS86TDPaFqAGe0kHPcgrzXjx57w2Xy6gLH2h3RWYHP4szGYxmVxU
+SdIuzcjKd+fNjVmU7aqpmMFWQAPpuoaf4j94sVHgOFGjDa0aJ/a/++LzpXOWDid
G2myGX46xhy9gjmKqbsJN0xAx1yNfe6C9qvyF+K08SeKgF752KP+AscmJUJvRQFB
bs2oedpfATmQr8TRKddwENsxMzLV63oxXgH1RQPVN/7S8yOEEQzXT+MJ3bngPhv6
a1LRgBUzBcDbNDU9dgPl9ZImlob/vdhYETxCIOe4M9G+vM5U722EuvFxA+vI6R/v
+0Ffu6slfL6E5MM2P8SVyOsPBboO73BIrD35FiKKqDuYoR5SanX5sRGAifZsucBU
YSwUweW3WIKinAR8DIXLLfcZXqaXs0yGDTaaCBh9Wwauu42fVGq10W3fABtzCZHa
yAXzYujAkZJa1fDci7dKQL6IjFRHQrZk44rdht6AQM1tDmACXQz0yBYDChi75eyO
Xws5cOYN4WcYbhFb0EPmRBRSLDAbAvuGAodNMFFUEr06ukmJdYW1hmWtkiZTaK+Y
yUBM+GFb1Z/M7laRFTsGl5Mvw+Mz3PwLthwn0PHE9+zyNtTnqjIRcyZjCGNe1qlr
xB8DsaXKt/dMU59gYhj/jiAc4LxJJ5cv3F5tAamIPdSIeAmIrAksLnK9e6vIabdR
V/A27gxfLj5Ov1bubAzYBAENjwHwtJtCMMf6oaRzwp8CkdiNgRV6M4aIyfP7K6ZO
GwjNDMBhreAtR5mCwxYERZ3oSYKAZSdq2dWeFv5u75fwwjgTn9mEhn0/ZieyIvfk
IE5F60fc1DNKdgVeOv/cLrbdncNVomLSaNmhWlrvgq6cG+k5h9v8FEabJTAQGXw+
oJGgXfj7UCuTDfGNwLNOKdhLnU6AXfDXnwV2Blik9/gfAzjQ5bkHz0rAbmbq/ejV
PFN6iFjQmrjj9YFDcs2ObRVYeEDYDFiIh3FXc2PwhpaQhy2E24769KL8M0nA208c
FoLhjVL8Meuy75GXm/NZOOEMlVz85/iOBZsd2RObIhJdtFCGjciRdfRcO+W/LCrY
TuhwPQ1qi7HUgPkH4g80LW+7uHKjU6XBuvx3curbE5PAqJ8R9nNmZfeRlryGUCoK
lN3se2Y3f9iiUiTlskHJ0zPnq5ZAt/xf7lCgDRUbIDLH1RGVxPIIA4klYAjVOm9T
GWZaSIbIFoE3avrOffU0O75OPf+HHEyNrXUnt6HThRyyVwmSGEKLaFcNoCzDUqB5
NFyqVjlLccCShmPMVRFgl4DXGEWvT0KV/D1L8WKijEYvI/fzmUIRbdtx1bbqo8RT
fq5lQvPo7C47+gxl70iIEYiFp3apjFrRbjchKrexcCbI/X+zwj2tU1PQEJ0OgYzx
NtIsgzlxhV236GX6F0moxhBw7IqhFdXQVpTzBanJzTmzbp/2NgpdWcn7QWPpVp0R
ZFYRTrHu8bz9ylsSyogj5HvZXK5bqdY0Oi8gF0fohcsH3hkwfeZsS3pN55+yLzSL
5lBfb+pEdmoZItAzJBI7ZUJg5kOxqQ3k6GlEpBSOxTk6xFxOZGjmDAVk3k7FYo9a
2/5mdepydDdQbGR2VQ+zxAZipoBfFAQj4dhfyczIrLwZW0+mEPh2iyVFQVxBrYRY
bo5GjRb01OHLnCo4cJb9cjdL5mtgrlciwQgrMkl7Uv63WitqdxA6W5vRlYxEIrtK
iPdhxaRnX1TVxLfREvDPIQ0/R+IXB8OoeisNxmGB6HpArG7tDyLNN5cI1ncQfvdp
X2ZtWjYuN3v4IC5nUsLgz6gfj0dHb3Lh/ibzwg3xn2QFLrmFpPC45CRSU1nuoLYg
rkKcbEKMFnuILupfTjFpo8Qti8JhnikZ6pI35h9fzo2URJTpMswTPZ4bDScMt2eM
iC4Ud+gGq0PZUD8UFeFq55TVGXuBDKiK7+jC2gfuofx5+xYB68oqTu9gm+dVbybC
kkAw98eIVbKqhNL+lPGhbeIjKWmdG1vd4crCqniq7fjYfBNMBt+lOYKXinsJqexG
C9Bk+pc7hasA46BF8Iqw0Y/TSHCNcFLqJj4Def4H+M8ldrCP/9G5otm3jmh77G41
G3slQBP9mGwhS7YcLjezNKIt3LngqrRX42M+nJntmuTq8lJyaF6X58y6+Pwsgyig
Ul+ZkJkTir3YzCQsgkvlv/QA3avkg9pz/Ey6lCZdlTzYXmrKvEvVJnvgZh15JIAm
PXyrW1htgjcLtZMQ+zHqJlXGcIZopn6d6G3g7xg6W7EI2J9bdZcY24PkjpOES1uZ
vf8MXvMp2YvHcqRBmmuIoewnNS3msQ0M+7oA2PjB5CM2FVGGoBx7WcP2iRS/DUbI
lDr6feypKyzULYHTVapq5VIyMJWHWAhE/Xb/7BvXkD5SrW6zECy4h/pG1Sd8IxN1
CkZ1XOX/UbhOV4Qn9/DcA8EQi18mETrRxqnX6rBRYxnlAjjRB4uhu5Ha3UmqwCb4
bI65K6P6NZ2mDlmYW2cEnh01y5oUaop3b8dV1PPynjy8zypoEy0PlGpDyN/oYk3D
C2HG/cmrTCnUtcoSTcEeN2UsRqFFIFdHkPX6jHyEbwJLnweCjKyqJaAACPZjQAFl
ymXUSeYCFpS9ZSyp1MIFsah/j93t1eLEyqadoHc1eVVWBFN0MrIpTzndeW3hIaWB
bBHCe92z7I89h9rRuamH+NRmXF2xJ84QyCjnl8t/zOijZCse9zdUzEjwoFhOGXCf
YNdWbPi6I1oIYv4LXqyuogn9HyEXUpIauis9pEGIzetaMTndIT9P3vFhDZic+2TS
g9MM95sZEtWwPjp86ZXImtoCFekti4tRckuEXL0jxNzS+6qnahRq9s89dHG5OBYB
L9qNUAc8zd/iFEtHUWOhox4JrZwIfifgz/Bqr/vA9AN9o3FruduoxkBO6y0xERYV
Acks6iFZ4FURhT2o1K2fHuuc8C5C4LLRLggGxB7Cva14aHGLwPIeDGn8dG69WSax
eICUg8b9hZ83Q6KY3yWQHjf+YGtMC4vaJcPamvp3yG6cRP4K8a4Qqa+kAdTEDWoO
zLcGuJJBo/XREc5umUhFQ0XvllGT1ra76FBSBwbdVNJe/DWtHB8y9Ivhcy+RZL+/
6hLy4OboPgBc7PZxwFQ3c6VbvdGJOzX5yPFIReYr0QsVb+7FvbISWDs5v3ypub4d
JQZcCKdXdIzKzl33e2WoVvFt4G+6ZHBgZJRE78nUFDR893BI/pIAJjsOYcClWtBE
mX2Yg9QwuRP0nBS0ngfN5oKbCeqjgGB9/so2afItf0s/HKwKSLVwO1FDgPRjRnln
hcgV/zOgStQMuOUD45SJ4HR6Iz05bE5Lye/BUbTibuQwNm8b6bAAFLt2IFEIp3Tj
QTX4SrslYPJtElE80/CLE1bhLCiHzywLmBdt3So5rtMmfRgTwGYnXjKTr8hBUfKO
lBLdd9rJBY8fWzTASRdp0uY7yL4YkQoVbevnXzVPQ1+bscMdOowQ1IHomc5ot25Z
VKgOG4fu/yaob6DPR9WPWQz3Z5ctrrrbaH2R23Jsb/cDN7dur9b+lsVG6iQZQjBd
4ChLoQ2lCyTtQI2i6PYJ9qh/I8xVhnkzM5TWeOFNd+48d17XhVOFG2/i7BAiPhCU
7lt8gnex8Sm+oEOeWK50GK6kll+7gRrDGe0H0jsiATAsiFssOm1iuAq9QLENjCmn
tl+GaIP7lXjyMZQbI223qddCnAUgS94aJwRBKQ82doRc5mPHqlWu8ItxZKe6W4R2
azDN1G6eJasMDEise17XuFPHbXFV2FIxLCNUC4Q2qiElXs7vp9QN/1sv/br7gmfF
rwaRA6VCfhTLSAePY0CDx+r+dk7yVwXyiRI52Wm0ICFX8KLyXacGCTIlR+WnPkzr
PoKu8gO4dSmjhHORGuHrq51wDaIchkJlPSSFfkZzVoLx50KoJjyy7PuTDOUkz4iE
k+e0rRkUHgrA0xZUmtvFXz61UsVYMdAcZxju1U7SsuNXu/VzOE900p3OuMwgAq0y
GO3EWMyoBDYUnQDo1beHAJuxQr3ZfS/bUKoEjfH7chFKDt1Q9ywNzyKb7bLusMng
HJ+IgTPhdTkrhuYfGwtbX2GbAGQjmGMZK1MpD28s/1tfovBunntRvqA5wLI0r41Q
T6uOkB3AMQUDR5waT+kM6DoutR7ub2ANPAk57+PhIdBrlEE7OcHMZ9mfZTZTF8jT
QwUiudMwgziunAhihQVAwLpkcKyVizhmD9T459IHjsI9/l5vOptvt6gXtQ8H1jN6
oCFFcn6u0zoeKRI1sgLJS4C5KVKgDz7icIr9wgJ+qMF7dWHgODyT2nGXiRzcSADo
6pMYNc75caCbX0yd/ROxCqOZka+a5ucSG7axOuBjwTMKzGIqABY4lStondcmiWxP
dEhAln4iMrWwBTTv75icVZ/GcpWKceMHdNhp/y/BiBN1nLA25a+vMvqwnujatnZq
SjDuogIP0QtYUY6ihi/bQlznSl7zH4SFk0gm8drpYWjZOWfLp58uBq8RZTHYth5w
Faaxb68kXFZ+hWUYu9tT0gGUa+pGQylM+rRv0ZtkEBT9oAntp6cyc3z39OjzzldJ
bU/4AjNSQ7dqIzcSgDRdg+c5UCh1mwLob+NhT5JpoUBYSL0zUwZh8Ar76Kc/20Pj
l69VQtwGMcmJ7GXRmvc+I9AsWq4MAa3PaJ46cp2yvDZr2ZEsYjmhz6Uz/SokC5Zn
bdXUx2MUvNrEp5WiIkoudYoPWs66pizo9QWRgWQhpS5gsTbNiunF9OUW5Fhbz9PA
KWUT/NCJYZLxt56i2EwmX8WTANZ/zOi3yhdsvGRX51ZueU2mxu2bupmFCENleZui
W0qUX/IgyWRO2cJVlBrdBt+JdIAvvh2igoXdIw5zjy4xCyxfKUeczb1eeZdZeRPf
O9873cjZsWIjhnBA8msqDfguhZMOaq0M/jEba/PE+wT4kj+m7c1eCSof8aqPx6tg
2iqwuMYPqDPrY4kZAXIGlT5nGP2UBlD3lsCPRJxlpteQX6YSku9RZMwqVD4muFv7
/rCipXtA6FM72zYudCOUxYX9C1tpiT4U6GyOo70ep8SrEkfoSeBw4QWJYdfQDyKv
4MEQ28LHRkha5b0jTNXXm15YmNBHVzQD7vSGZuEPek0s9btGPYExd0ybm0glihOW
kj2niQmwvLbBP2PTffqYhS/KjVg5BGdmj2XBJzdQb+Z61frRjFFHLW0k8DKQC+QG
xNBNSs2NnfJ7eojiYg6BPFD+YpQIgmOCG+N5wG/C5lurAHTORmLHiLFCQUCSi2dQ
+7weHtrHCdhqh6nTSe10TNMLlBeK8vx+mhRmoxoD5iz54gNtT2tIjH81C7O5HIgV
G703ygKyzTfx2TiTgX5knMXmPj27/TbHjNTgBZYGBWtbVP1iN9Oq3w3h3GDskqNi
zzbTN/M0DtJcyKotfpQSYsHg1IxtPYuwYTNoPcOQvXHeAB1xVG8T2Y0/LPfjk3zP
IprA8PzJjvYicITaxdpep27+ijrpvWGfyDOxWBN8PA4OsJkqRF/1mrt6b3goJ65f
WObz1qjFlROKPa2/OMpGrJX6jyhb+SKPo8KD5Z7b6c4iygVCa5Cytjf3cEAEUJyG
8bNjyLyVVuHGh1cikqFEJcQKTuyWT5sN9JxlIb8cpVTFb2LHwrlKGU300iZJ1RLg
Ef9hOsBnkFNrWvw4M4/cwUywzjWhrYbF2F9FKRyjMlhCfXMh6CgwsvBnSnHWeH2x
Vuq1WSVjYk+HWUg74aPHptRi/Yp39YAE4uxXoZKiiUZ61Sl0Xo8igUg/w3HN2b8P
WxHJzy77uAwp+Gqlm67of7IehiDHtaoMZEU3wIcVr9TkrV/rcieqYIYh0PRj3guD
HIkUAgGq3wBFdcwO4jebCVumdYo9sYj3VX9bxQ8q2scxxJMF7bug+qBmnr8OZpZI
du1w/RANbTx7bHwxrO0QSwWb+xoT6k77eiUum9wPkDWhik+KpEKMmG0BP6P3GLrD
PmISDuZmv7UTr5PymcBfqMmqkMl5KSajawRddCeiWSjhg+K8NLS8LK9+KNEQ4gyG
QUI2/PswO9ygSs0lGOqUAg0Fa4q9WiCh1ZbwTNNWkpuDk3DRzoL4SdrIZPAuhs8Z
foiOl8BVUcWB7keQiMyd9SNznFSBKvzoibZA7Dj6Pi6ZX+lz04rdshuUtc/iOsM3
vGDdcZk4o2ZHd3ZqFhRhvRPWbC9Ig5ahJqkbMpQAzWfFDNLkSvWK6okY0LJPZdSZ
iso8kpuXA11h0mO+Wnrp9CyZrl5c9Bg6vGRZevrx0WsgnQ80MM6JdQ0axBC5e4SF
v+PnjFC1wJakAomLKr/FV5wMhed8CMKgk0Pdl9BI3zalpGWqTZODHIDbyW/OKOrw
UzFI7sKQWOJ3EEvzW85TJdoHpQ4HwRkGC4OEv8AdN/Uxfqgt6FMObUc2vq8PS8jz
5QrTU9G6Y310VdOsGhS2pA1GbnmuT2wT/jxYALKSaRawgxkb5zAYhgxIdXBo5Hzd
idMU4BNPdIGDoUKnn7+5pA4ihWNUDjyJp9c3tkpWufetAGT7pV1bawSsxTzNQgsp
vHldqVslVC7QQbIAecbIbkFig+gIc3+BCQXQV911aDJHlggEqXl6ZyeKZ9D0DgUI
Zdo49BfAR1EDI+JMK0HWphDMCGgkKEpLgaYDywEcrU1eKGSpwqivFs11zuAvm0lA
vz+b4V4KeGabv+b7wx+zGTBJv3T6vc5SxvNfYLQU78a5IFamX7FCzzL36v7nJIWB
iNj2y7SDUxF6y3ycayyNQUH7EZJG/B0ax1DRK3OuJIsRTjZuvbOqtVw5xt4/PmIY
S4LkQWYlZr6Tm9P7lJOicC9bXgjrtXLuo1oHX6C9ZIbMEeXd2eO4W19IlFc5bqsT
Yme+mQmM5jhrxvhNeTlYkkZYGyan8fQrP71x2gONc10rCoQ4hIbATfNCYuTH4/sy
3nAibEMEkXIgeM3/JE7LdbLXMPXnI/kdCVjK4WWVDaTcOi8azVr2BYB/Ntdu5rT+
cKCGmYnBKfSxFqeeSPwYCDp9tKjVcURpJLgYEnALmixwyZSXGjugMo5meGe1Ra+5
oDkeybRSaobSd1vukIOLsGKAi2Wo5+VDXA2vomPln8+y1lpTmz2hPZpFd5G7trCM
6guOcXB3GrbnKb4NpiSH+8SyPwCg/7Qr8tFOUdmQPP1qmqFp3fTsdnrrx9+iybnf
vDN8Nn1mKTdZxQtYJCPli05E+UEoX/53C6AgOq9/WKSyFs5ql6NpzavM3zzjZEeR
ZI9YSs53Fv0xZVDiLmXSAf6a7qHExjXPsFzeYMM+J9O2QG4Pw61Cq8vcXkwhrul4
uboJA3ArkiQCLrHexHL7zrArHgyf9oRZ+fYCBIrZjOZ0qx6nKHh71yOEW7a1JfWr
3rgI7jEnJBu3NUtUqnQVdk7EuF5pPWEzivRFUQOR3npdFqytlEvS4Qj3fWVn96Pp
xsWtMhp8c01ZtJABsJbaHsra/3n5KqjeBt5omArWJBbXxCVRfwuv6wIEK26o31Pv
ddw42LOpsQeDeI5kdVtTodgAFQaOw8Igs4We4CVsjx+WLTGeSCdVsEvEYvsZDvcu
si2J0Q7350ayxvKsP6XRxghoKIpJ/P1wUzJ/sJeUM5l0BY8z6ofMCKaic8KqKBCg
3Q0taHN1u4fqXSLg6CvWYOcD8gFUs+OJyfV6NhzpOPx7e42M3sI835yQRDI80Cyx
bIHzhM+t20Sqb2nWkdwFVQMq/+i6Cc9KY/DuQhNvOdCyz4SV3XiMzqQhXq7hGdny
FNtCnFBx+STotl7oLb/1ADMnj13GdQLJ9NtAgCzIZ3QeNq4J/TtkIkQUuA+DHUvT
KaQzDmDH67ltWBU6jIFqlQ2ADUJsMoIdghdcD8wIJovGZqLjA53ErBfC0aGLiQnc
2NuT3r/Akowj9YGUuUKaFbf2fYTYyO+NLDkHYHtJ7xu3OQt8kPNXv54sKRU6f0+0
Rp69fZ6WdDRjMwKcUFDn57nqwYbst5NdaqIyFMonsJTQYt85V93jR37NiQiwK+yX
TyqxweGaUy3u2Ds6nITTBTif+5CKoiN/dgZ01Kk00JYDFgMf7iycINQdWwFngZr6
hwS4pVThhtmtczskRohaiObrlyiKqPMnGHT34DBpL28CcGDs0XsMSZCvxGgxy+3R
gqOi0a2/CKbZsEoVfIVTH7GHCbpiaG+Q3jxaLO3b9AG4kj9AEg8mv50PZgF4EaBm
JDIKiB3bAxNGKTBQ9Ll139RmIKHGmRpNjWybW9BvCrJcB+7C3NDK5Bta2rxyXqt7
KoxSQF9e2juN7rUl6UoIa2Zzq9MVHnpQxMc5Q5CJ7eMGL8P74JPFCd/It6/v6FQK
uG2a4uWmF0jWb1HPowW5GOoXT47vEmyl5wqJUj2afEMjdgXgVwOQwpCPU8e4LqOt
JLYQbEhBMknURgZR0n1ENUgunnQz5gfr2M3kEMDgYYzZjY0OAMvfGJqLWZ8u5qcU
aHQmdxkFKHYywM63YjyORFdMUE0nb6AdVKYaDdG83R5+nE41GDObPwSJf+BI71sT
SYkcn+IfPnhXJ4M6oZ5fpmSpYJf4UaedyqlY+exsUAM91gyWQkikSRyzrxYTHK4R
WDhATflr7gqYMzv9BBgfz7OxP2d/6Wa2ZioR9z+O0uCuzWhwkXgRYy5ro35NkcM0
KgJbyTVyhrk2M7kPiTfJgq3Zsr4l6SVxH81frssGVOcPipafpcDXmokdKhvpqbf2
R7LcjAeyFMDOvZI8UlHyrryAOtkbsEEhnSjdi4Ztb3CLAEhMmZSsGKJpxWcEc7Ht
zRk7S1vQiaLO+jQXVNlg3Vrjd/O/7oCzIYwktRzz+W6MbnQCj9qYTVO5nvhRVonA
Q2yGLrM1ZP4ftoZ8YJig8lwwd4I7AEif+aGFmTYEcq8CcvvWa0B3/ER91cXr4i9r
VQW8XUpfyxwIi4NmETdS6NpdcxWqi21u86QSqR5I20qRCj2GFGSbebbSJWfEhOQ2
2OQ2DknmS3KbfVP6QWGD77HTyEghuBjVUeDqw0ayBNKyEg1Q/CE6W6bo4uWr+Y6Q
gVTIYTjb0WabXOno7T0cG3PvajWYGy0MiAHNvIexF6X61YCoBczcSGQPeRPMN8IQ
PuSTR1mvsot6My6iGZZqzEZjrmrK5UmgOOwtD8wuGlEYbGV9YHhXQOrok++LA8j/
1F6J7obw4f7aO2+iEA2/C5+Lpz4Jdh7maxqVIIC5vJnkHRJgHeP90QhlgKCmEk/w
enV8mPaX3MYWiPf6uqpcJsXVwpuhudxuuiWTcmhZG712v6q/WxvWR/wQsPMqRErJ
QzysbxxLiqAQNoj2YiLWTwZTJqWsw53jOYKilfDxcSC6Ajz4Iz5PPAoUrkXBnkzE
qGU8run6XsWi1hneFHAlciX1hVNiDirkgLVnI8THQEXzelEXHPdisAGO+iKY7l41
zjD/T8DXmkFi3ySWkaCJc6XIZPrJaGUOSgul+DC/tN6/m02KokaoZQka8QIx6CMk
cgOfVMV2/lolNYPbMQGAh8Q3/fZCihPQLQFN8ItHDoisaR4ahWG/4QhRs7JCbb71
MbyNhnmHjtO/n0eBVmPFY/RW4uVoBK24s+8fCg6SMavoeEIwDGUVUsGvJSVE9bd9
MNSctM5kbjhuSt47jFPdow279PUNbzAisqBrrirFy989nj0zJa9tADXU8cbzGjr9
ngqyRqAQMLSsyaMoBEMjdBSKeoWYL57/A4fldMHKDQuYY0RcStx8wEDoBuc5uW3s
o6LxtI+gsiGpOukZR7iXe0rKCMgof5UFWen77W2qdt8sN8xRZQsqakLybyIUsctH
kSK6Awu6VZ7D93VGCfDXBtfNLzz6MZ1PMfx+fbwqaii8vVMjw9/spbD+4SWs6VbA
zi3LXshNIlf5j+djga1kdKH8KfutZz9S+2AoaV5D7767Uqr0tdV3iu81Qf4YD7fB
AzqpxeiV0hBMc4X+LXKOaFkckN0qCzyAIZRD+tgK9XUsHS2j6+GkYqGoFICPTYXO
S+oLQsC3nAruwmmSD1CC0fmnK0Htoe0hI/0rWv4nUmLY1DmuFYKW7ofTxddakI0Q
USEzbLrxapoH+BgvRMx3dnXImOvi4ootSEJTFobiHdClglamXawntfJvwbjV8jeW
A4W9Jz9dJGfdIC/B9JS4PMs8rfUeJHGr2yE6xMivTFRf4KXdVwpviFKEJyxYTcLd
1peEcbjDl3J8fIH5Fkxegc6tf8I6bvljcO+M9bKRjALy876js30sHPPa5vnKNLMO
UyS7qRv21zCCkWnxPxvDV92L7lkehzPPe+TI5Z7YABJdjtzu/aJ+9R5qqpgskRUz
t5sTlr11Pe+o0zhdOZa2+DXds85aY5NEBPGERhFpY/ieyJu6eXCaI7AqBw3iM83v
LtVmPEPi3BcIrd4wtUajTagO5B7Mx8eAW9o3vO97jrpzz2YFVeWgVY6SBWWfVlGq
rMpkdl7uLTXhkN5FQfd9Oq2xnYn0jBexgAJPa/wrMsb+OcZKWdDL0GX/loARzpoS
9VZImU1p3yEsTaJdH+3OxNVu5JajJctepmV7a+9ulW1ojHAycmuP5o78bS8Ffu/z
rNlG6FzvWCPwuhzCIbNGbsqTJPaq177qAklk3cAY5rl3zJwSU3VoII6cRT4ZhFbG
T+Xa35ObBlNLCQuNBaOU++uiKzK+uX688ka3uN5rxdNdiddr5OhhouH4ciY4HWZB
VPMNQfnrDa5USrU3BKcIhO5YcbJ1ujFDuJKRsT5UkZfkVROtzspIBUhASqq2OP3E
ltIcmSpsvCQwNvfCd9pQDbE/lux9z0v1M8zJ1NwIQhCoiPqjSzGoZ9qIoXLeaXYW
TNjaV9V8eU/O9wAAq1Jwk3IkkkpGqTqGWi74OCsGWM54U7ewP413YySdzbjCQs+Z
+Hwdyd0cBLjMGD+BR2pr9p2X7g0Gs5xmaZKTNtRQaICscKbVseZ2TUrW4+hJYaXg
TZasUFobGTVvu3tsy3x7vb+nhaofQtrdd7mF/d4T5lyHmfWQcKilnuthTRlYodBt
QCn19YxoaaQCtXjoYB/F/CEADRRxTeuK9I6sd3Cpg8QaoMRB44WHVfDetN1/Ql9R
iDQAg4xNs05u0L5lqdajlCLNjQkJl09N8KYoZxntjMsTkzrwQ7IdJhKlRrDaWLEV
1Ppak1Eb1rbmD3EnUMQWYFiO9eLqet2bvBG9wUgGiJAJzQp6s9vQHN0ivPMoEOLv
QGa/hkmCCXpMLc8PbiQoYBVZLYL26QgzMeYb4mzHQmXQsfjwE4UVSKk5fuWHz86O
mvkUgzrIOp18d/yW9R3P2OHWTCgj2PE1hJn9UDKXE9oNj8gOLloZvQxYVn8h/6VK
xyq7zYMgnlbBxl69o7ytDhNZDUWWBZnlsg2tOT68JoMhSP83exvpDoxzgfyGJLHT
FHP8S0JLUrSrjsgp3AHRe6lwInRRihQAoTHHSztVOGlw5EFjsTeTXLsUAovqu3B5
qNJLMWWoVihCnYcEXt1ND/g9MLDLDxVZB7ac7WJiM5RhZe0mR51Fan7jrsWbnlK9
iPgaH/qD1MRHQ3RGq0BsSkDcxASd+9hfCX082CoF2PSpDLXtcTj+ofv9vhsx1ISG
5UnWcE+evc1AjbNxyvgVGjHbtU/TdpprKCeovKJcF6Lw+lN/zPtdjfXoVP82bO//
5kHBpCSmVNlvxZHim7baNCbL69c4nqItyiyCH7p4zox9ZrjE1v6Wc5xSACxh5qYZ
UnkDXEdwUdzGuQkLa2RLcV/7pOAhP+GAl9KnFZt9RCM/jqpyBGbCybglcXh8bwEM
03X8M9Vj0zZQ88jvxqRoP3Dtnt+cmzLdeCi+oltxHudv6hAHYK5N8lH7Smo0zITZ
m/0LOGaWlwWwPAQuRkz5z6QPuQWcxgvBH0050nwN/y34/9tTBk4PFeOJ4HFo+wZG
1T19PQ3zuyX0J5IEb0+OvHjC6i+pXilH+hk7GsGMIUAK20mQn3JBDlbZJ63WCGjq
a+vDdcMJMfzZ1NJCNuE0NGR6tIxufEuOA/GH+w0fcm19AHujWJ4klV5FFpp9IoDI
VBKbzm4vvFjlDBsjjyS6/SWa1d64tc3X4FufqIhFYRq4kGAXr3LOMCG7u9QPLI7P
FYpX/xgEU1raQ7hvSsp786DJ4zegwJkkOC9xEPNE5d6Pbkot4mmd5ParVpxHEeV6
e3b1gLxHhbD9uI6WmIUiwIsDzZDmb2PGRgycwlyLrEgjTD5RguWjleqHRq3Dmo2N
A9thrWP/O+YlksfB18WWhVp5dNezk3f+jmo+1YCQKR+ablLNfH5yVLzuVJk9cfus
+lfolaaILbkMntMlWDFNh9giEUoqMOXQ0GCIJoryV20+4BmywB36NWZltCFRbkXy
KahnJf9j8WKmliBapvhBzSvFVQwXuxXAjQsYUpHfY5jThQM9hZsN87hQOYIEQ9wC
VIpLMj5+YEWC/nx0FewruSRgujtB+gVDFFJB61Ai+y95KMLHmvnMwN83oek3ZIvh
pTOiBVLMqOuJ3Utho4O8aRSRf7sryK7tosabIIqUpYltUIl1uwkW5yTs/fjBCGv+
ee2vtlurqGNiMJ1D/YwLvIsubkqPO2u3NTT5V15t7dH6Fj+IZfGnnJYg2VjjHFeT
edAlcjfppwhuPodfy44WwmHcAsrEWkL44qP6zJsRKWqGxu9BTn00Oe6OgMP7aZyR
rRq08VKE+z+DQ54RCVSP31esJW1kICcRoh2G+zWFe66RdZ+QB1IB6Ia8THe4lATc
+V35BWqb3arkfZFBM0/T89tjhJpEWPCCjvte+RPOmg4uWeetx4yt1kJpByr+yMKp
q8xwmeRVKR6Rwqa30GLXTt+s7MoWIkTHukSxahuyCz1r7DBNIcjR7QZ9Im0oXpia
4+Ldg4UaRanF/qyLAD2G+nUOaBt8Mal3oogPBjaWX1kvibA+luv10J3ckTEKS3ek
vID6Rxh3X8iJJPFgw8HGNkWpvgZTP+7eKs9luu0UFfmMQDh+GHmJ6tYgEcsTnUWk
gRVsEM8x+n+iUXtous0nWKkCba0rsK8uHj4UTdxOZ9ncfm2dRnBLowlRcBUOgx2R
GjV3axewLLddayaCvhisPI9x2a7tZMyzWvRzfg4eKVpD1MP2WbyKoohFxXI423qT
qx4zKKQJ2NMUqL/NUAqX3sneJCv8RtfgOpnv+QbHR4SKB73lZwakiZBzev/w0KGx
ZhOWoDAmYt5hSA6Y9MxOLi4GEhfNe9kjpRPgTe69ELoFbBoBlDkyt/H2Dx2urEyq
zGs5CoIX4/tu/ebMsVbN2ilvCZtYNAS9Aj4jl5tlb+LdkiI6vHukcOOmMdFy3+f0
OSgGGwilbpz03PK7tn0dv/NhVmXgde8euWJlrt4qy6IhN8+A+uQ0w1NJrFsf4QU6
0NwOPiMEb5Hg4LpcC5crDeB4bAhmlfYSIebRF5fBn4b7bW1C6/JsQ0AbELg7/f0f
sajXKevoRg8MZYxVKAX+OFJz/LuxO+W0lxWhj0DQV9Ow3gpy35VScqLlMGnMn120
xc3EbxgqEItOZZCJYEMfvF6ujeYQA7yCHMFsRHp44vCS+YpbdhnkaOvTe7TpRdIK
vhAuLm1xNgXbfr/obikMkP47S8WK1SQZIouLcpWFS9PPXVnWra5TsrcvEBykiVgv
fsJIQfpRwaZOhSLagRvLAGO13AkmbTsbUa5X3UOU+gwzYihfFiqi/ZNvXKX3gYyz
hiApau8iL6AWvHqZqGf47rnXQixsyV9WLWOtpf7cbTBG/8n6PZ0duYmaeDbDdF5W
V0a8SzxF1GjjEFTWtT/qsPaAQJHNB7kJaSNeH+tQgN+DeVbXlH7LeToFe0WOh7B+
ihYkaNn1mtZt6zpZZOHMVh8pucsA0EvSlJn3IW50W7rulFOZxzDRTep5LkZxxUkm
KoNVaeibyH9AJYDW/avbFnfjnYMiZYeMtt5g309Oa5dMMAbUrrZvIt+4J560LCTM
pTIi3eNs4qUTrBFKe44MgIhsMCMhFmKcueRGpIDEJm3rLGq1EKXIetQx0Xi3VPGc
jKt2w+kggd8puY4VRLljgMryD6NLXON795RsaPJ/6Hpelz6Nk1UxPm41zKPSw1UI
YipH7oYpbngJlOg5MqkEuRxkixSmsfYzhh7FJ/su7zZ4YLqiWxK5G02LHeT8dd2l
9X4ZttGbiF5IcACEgRZZqoJG7opRJv57nBk/RvRFDLCx2FBbayPvZVURc0VhE/xG
NnMwplcGqAHi9RBTVnLmHd0He2MeCkwoHQW8wub/e2ctqNHe6InzXUJJE4SCCmgG
PKuTgbSo8JBFEFiHkJtq9tb4VMnA5wDzBCARbBe1+JLZ+CWJbz8Ai2pNyx8cMPva
pZllKicO2K5Of5MJzPiZxapy0iy/3ELKUOTVUdCwQ/+1dal9sSEe2d0l34ElhAxJ
oj1QdmsfD7G/ebwEMv9agnm3UJbINB44qLQKiVi6hdjEgEKRg2U8lHiitD7uGxf4
tH49YdGIaiWKmnkdGQ9WTYmROjcgZYFH4HY3nNQ4J98YulIhIlNf6vTTxrd0js0c
CiXKBkRu5APRNX0J72SZUSzQ+rsSr3ov60qiOJuIciYHCNyOT2C5XwVE+n7eb+HU
Y5ywDVSLhifv5dmTlMlmWtgP7Dn0El4Ibq2ICRMuc40wRL8tMqEB/c83M/6i+iZ7
9X5dCllYLddQ6WJ1WUBJ+rQQTUjDp2ywHEJGHJYhMzd54X9F3f1zrsZ/lutzRd9r
gNUqlU8s9TJFh+eri1oTNB1bLRO9xIUNDMOBSfE+xPh1ilJ6WkeDTGZnliDgv4wF
ye/znhJQYL1Y+w3Zvstbezcy/Y+PoYELA8aZXB/sSN76pJw3C1ufTdfjKEDiYyfZ
huxuiSfDMn2fux6yJQKBSykvE1QIXFx6ZfgiSPooHFE6g+bUmhjmMPzZR9f4kUTV
KM1R4iZ1/q+7gwuCx400Wl0xflp93w69dzVHly74Aknxg2rU9HdtneTNDhsCl07S
wAZ22dL/vOswKAFdMSZGM6BPJa6CROThNKjakpa/8DQtuh+kT5Ml5M9GEOJCqCp8
0RzRa0xniNPbCs7fQ9o4TiX2HRHgt9T1bRhxEQ4scKANdezL5jaawIa/l1n8oSPU
/nMAFznKIu00nqdcu+LecC7eSQAgHc72uFG+MwN+/OjzIhGsotP5jPzN7qeHz3N4
l6dTPPYBsXlv5k0Ilv6kx9Kgc9xjCevmXs0llSoOvL5UCxhHIEUC43+zyjT67MT2
eClneaZKX3E9MDx2CpQQL/HSqaQEqLzrbRDoGFwyxDAw5M/PyDGemUg3N68EHlF3
SRxd5QUw1Oweg+85g9JFZKThTikoKMxNuevlZmb53di6a975idtUBaHQq/gjiH5h
PLID22FsAnFPOvd8iF3oLpsiL+u7HqsDLa/s6N5Xqao/EJkUiynyu40+81Q+2v/F
I2lak3Vs3en1WjqJqmQDpmMkPUbUCj0vJUU30ntMb5FNfl5Y603rFZ7LpFFtzzzC
Phkeve95whlyus3Fu+g2EgCAQNYxOLcnjVEnDJvW5B3kA8YuUhO1znDYR5/UwbbW
l94PJePARD8nKs0YyF9OUE/XJvVnMGmyMiIxt8FsxrzoKE3snJI0Pfl7mkgEYDdZ
10YBemD5qPgh1pz29NQlzvNLC1r5ifgUUJnmo+TeGAdGx+M2/L9uYNe/OXlPLjq6
8omncCMvOgU4P4B57ouDokGK0BAgd1FU6wziu84AH4poFbK6mjEj4T6Hi5GY2MRH
xVBNgSaeSF8zmX/lzfrYjpoD/g83G3dzZeEt/QlvlXS6SvhZVKG+9e8S8As/aX5C
0Pko+PUuAkkVEegG+SqSkUoVh1c18e6GP8Ncr9CtZsj4x/tmAJQMQ/QGQTTfD0Sc
CW7UtJzUUSaY34eHOWv4JwGAg3SJIOHCou3DC29YqDuYNGZ+/M5M2I/fB1sZRDTF
/BMB4p0fT6ojav9L7dYtOOk9lnKnLMgYSKLeCUC7J0ujWN7F4xU9AmYfIiEW77L6
O+wACZug5SxC6VGd0hgAFwW2VVFwSJ5pJGHduqFzoleUWazO9yPmk25qcD/6taLV
q1bdPR+aGSG5Uo0y+RoSIQsxBoMHOBBq30mhtvUTTIUlX5M7oDsNxJ0JE4r/7Wws
tubNxiiqjfDj+Bu79izI66aR3rszOatfyBi8cQoNYtp31TxV+aM/hyb7nXm2DyU2
4TV7Emswi/a5vvIcNqKtT93XzTzm7lqRJ99b8MEZ+XeW/hTRE9m+eS6UkUcLNi2q
ozz5YNIUTmZr5SnJrcqMDKxVCg7ESTMTSm84JlewFKAgUOWo5GTofQz19z6i11U4
wV9djXrTgzq4MxWtk5/vqrh3U3oic+M0dkyujz2+4kYJQDu22Y7ECqlZMo6vRNWz
R/p9j3UJbQRbVT2kZpnp02u+ZOao7pJ27m4RYgYDsKmbGumEtIsiYgp3o5qdH3mL
aXlXyO6EUympaUwSl2JntYUr9XNWGZ0xFjSBdEMOVybpox2P7BQbhpqrTaW37fde
FAUw6VIobH0//8+kYKSJjMmnkJFJJILykuzwSm/+BpNuWroK4E8I3hOQxqbRJ7oS
6s7TtKFqpAUfnuycN0bE2Z7aIwA4s1l8hIqv3Q5abjBLBXIo9hh3+uzwzettDKnU
wCcUuQZjopS/1Y6N06KKKK4G4s6sNqYBCWSl6UDo7UkzlJbNIQDtOcDPblud959N
XJS5f8I3sziyEnCMvHtTRN6+B+bvEXZZSYxck25nckdiZeVnVlD2xvds/A0hgCJ8
eNXQIjk169bBRdgSj5wfZ1IH1B41yglr1TW/7CfOz3t8xdyB/yMeLMVQKYPEn1gb
HFRGugQoDKHyqPtk3I5SF20LRFFTJCLCtpd5nYOGz4HCr5PEz262JoaVjwKAj49A
piZo/9wNY24/R0QvHmw0w9Ygr8qO5md3w9JeCzFiavCltQAdjATeh6EjfLTHPd1/
a9EbGTveEJa0ki2lNbIikE1AsOAmLjRPNTpwRQiYYX0kEgWvgAjIjZN+WmZJfcgq
bWeGq0+45lf7frkQok+lgq6PtWKHUsRAXZL9933DRhKZZdFTD1aLldwWo/kb93sy
tUaLDDOWIq224Efr5GcifK2sglWvx+F+YrwmDBeMq5oC17i/duhu/474sppp6xOG
qNHBSrgJddKV/2zP2sS47R/RLE6zic4bR9mpCwOdzjg+Yrdbx4eperxvu8xJdKhY
78hNxk6H8M2XMmisk7sFMPL1VetpYe9wMz59fRR6P9tt+C5eyKMCWhGUFu9JzLS3
wHbczeSTbg8nez4PAu7mqnCqJ/8yADMswfblWVeYKL7zXrYlRHGrGugdKeHk5gFj
eLnHT7GzPf4eWT3yBJ64O9tkOnJl+xfPz4JAkWJcAROw/kLFxhbKJrRIVCkbJ4x0
Qz4THPSPAb9us3e5DSP+MlRcoaxS2IYDTwBVyk/5HUmd6E1df+379VlBjLAyipTT
yoHK9T67r7EFFhbpW93NYiSrAmTgjLcgAbDZuTtIkFuDAiMPEgbF0CukncaJWN/j
gHzVnU650VS4lMRY5yCweGNtSbBYMSf1gPcyu+zs3w68Qep9rt8c0+oNYnoNsExA
DtQwGYqVX6QDgIgrzg+vlM3Q8WiIc2SXRuz7hehs7SWFU0YJbXSa08iC/asWP1sD
1tB+M6nDl1TT+pdFHWyiwj/Oi+KtpcYpwgqOqsblApdXiJREOgHuxh08jwzZtiJE
5JqkXAIFc+NUvl8pohmoRt5f08zpNIqIh99cmms7Q6d0PZ9AfsMfal0IitVlRE0+
E8payMlrOPawgPfC9lZjyKbSFVigr1xIy3k/DGlu+M3jD4S2P26vHkShfngaIXYY
aBb+19tEB7Qq0Yr4BAVFP3WNiHx9T+uG+c5Xo3YrO/vJGTuwJa+hUSEswfAZWZNz
pu+kBpKqOXnxnEGr8owrToACdSKBdmX6A3aQafX7JSELHPsNzHgxzhVVRNUkFcUP
i5zu50jn6wRg4zDy+S/VIeqP9hsS19VFcn2MXI0TiILO0iBFAMveQvCr8zmB3DPz
GoBZE7Gi9ylyMSmHDH64GCC2zL9oZmFLDoIST9zbnBgbsYzP9z3oJnzcwOmHIE3d
Ooi7I7Z2QYfeB41B2+kVtsYPnyNV7PTM/IKW49zfJLsafvyoYDJrHnngKChU4fpE
rWicmBS1GOkAUVnTSWMqq/iAdO7DzZ+hL/EA2IxLYc1wBW3MjIrljDKkIFYDfK3s
Y7kPEpjc2kKldlLqGymlnzHrsOAYox6NvRcr/Kszgdov+8LO6xAvxpUqr8KL1GHe
ylrDoZAMeNFs4QU9D40ECE8kB1M0eetrN28V3Mc9NHhuEOVndyZ/dyKpKIqD8V8I
seIoNaOvDCj33GDaKnrxQtljXve2boGImAla7TdTOnnWFDGMVoW/repRITwqYLiB
NLK7ch6R4lJvebSC6Py6+gWrPFSWTOBz3QCYMr6I0MW2M76yyx03thQ3ygY7049d
R0PUf3mz29Qwo82t/Fdl3u0N1QMNpJkn+kDEjO5k6VSg+JCPbIVgh9yoAXH+OE0U
QZlw/WV4ZBTs/K0CFKRS1dRPd9G1H89MYrcLHEuG6w5/BuziMujyYFEiQqE8PDHT
SkEoqHnYD1rP7xMM+/5splCP11lf1tp8xyStib6QNBTJAZsUxRoFYBUuD6ijT8Hp
3M1vzcZUtcHyFgtubmSXR8viqFfY5ToQgP+URLE7PWwarbXtLIwLRkeWLJ2IEDas
eAoW6koRQPb99+6Fmmtnr+NcDfK2p4rXQT7p/HMaccDGtgp12riMcmVu5xZ7KxqV
aYjoTBpIJaxxd0NMbbGopHuyHbJscj2aCusBRGRgvaEGNFY5nRuu5Nnl4Zn5MEgs
vuQZjCXLD3tv2GxxvYYTslGwX2+cfaAscyxq+7eseS34pGZeKvXx84UcXT6CA2Av
mi9CaBvNr2BGm7GSP/k5upwfW3j1OEHEgFxfLkbsHs47ovGQUE6MrI+kH2D+ciWc
NpTw9SPGJDVhTDe4bS0c2qwRJzTNvUo0WlmS0uv9htBCFPG0w5aP6/VuDnrGjI7H
oH6fty/z+OqeAoB+QEOm/pA80LtBh1Vh9CyYYVY62cK7F579+HaNOzfayTUdIRsJ
r//HmsJacDXT8BiYTPToyRNafxThQ4tBoiODdozJq4PjtJYAwy90ZEWIg6CwbGTQ
RBzp2D+L7REFzoQO2uTx8cZLvvPQt82ir3V37OOR0BUMJBTq+ivsVBkB7EADRMVf
hUrkAwHTI2a2TC9HFgAxAa9GK7TI0nDy7d42ABG0vLo5YdSpo8bfwf8KFDpIdE9c
i0D6iHcQ8Rs+iu1ahH1ROXMMg+G4i3ST21IM3PC0Ls2HuvwxtmCkw+QLoIjaUPGg
NFd2iJDGlP1htbxyqvgM1Bxw66KGDyl/tJsPS2JD/ws/RiJJoZO7sF49QW6va080
yQiXlbXKGwKC9HDLkMf/6SkvP+w4eDqyugTDHcx4M4soz48Wn4pdTyoXDQwTd+TE
rx9SvkSZoGq+h6iM88irnkSSxbBnwF0Ipl8XI3x63ezhISWW8b+60bgDE8XAqC5T
iIffpYIKyqtZuHWV1XZoTwslZEBHugOA91jDhhTLk+598T5NLLKNrgj3t39sP5hG
GB6pDXIHWkCivIqWJKghYbPXNpC9PlApHilwS9WkSDNMxsLXwmqg54d6dkUkuRAi
XpCNUpq6RYMXXLxRfe0Ddi3MyG6ZWautWe3wtaU41/h1w96ezoZWhLf63MPtPCRV
b7XQxhpRQBW3dgKfQ3QB0G1Dn0aRgs+jIeURereC7m9czG2kfsGQSbhiyGO0hcc7
dJ1KQVjyvL2ru9LUc/CmDg+jw457jQHLfP/frVCZnawsecMIhLPMtC9jEbT1SAqg
cU4Vhox45yMdRFdiqSmshb5n9knSId7eP5VxrEVAD5ojh8R7U8dIi05w//vCF0iL
5rd1hZR7nBTsyHhE7dFsHvR9CeAGA0fwhtiFXiPAB/xjyPJEvTRzidGbr2ZQO7h2
S2xRsF8eHmTfptfEx67OVcZMhnZGVX/itdIvDDn4JhuAxS90XCIaOJ6Zp1sBeH/B
gGYH4yjxglrdxpzCRAmkf40ZXWGozq00N1k3uTmtZhMwIfFknOu3wah35gxSRX1h
pjxqLC1Gd/i7RUjoqiv5QiOltrlMV8NhFYv9u/ydT1SAR75roY4qflkif4zb0mDa
bmZZCVNQlUgbQOE19uYh7uTBR0LQ6D15gkb+50fOrsYBdiCAHbpAt+4Uj/9Mg6q4
6+7Lp8wmg91OHghq1cVofhg0R3Szh6CuCEMrVwRgr2FvsXT72o0StOBPXI9ruk3b
bwceR1StyNX8wzs/tRW9Wek7TTAXSYqntTvhNdjJ2jc8PM3PN2BOVErpZeIuekWO
uRTQXObxmIdLIxr66H62rXjbZZAwAwqkGhVOEypExrd+3R7CXB/kef59t+C3JHHV
eyBxDqwU3ZyxHwbfhT/QvvbtUIdfKvvha8NsdZA9WYLQ1eiIh8LlX6jbGZr6KcMU
lilPcJxjEKNXNFz0kAjRk2pvEWbA/0n5pp8gjeouinScc+TvIGiweVJHUh/cAYxW
WK89HcvhAgnc2dD6gKD3IJqalWMCOToojm9k7pEs11CcHKQ5yI0qKU/iJtqwJ7+z
ffzrKnwpsGlv5XtseVltGjgYEHhs0hsubsJmxYnOXAfbggm3yD9fy1u10RVpm1ha
lF94m3f0+9GS9zXYIiSPmbfR4VXwx0GjCdiqCE9q9d1ZB+wAf4FxZ6NckkOtg66s
M0z91DQsSVGu7I14ZunhTeF2nyIQm5ZCUD2vjF76JSJNklUWrkCOnxcwquWSUXzU
eYQR3kZfEqZ4txp/sYi5oMfI6rcHpZBN30fEA/SWzn/+ZcuFUECjylUv2Yq/DkOi
F3MmkPRcaHRHx85kD+6AU5UBic3fd/nEl2ERTFhIQzFu1N+3wiSnNylP0Z9ln6Y9
0Kt68ld0zHxLeEWVGrmZaw67GEAbCTeRvClAb4ouT58fl5JDhj50/JAyXeGY6eSp
yreP5X8TELngcZqvi6oZ+5eLzIm8i1c1VZIoZHGrZ/e0PQ2WLkBStlOt0s/IuoPA
p9kytgRxTQ500XoxRqLFpwuwyPI97fgRhJJrcj7iVbfo5evT2ZVkT1Z2A16sCHj8
lA9YNzcc+yUCK1CAaGsSHBswMIYr3JsysSFBJMtC4kFXE5qhWRnF/k83sQpqIjVO
UyZKkMT9aySGry0yuObSyOIY7HDREE1tRj3/vR6yuV8Yrum7SOG/vP0sFtcfIFXx
3DRwhfnCtRxk6ZBBF6/eFEspttFtb/+p6sRZAprDl1Ou7SOKgKyX6iBs6VDrD9Wf
lMDsq22pgnZ/hdKAFNHzmxMjbOfqeVZAV+ablXKwuv40E8JLdtk0kwuemKn46yNC
RO4LS40oM5EWpS09vED0dZ5MpKkfByID4jVlpSRvxllm4vFE7xw8Y9MuigVf2SyW
0JaZabAG+kia3r1epHvMmo7n2HfmeYfWep/MExzKai1WrPeBti0UJvMc6Cow+Okz
Q6ZHcR2Fs3VwD1fXfLM5X0v5ZRNs736FjqFsyQS0YDFju2dW5BiQb9NX+p6dYEnJ
srLvATfAzK6Qf2mfBkmWUELO5AMvDk8AH0KuhOjEDT0B1KDmfzedLZvDHGK58ZS7
55enucSm6RsrNU9sv/TrlxqrUocXvK09seqrBJYsGz+KhzT0PqF6wtsPyyq3wtc0
9VflighNQ5GqKkz2PTe2LFylUewT39TVRbgC+XGOGilqS2Fbilp9gnMQMYyW2lzf
beFB5Wn8KI9ufrBrN29fQ6CHKq8WjCmEcEyrq17n1bPu9T00KDVxld/YtrZ7oHWj
RjpouW+5ZXfyMFH5XtvdLhQ1veztQhOx+X2FesORKd+XD20oz/FFZcSU3hhJNLUz
w0wJJAA1Z8xb0sc+KrvECXs2OCnhYMDE7kkUAwq2yCHyoUYdntzHJAtqPHvbkVHC
HDYn4PnbbqGvRQWycj4pP6B2X8DGPGXzRnifAVc34vzaH0KsUUDLcQnHMMR8E9KZ
IuKK6eo/UI7/bUTaxYjjoOXUsUYxdr5UumnHt3CVg9jEh6XnX2lwcHWkapGfJaTm
LCyBaqZupaXi9JVxIcq/3KNRAH1ISYRCq2aWCzWULWcmL/N3iamnZD/My/JwUli9
q34acCGgf27nwu5yKJQpnxwENqqp8yH20hHcqs5Qqt/elSg/X5GYDENCdhTacCdx
e41YhO5xwyCmYyKimWS3gPezPjDgtltU1k+BZFqBdjr91yDNIaFj9smFLHWOP9yl
HK1d6Qm5K7dAXASumC1SgFI9gxdaFkuROVimVwcP0bAhfvALRMXc48Z0B1DnbrkQ
/YiXuWxMTuKe1Sz+sCMu3poAebTjzFc9Lz7q9N4JF87Kzmi/lpDWltBbQWyvMJmG
x3I1juL4hVRhefclCSuJddTrJHiAVDOKPg++tKOv/+7ERnt3HpQT8l78yJV3XwIm
56uQsjuOTHpGBxxrv66ytGzlmwe9helPYHB5gYkNyEoVTXlfMHheGGg2b4mB8W7i
sb1aZypMhQT8OmKkgdOO4OnpUaXMW8eJSokXEr1KxqGDfwWyB4zoyOOSNZoRmsQn
mT7ul1is5s6DhNwcKzIzRWYf4+1bO5jTA0X5zCHQI/0zdG/cIyh1FyIDGyv5JgF+
9CeZk3dDnRd2ejw44+TwzBo6/YPt/YfiG78jC5W8D7CEXkGwIYbStEopc8yo8O+/
3dthhSghbIVvU9infMXeouoS4jOs0W7BC3nzcNW0Id44S5EQiSKXC9rflJ2b6ft2
+ODuNtKhjdgPZL6jW959NMAqXC1l0t8IMskYekLYiZK1sdqldib4TMigX2sF6Np+
v6Dkf9BrI2KmwXkfUnrpbx6Uo8X+8RuulTeEMgXklwQBvvYbrNQ9+0iERhzEOLnf
8ixVH8EoiEUrdz/0+NP/6nrFDXohrfG36m5N/E/qJoj7VSagoxR7K5/rFGa4FFgt
fjanq3D1/x2xkBN1i+d7ZwY/bkHyFh0C+KgIan4lNHXtwiP/lmWucURTEbVbRw8z
2Pdj+ng5QLEVWypuGDGflIjHWsCz/37o9819mjc9fDqZyzg6JZiMQk7m4qh9Se0p
vHRT07XM7Z+p5DUvLdH+5ZwhYg+geqN5uDJvXTcvY8qROpSTVNLjPESmLVbJUdEU
UqnpCVoenTvQ8v3q3Yl0cpQZpUndgvEBbaW1oHf/4+j0HNFO6nHqKoqdmCahb9g/
z/mLIKM/cBxshGCWnY3uUIGecJRptXw3PhsEpIKzfKknaiL/2e9Nv2yOT83+icaJ
YzUC7mPMGYE/qfz+b8FLhoAS7BhFvhjRtUSjaqk2Q/fe3HvDkfXIAqFzksR8WUNV
I802GOVRgtQdE4/b6dWxDUaYdtwkpLTsp+td6r/v57KgglrfFl1Mrm3WR9htTORY
hc8++XGMMGQc2lZfIi4jawU8IB8YAfbgClqbJXgnJaR2laaAHxwLe37nXoR6piW5
a7xoPnmy0zMTfTG4ADQyJt24C278ihqCSkdbPgpG/vR0SXK1UUqOYNBIjrBtg/CE
O/vZvWwagaVTv4IIYEO76ecjLFUR7BGyKQeA+ZYypO5M9mvOoyNVTRI29aZxIJpQ
x2prEeCMQSX1s0YjptJR647Zd8aZ7KcKqyK7U2J5DhVWZs0zlUex3NKPsyXys1vW
b+JxCVUkd5MRZqrXIIIQT1NF2Op2pHCGN7bCHS3TTSjXtB5SGZETPFX+8aAh/j5S
jV25ekBqR8OV8O6dmI3gdEodiWVbYzHO+o69uAZgJKAyd5opk6O7UBUgWJGA5T/u
6U+3enc+GTE4brwk37rjA8FVBnIicHfKA7F2osjBXqcuolDHVTNdpUT0sy9Hjsph
4QkAIfGOOdynSBKvAjIZhfBhsMK1O0gI6drCcT8miiH2n2tJIwqi0Q03ws7CDPbG
r1RSWW2GeBD+pCSvY7/eYk7mQdBnoZn+b+iATcckxlziuC/+sxdI0xFKAbM2Oyi+
0thdo1Tp2YHrtp0krQ4Ws37nKQWFwl3S6SqQTblIfpSVn+48IlW6ruTM7UMApETJ
CNZqcRP3xjWGGbnc/WhlybvJDYFs6BtoF3g1IfVZPZ2brnDimQdXIIryz9U3zCd8
rve025URASwrchUbokqA6jwv+X3RqEgUtNAMUi/3HQlErNaTbC7p6UTLwI7Vxuec
Ax/55O+ElFkWnLlov1DwvN97LA7E4yrPN1+bvMh81QD6WO9O/NNPUoKR90BkvjIE
Lk7dRzFUiwltbt0AAnMlNYsvi4bnYhLobQBihDWDMVPFZ9WU/+7yL/l18bCnNGfO
z73YV09twX/63NfSgqxRzSWZGhQZVIvV6VQjJNPyizQwtpiQJ828abmK+Wa2OShv
4/IuXZijWh+A8GhqKijj9ha5nD4EZn5K04g3OcfgizKexgqY2QW3KDS23Ge/d/KP
+lT0EcSqxJLyKxxQoOjNPqY8lqmnNOjph2cLdXrAoz19u93LMt5kYpk6kCQoRjBD
GFwZW3Zun1oTxjC81Wa5LZIYN9XG3PFg1siFGovJOf76nRdR3nsQH52quf+W+chp
zqjzxSXHggIwBMPQ8x0HcT6dtnw0mIgh1BhNmPt88TkCYemat2j6wil6rFvTxwmv
DqhL4gywvlHSUkF/pMgOyy9cuCKLvryFcPlelMS/UcKUPZWWQ5XLisFSfWWvvCMu
XRwaLXD0cMrMWo41j2JJKVx+U79UfBFaGDEZKopNGLxBdeOwhSZG30PFnFaX0onQ
9cDfOtqiCA7YDnL65UJx8IsN1Xd3d7nt4WNNg/W3fIFPYZfRAW/jNILJMCkECVbj
//4Mvf57P3I1LbiyO/JJFDU2PtVsZE2QLAATLyPdoRkTh5MEDN7libQppuzBdPiX
20lUQeiDnl96pvu5O0BdEAqLj7KT/7Nzl+TvkSqmX5wjj8fbTrb4jeE6cK3Op1Cw
Oa9Tj2VngAFKSrZL8UU/Od/EYvUc/jevx/ySFL9g53db1Q4XUbyhAzBQZbV+fCVT
O2dGZt1gvJNESD7uKZwOc4cD5n2QEeRq/YfQUnMdppZovV3n77X9uCMEqTjzrrfS
SsMwirMZfOVUeiuRus1iJioNj2l6G2P/HarRWCS0diwGzwcS6+BoX22cN3RKypC4
ULnC9fTQqYPvn8UKbkaE929vGphNmdMo/4w4nJS4nokzpdU8lArWyFLiP50SWTYc
zHgiiPmBlJOM4NBuZ3TrRK2YMXo5zEXihIMvGVgg6PHcYKCcJ4/YJdt3w2Y6C8q2
l/YfPCt4kVn7gbsMAaI5gIwobD9Ohse/hc8cEzZubzJGT/Bo3ufZjbYyqr63LY5q
uuLPcbb9H/pYqJNv6wEzuQ9owueMV78qJBfLKA3anmg5WqbcD1R8K+ABRYMKr/J+
Nj2b0gST/OkkUHxb4BEUkGZ2nZYm6nt7gcYnSPfA4wVFVydfiv6v/1DC3Swiahzz
uivOEFHEOKA2ImFBpmp+EfevCMwJ54oYdiv1hxpsg+7c05kjM4z3WxuFevvhU7za
OrSlfPH47k78zGpMad5HrdGB6bOtPOzNBmPPBwaWcYE61pfItRBHTxZoOKfBFqsr
++Qi4o82xV3oCtUtmzcEvi3lvlqx9zvbQuccNSx1GVVxteuVkvcbxWMUvc6yuRFz
0LdhQ0MlyEF75bkF4G741L7Jc9NtV002jez/S7fhOJh0CTlf7wvZqfqwM+kQs28V
LkIjUow+1inQ1npiQzukC9KYxwxci327PqvsBGLOv1ar8p2aXNj/lL6rNCOt9vXN
msUDtQYuaSXBmK+wodF0wxsElwA0FRAnOQAM4nC55LA1uv/kTrgrCpf/3UI1R9/u
mIfSkQ09I9NTeCaSi5j1d97jtO7E2OuJnbh25fmz8fQCvJ9Yth0BT3oi573n6MBW
l/aLUXaIXCNVO7qzLEG8hQnWgVKugk5RCWB9FObwHygpb9NgUzHwnnnMp2Pm/g2D
NH1Fv7HKiQdYFteXCKOqDUUk/HKlE/JcP04lhIjlAsMbiWUtT47IRUQGSEtmS4LW
1GEoDZLdxXV8mpTyOksh6PjtHsO0V1wkribdC+jJVbrixeqsFlLtfYEPkmdb2xo3
BBWQiqFXXN4l4P3zogyZ7zmuFwVOQVxeZ/xp8+TRP/CH8bJyp6SScu9g6wb/8xGJ
VIDNBKQ+hnq5pqqCgwGloZM9w9pHb/9qFbqpjSWVb06ZG9WWJLIOh+UAKgJdPpL9
lQyCdOWjZHoOViXqmyEAKsm0DiJEN1PG5hz2YUNJD9wQPSWBAUnzyZS9eY/3x/n8
D96nL26dJbvfxJHwx+5HOVf6J3XQ49wB8ys5w7D8Ab3GOOpVWcAnGlOdn6rohcU+
XKA3urc9VhUqH9wQ20hZyewtmHibfQB4mcpYzDpknMCTjW7fQS14KZfqgRDlGCOs
b9hBwcq6KWNrCzYUo5FNSmm+pYziZAlyImmGV24xPKISbYZOTKU7jVW4e0I6pTq9
zNFqkug2fJeQQkWbQzZJ+NoLkemARB6PBSvLzAqnic3oTmuoJvQUOXz+A8v1S74u
sSnqbRIHjA6NLy+gmI5iLT3fU3atV89nCwg6+HzDpDRowVcNjl7mp11b+zzw7qfG
bxflNJ7oAHOL6labzoSAWD5510VCiHPiRY7cWeIiHXyEyCoMWkktlJN4bz4Hl+C/
1L0RGOdkM+up7F5A6E+IrwEkDViGzOJnhbCQ9zY6nK8m1t8FOQieD6JIYy05wsKz
Z1idVXIMko/Rcc950DhlcNp1/CgQMhAxuVpaKP4nwuv4TCqc+9V6s9PEKc0CDOpX
HFbB+SnJRM8h+StrahLwEovyJTtQz1jA8FkacAcRt7XbqKYsnPzaZf1HiWFJKFb+
cpCCFhPOy64Do2B0q4NlIG7BSFKcCUJof8MpTnmmPoHPaith+7ZS+p8G6EeH5rVp
3ghQJWhK4wkHg5MtxjO7fsDhnz8e3wcdSwjxb8Y0QsF9upG89q5Jq16XXV3il39K
aJQyoa7cnmL5JAgY6fS+16tsquPcqZbDWn6723QbfsJ1Wguf5dG6rw0r2XOUqrk+
JzOu89b872r41E6UeH+DGSF8vpIu8noyMoWcF79mFzUkCreqzCbZlKBavZA3Y1NK
6PEcMG8O9ADFfjeulB4fiWpf8dQzStDJBdMmMSgCkRQYoFj/MNAMidb4HvLiWLlz
9VuST0HidVT89iqQGZVE3zD1FRXko37Og9GN2kA8oAMiiDoA5oUNKlgIbMaPjgF+
uWUuPE1qd8bqmZd+QFtVLXf2Xtn05pndtMSxbDzJs/ctSYj1GiH8UZR/BP1B2WsJ
lr5tKAk6ZAGNN1tWiz3hm6Z/BZNaIlBgtmmqwDjRt2ThoJ2uL0XCOb7jGwa7ah8/
orOo6zuo9xXMl+641z6Ae0yf1kVOpfWZaOyDnNaJRY3+S2xE5w0dByKZY91WxYko
O2XTm2gnEV2R+NyrWX7hGFRSac7xwOlk5ksi59Jdli1w+uaQfOdqazozINnnDsC0
jR8FFMbAObxGb0lji1CuqQhQzhhDiv+N9Kd6HIVcsnklQsH1BwPy6zlpzNLg8v7E
BgCgg+REbuRM9DaAqnOoxdUA2VSACqDpofwDMrdHD+/PHvTpt1G0m85u5yldhYkG
jWaiF1UB4D4XXIHtRdM2G/k2I6T0cJ0u4HbmdziQWVtyPxqn57hb3rL/DFmTm3jP
g8lUKaYaaAD8JNOnPKaMuFFXs4/FtcGbET8LJdfb90LoOGolqGP/Ye/mK0vOJ9BQ
ELkPqT7AgPXNFtCj06uiGTVan2/4NvB4Wd8ECrk8mD7pt9bKs3qazyxcQZrpW5oz
icDBsvDjin0m014zV2LLY7NtQBoSLzc/NTYb0Q3rqfs7Trn1PPf5tGC8cc5YFoFt
x9U/0dQ8lVNZ1CWpM67aIOuKQ19FFdG/iYBAHhT4S48VcOPRM/+mSPW8+kdCkcu2
ScQt6Xy99t+gbs4ZZiWVWvhlpgFgTgu1s4NtwMHEBJ/hXE8h/Veu4tpgOH9Bne98
O4rsYe4b41dHszUgFRGYl5x0ylr9K0dpE/fFAlvZHrHwDKuwx4XmLXUrC86RVqQJ
dHczKYY/iX6zH01owCDY5u44U8Z3V/kEGz6BcRMlU2x67OQ0LMEzWdYIjx5Mm0yx
wdWd9IExc5iyBUdxojFTPAcEWfGze8yVtPP/yS1hZWzS+/L7tcAJLbXF+GAXQ1nZ
zki92pN+lULKuSBI1e5qXVhJXRW//Yq3WR1oIcmZMZ6nqfh0bwiztCsw87ZPxtpx
bnV5C6pB4+BhsjSq3Gmy+x7Wu2koKW5TF3sCAylsDCzXQw6bgtObfqMxRWTa9zNz
blJU8DORfy8Qu6uaryWnbeuyBFVSWZclYwn5eP2ZhiWpI84JlkAxJ94slOM0eOd/
e/w0nBO2nXdgDAWJDo32zdkuSlHk7hHkdbugsAnZhZt+W7RHac/pwgrwuJRy2qVZ
JWtc+IMwGYNvdAiu5FrDXKn2qH7OZo6fl9pMgvEhz5DwcbXdWPf//os0g9jMzrOw
MCyYEp10SogI7k0acrEWG9a3gF4sjpBvmBAD4rFXp96pcLmrzbovaJk7lwWn7osg
N4+WfeUktNob1qmlOm3QRohY5Du4EuzcX3UEYOPNjYTlzrJc1ijw8hqvbeJgDkhk
n2YJ10xdQa2Vb97TzOeO+KrbNO1IgCugX6IY6lR7g8pT6IqxmfNmotxVId91J18k
SOicujSgRiLyosZuD/I2bLjhef09xYkbNx2fOrK51IZSuMbao7kauy8NaouvcEqP
S0kTcExZqE4MoloelfzPJBt4J45XBNQULjeiGITKU1qnmUt9zJu9DARIyvoabxXn
Sm2synIeOMGhhlofOVW5W/iBMWDMGtqT1hzfppTz2YPoTaebU05kfdvJ17CTqCJF
q+TeWgMIQ1SNIWEL/LHVaHbGYfpxO733/c8yc6b2swlqPPhnfLmVwysg5SS3buRj
byXvTEytsFPmLEOkh+98OUCx3H1NS7j6kxC8nzJjMCu0wMw+eA3arHaFKX2PeKpr
cy/0mIkRygv20bS2PW14pjOd1svRMJq7S3HWgA1rHDO8C4h/Wj6vhahjeI7r22fd
u0h/oCMWYa43+SbAU9w+x7Fz13pbJjEdMls/yJ3DUg/ZOx1qZj9Vt+7As1+fgqv+
rg9lQQPROil9QaYnaVVtFqmzFcO/N5cHqBl+sccOef66ognyp+ZMLmseH0f3BYLh
W2hBZnLIjgsjGUlkSbfLbtsE9C6E9xNeEBfG50mLZrVUqvfFat/63LFiJfdfXLPX
hlIAvn5y8oUpA3dd1Rn69EdFl0OwpbExgt/OT4j+a/1jleNV2HFItPk+aIeK+pJS
kU0UrmPA/3v3HrYT+UOrLanKQNxL0veW2hkkhczSJSYMMVtV+K1qnVclQmKcQAik
7NNNQPwPWsSA1NtRWb7X81iufZEMNSaf/K4DLmI63y5VYhWciJWeXrYjkOjCytjm
Pp4aYatCVq9/02hA5fJfMOvv+4wY6jHCSWvqUw5Hxx7VhYAPLg6O23pT3m9xnK9C
Pr6V+SPGejNTBIAqHL6gyvhdpkMF/hcubPa5wObheCSGR75G5ns3CWZuEQ4h9xpp
lRRUjdReSvAH8lwTkyBs8LVNmzv59SBKxSXa3QDeU1YaYgOZEcZ7XGZGLrTXBT1H
u3Z55prGF3+hcbWpTYasP+dE832SWnSf7AaCD2kouvfcQsR3ox7I5yqU35n6s6a8
4j6LZZJ/BR2iy9+8ET9Ia51htIAbjDDe77rN2qSB9SruJSqKS8eloZDYzEy4Qphy
vjHvepd3RgZ0Tkl7BwU8705QC86Ouej20bWkSYDMBvgfqhp9beSZkTc7WmJclvwW
spd32oN2sPD8A0iq3HfgyxVFtcJgnpaFUKR8PYYotHWCTHoqFWY7FJva0fZIa6gS
0tT7FBvp39iHxQILgxlUZuUqjt08YWnYP6prASsNT/LKdfU5JFZ2KKGhenlCi7Ta
JeEmD5/K7H1/wUhMALPTBvl9+kGXtmdO4KZ73z0uVLob+yD6oKR3pmcan0aidPmL
YVOtnhNybNmIhtG8LA6MUs0dUPS6GDOwtv6o4k6pDjcvcENg2+3t+WKTE3HlN4iA
St79ITdIIoQh4H9Bq8bKaEdh8t4j7oTg9O+PhV4A1Sb2c8xY0PC1y9O3ZYVuNCn2
50ZKaHUq+DTfiTj7v3X7Q5rq4HrJh5P8CPc2feIuVBnpuh2gdXag9MXyGyAj3vY4
OBoqUgdu+a3ru84ZbR7vGQl6D9fgl49Ut7tynm04d2r4PfwZprciEt7jC20ked7w
9j8jYbpbMf5HxznSHIGcUiRmGwYzwVIWjXZXHEvGsYZ1rj1mOr2Yr9yhQeOqVRrX
xNnxLgDzwZekbEp4og5AEdyJVF+hGJdRvzAQhJY560FNe0suoRknEi/3jj5AqDCK
2g5WBkHQd3biFceZxwzk2nwCOb2y3iVFg5xlRKQE5POujtSbQ+XFXfvJctCs3WTN
wMHmekYUXJO69AQUPCWwvHMGYQCKPQuz4/t85mQN6415W6wIeNZ+2awByMVJ3TSi
NZ/Ap12Fauc04clFeI6RHn44rTG3eW7aTMJfvO1X4xqsBwkYPGVhhF4TtyL4lfLx
SpJFT5frP/gNVC4pkiBdikCVG9Us/vtCxnNZSFKg6+2laWVOLlsafVOH3hXBGxlN
p/B1Ty+7VZKE88vDrRz0fY1L5vlcazg6E37S/DN5EDuvkpxo7TeCXhFK97ZkmPKI
TTeOyxQXKgNGo8ctBoCcxLQrLHrJGHLcTHcxDVS6olKYQ/Id7vqdH8DxJc4BTUZu
MgAZiuJ3zgaiGeTO932qPe654EVo1AvyajuItnhVaMSLmLdzkYmWz7hAKEjTiSBi
j6EWqaitTJ5+Tw14IImadI/MxPfDdqJZ6jOiUYn6KL6R5p1s94Oo/g1DoJ+fuseY
MYUhyWaj4nOyz3W7Qw2oTt2odV/tDgZg9sgACtEzbIvYybTw4AZV4JOp2owxdgHO
MiLoe71OoGpUW4HIDHLHb9LW0jZ4qi5uEAdCeawRlt4SPTDM4JWANFs+JzqPN68S
NATp3iTQf6JUde1F1iNU/nQxHk10OdJCbRaOZs9lzxrpN67F9uYujXdvNjK5JWi4
JZfGhWqNhcsEGaFZ6YUTZRZh1Gp/wJpskRGewxOrLI0liCjeMrB92+d0SgtCAxzK
Vc24uW9xDRzGX3icQ+7RDEKIZyIhFuid42dHgYQF++NTwVvG+2qmhZgHjnT5nqgx
+AECjU7YVeEzsscjnN9rJmXaDASg8Qr+bKM1AbGhWP7259tUTLtruOuOExBl4Heu
XEblh35ksD7svb/vNt8JNq7RCOLDNY99Rh8VWwJIsLJ7ilz83/QyM42PG7KJz4YF
Vr9yQDZgC0sA0caDeFLBlx9RSbB1t8o18P8eG7ujvObYsmcuK73Mjim14Y6MmD7Q
PssQlc73MkmK0S0mQyegJ8NU9PMiqg6TlxpJP8DSQ2kLuQ4KRW98bPdn9orPlh8v
LSp73Jsl8yre3vslmzjJAshE3LwMqfxc4pV2tcTnrVKkXeLRe3cJuqkPmGaCyUKe
wiNifvfu/HBiRxY2nDthguUublIguD7H6zyAjVJlVjfH4xWs48536xM7eQZhhQTH
i39Un1cZzPrNgGFMmA03sTdNfURXnkG+HnfnmBPFEbG73aQIqegX5F9KA+e8v6O9
JqtUGsvdkPfqq1o8NGl/dbD8SCU8Gt3RWoWjYCfObvIYd/F4/CRPs+mmsWDsBr2M
rFkyT+eGCPNFouo2pgGPtbByQc2xGQk9TQMfKMmucAgRonZIlYYMjpHekcea6I9+
uNoeI0D/xo41HbfQIafq6R0H83gAr/rX4u+rJK7cgu/+GgmtIlNzXsN21kcE4ZVU
NEs8+I/7kuMXfOeRpvbXMNi/3Tv4Cq7/4Qod4ZIDGJTi54YrIk5b6ghrIKGGNXw0
8LM+MouSSIzdEH3J/jd9gjRqVxI/NjXoudlAL4XPmFjtst314cjkNbkfeHHtoQM0
47QWycHX2Xi/xiJlfCLuRV3/cmLl7MDzc41hk0iuP/HHaNPEOxc/QgyUiaVYjSMQ
ag1BvHzzj2+idiCQhWGpzBIUVQi3/aTqp0ml0ic6ujyBtLhzYD4T7cQW/R6bYFDp
jUUMDBoz34jaI/zh1Ad9gjPdJMXEqC7fEtSkKooFFqKYa00WdLXZnfSfOCV/jL6X
X8DXRZKPUHceRn6E9kbvQi1K1OWHnb5ErE0KCU/qTEwZpNv7BuBR9WeppUO0jgwJ
lo2+Ys8gLs2Syq/PA1mRfFCEDsOvml/swjBrR3Y4FgBeV+nhmlp74HEAsY01WF8D
LLC8sQen/OlC60ZRvI5dnEoVrijFSSY25R9cYqrgCrq1dSxxMaGg/8ojVNl471xP
c371IPOPN2BUu7Q8oYyG4NgHC1TrHDdGIj6BOIGtvRZbrHEvnqN2Sr5LAGWfFjev
YwILwmkD5GlViA+OW5owcE03IWATiGYtznFCxEFLeqUnQpkNZvksGIuxCP0zXnsS
WE5vGA/VH4JQr9NcN1O4Yk7oY/y2Ekt/+ex0rHj9YVMaMY/i2UlK45zwc+Q+pWNd
PcJMKVfH6GOdjysdJSGg2/eK9rRiswQFdOSfWfrSatpCv+jroziDAbAdL4IHlOyf
tmn1TJs1l51X4EEsT/vg2RU62CK/QDkfMwGkdXDEc14L2XemMED0UvexChK44HiH
kV9Wy901y5V1RDDhMyk5BbLTs2xyIBQQEMS0Z2swyHkMMKShjFZKdEk5PsWREl/d
kv5ok08nhoHDUNx/6iRn1JDqKhm39SsAgSN/5PY5cHBBKpBEz+rxJh52KoO3faZg
7giIN+VBeODf+LN+IjAibsw4pLKHo9GKerkb0pUUEpd9Kjf86YrHIwLYWK8on01N
o+DFcUtpkr7Ypx9pPpkgRuZuaGm1e5kt+JO443ZPdMqtLyw6F3FiPRfy5jaEcBQ+
s2fDWEcbpPThKQikOtJhwrODubRt5Pnmom5FiUqOKNkIXtOvZfw3HJlQ44d8V5v2
usb6UzFYWgSXBQBnxIexZLFFhrSXqMc+Q8biaKfeTrQE2JNchO3LNy7n5syUDXgr
nIvplcA4bUM7NmKDniyMqVzb5pos/gUP8YgglfHB53a9rPhTeFt72vA2+ZbiCbLi
CdC6HPtPXuhLKWc01g0QaVEuGfGcl+moxIdjcrc52s3MuQj9rYFZfNfqgI2fsZ49
0SWO+mh2iXMZl2wc/PTZXPsCyHataTD6Dun1gQtdhVqfxuhMSU2CLxPY3D/RtFFI
mCPF7wt8s9pNhiNod5pByHMtQMPdnWFjyCNp5I6yeW8YABc5e+WEzTPFB9K3Johk
zrU5yKvKOBnGuS9wWshTVBQzZIUDzeF++cwqGQhXJ1Qb5ramsql6kf1HpbmKGzhj
IDZVIiDGaxQXld6Rlo5fE6tCf2/WcbxhCMKJBNm5kYwWv7aYMBE7DILQLSIWNReE
zRvREGPE7jcr3jCZvXQSq/AljnK5Jh5eNV8xzJt0og7SUUwTJNyUSz3ur/Qg6Rvw
zzruPCSqjaSRaNduGUslVyxmybdojrgnQZ8XRu0gJCJEhonqkmxobq6eloQly94O
fkHo2EzTam/yhLt+3SDkimB8USC4NorFWGMdlSOezArrZWyj54Xd/exMdgyKcvtc
ratWWB6lYotjlPbLgynG4bIhVAV7WJJPn2w79mMs7vuDTyuZ4I3geZOGncpgfIHH
FZj94JIYEntSNNO9Mpts/5gP6WB+6XKvnG3KGePYAuZ8LBPeQk1gHRUnxL128yG9
caJ947yyoVuG9XQUqlilvVigLLhwBB9Fktca19rpJl+NMbmym9QIHQTtVuPYgJor
vVEkGUbWIsFylHJuvyRnsTIr7PrC8mmhcA/FfB1Qmjg+Jw8NSfeGMUfK3k2IDjbQ
fmFdW/anOYXR89Id+sUwxZXlOffscWk7r6Bv3Lvp3+DdfR5TQgWeE7dSmYtHVup7
BCeWs8iSWuWfQY1MFq9QXbRYYymjLp/66Hmc5JE2vXcw5pKOWiGujdBbsk7ZH2or
ji4c4pGldOs0aTp+bN9S3DkG77jEs9fRkQeUCxK1nVqage8pVu7k1FnAZoRgkVgO
8Bez9IkRY6g6P/KNvtII8Db0bB+rqZ2jPNQVhaKHZRuKD7h4Wgqd68oyeCE7j+mA
MIeiXJ9AsKAm9aAhwZm+LNKFmvQ+zuxNAD95wETy8fuvGiDw/Nz0x5GCrUOY83FB
L07DKKhHqxy4L9kIkzMi4rcyFCIBjdK8ZkaUf7z+os8oI2orIr2B9qmBp/9YsMvK
mf4mA6gsBK/BPXhRcemE7ym0uM/AKmetPI+a2Jmb+Z6h8BV6V/bLFt9+4Ar4ygg9
24bo6Xo1P+5m3LG5RkwpE9btA81q9p5Ldxn4cEZ49An4I5AooomkRjySm0j4tH6Q
3NP9cpFetNSW/qVI8I5k1W+oPCx7hf1PF13j14UGWcVWksCBg3hUvfvhYXiwTbMg
BHzyhM8Jd8Shh9wCl4MkpMDgTprd3/CP2HMzsc8owXVIPGPTpyVjrUhTYjZix2nb
PNar69C6dAzGXoF35ks0rfw8rQA1n4f7846hA32OP1GLopku2LFniQ7n5dmmydHa
rnepOvhLzLSsSfLaRSp2Kj4JOf29678d6vIW8r5juRBLyBbXnn76MzBKWP5zuQ3I
ULmK1ZWeY0c9y3byUx5Q1NkIk3VA5c72rrtPOmZdkdMrlW8wgOfPOEUitKO8UMic
/ol3Kx4E567rdsC64zIMyC5X/e+J8TdQQwCo60aRRq07tj35KI51nIenTBrN/fqY
te4mQwv85/XqcXIgRsl4LjqpRGz5umeGke3KBCpUXJ+5q3HMDzaHKZ/QdUcpIG0E
XPcsaUBL/R5jF7Jd4gwkWYjrXgFdtGAxiCk5yylkyyKBTR34YGs10tfx7Q+5Yqei
rELK9smJXhs7YNW3aGqcalg7Lgb6TZljgihZrExhl+/sn0QlsRF8WsQvCNUd+sd0
GevFuRzKUJzxwCmPEw2wou8Ru52h4R2gwvlp5rf1mAsTdcLrye+ZfmZZX9O9NcTz
vpCJ/hk7OUX/u5QkzEMjcdNgI+9NuToGgrnuHyEUl715aYZu7Osxw5rwIbw3ByNX
EA5cLqBW75XBV/H6+izuirS484lnSBDpZdJhb7fdc8kArSKyNL/Q72SvtyiMiwgb
BdOFfOBqbbBhMskw3pK2BCob7Dr3ZRjsbc8N/ctkjYMLgbOxJddEOnt1IO/UmSaL
sgPJDCucgNU8d6ly85sm50nf56ePeNR89Hj+3O4J69mwh0SYUPpNCuTxSHYxszaq
dfGVNN0lOSHr8pmNEavcloNAXtMqVySuB2OOv449cTwHCheYz3V0b33wlZyKJR9j
dWfHefft+C+tNNpEiOGdVK/RZd1qtJoE8v6Bjt0G+se9bYjPjMvaSxOtCbndYCn2
yP5o15AW3fVi6G4lsAoe4EpJSrnDqUR0cQY8ySq1luYsC/O2RGlbXzmr1MdvvE1X
pKeoG8zBBj+zTQRJ8MifEqaMn+MMMAyThTV1kd1P9apfcJP7VxXG38SXlmB1E18M
ODteaqLHeC5oOEI4qlg8I43gQkfQq44/AgHaJQfNnsZYEx83RHfTF5twWfqvxQH8
O5dLIF1rA7EB6kdPg3n0BoEcJO1Y/WvgnsEUsQEJ8NrybCcUbgbsQeYjeYrzhKbf
U+0Mk5J1Sjk7PQ8zuP9PG5lgoQVNjIyPtUmxzUTGPBFN55LOM0wraqcXr6DAB/7H
rOnQftnSzfTC2wyydI9li/sBhSRsnGmB5lP7GXIZU4QRkUcqkZ8zQESEfuB0YNH7
rdyCdl3094Q1pYVli+6APhbv7A0AFrWvHNOwl9NZDwhgVniHXZkjtWZg6nfNa9ZT
oQR+a892aKYakBPPMkVIt3eo2oDiRXjBZPFUW9zEdgJ7XUSjPOqm06XEa7m2ty5Y
Ednw+jSoATYAZKLNsJkmo1j8b3OCcgQY43sc9GXs7tSe7LP3T/kb0arPQa1Vuet0
+z6GtXuwnkpaSMwzYnYfu+p9L5Z6BqoQxJcl128KWESOJ05n1wFK6MrWV9hS77Ag
+VhJm2sEtgqmtdETwQQXpXU59PUq4sb/iGrEjoe9SVqu0zyGSFJCOXWgF5aB+JDa
ebvCdtarRlgcpZuzpYh+oSzoaZqZp3P/zBDVUMLt2r74IwhNDuS56FdSNgwEfFVK
AN2rJ9lqh/fDLYTiI4LevoBX1bgYqQQ+mggwkvjOYWrdLTScjxnk9XwXjfMEcFIG
ySOWL3NzsuH23Z3BYAKPUueNLKfgUjqOKE2qCo7D4gaiMPxT65E78mmZQBRXx1h6
/AaFD7tUjK96kEa2JNEdGFTh9vSenrm5Dmdv4Y87u5vBTCAtUyywKiyYaNH3YRwU
wSKX3Tc9Uh68c3yo8qf9QO2QlZH/3qaiYHwfaD20e9MXD2WwkW3RCOMPMu1sZ8DD
NMYYyKHKh1VHRyxNF/kTzo/uMHPhovE9QxO9vaUfshOLAJEHB4tJzgqDDw9c8m3/
Sj24CsilG2a8mctkP7De3vGAy26TGZeUd0BU0ItXF12hqGTxG90zEoqxLZOTADVI
BrCgDPm+Omlk+HqzMhlg6uUOrynG6FgO0yV/HZNk2BrRgTXqZfjdWv3HmPftcO57
7LWTbFk1uI28se3PFG7LeDRqAVvpUm5691UYgYMhyMeFWmnD2ZWn5comvmIUmjSX
vcDbVbh+ccUJ7Wyqxh1vo0hmHIaVXaUDdVN4KPZ9ol4FCY/8TwcKFO/9feWETvcW
oZF/joJnqODX7y2eLG/P9ksIVs0ZZwvGfBeElPewRlb1OGQ3TRgdzUGvKuczfQlQ
R0TMDjxOYXqw4YQNS3lV5LGZKfIUQwt6OyQCrvhwaCsr7FdTF70cshcPE64/LUfX
QqreyEY4dUfHsN1+z3vPQ9mHItyGu+JMCEk1OVQ60+wNiRkbmFXd152nxYzl84bq
VYhNoAsD2xx0G9n9iazbf5yIfQ/axkEKhx5tnDBX29y5FDFtnADb3ztgJrCDAOnw
/z0p9Kh8jFjHU9eAQSSEHZqYf4SljSJe462bqSv7q8E3c8t4e8/GpViIRk/nmbIy
jv+MrwvaSR7HrQemCExLHeOSbOLHVoDhlANUqSNvt//XpdtETj0trWLfBeZHSffh
VvNZ1tKraeZLi3pXBbMHF7q7NCdQr9fmeri5+bsSkr02iZ9Mxv1fpt+YZjfrKLv5
oQa2Q+2FVCepSkMmIug1C2Qgjbe1dSDCBeMdp2WtZgeWk4BLm2kCzHQFc/quJal9
8UIEwDazlbWPVZDb8gNbovYCVPJ6kMtURK5ViuOUopPe5sRoGqXhwcPp08meo46K
DOmOE//1g8/jC/86NZzrY7SDTPt2kYizknU4XMXJ2VfcHewPUFXAtaurpC0Bl+5I
ud9giqajNs+si9ugYlGlHkGK9Spbmpdzg0J3X4YqQVQZVAbey71TlKSEnUqY30PE
/BymwTfk6veUjL2x3pXNYN8+H75TRQp/G/ML02tNqH3k+6h5FNltuAVmnQ/BHgYr
0ISPLHSgyUrPLoE2dRzRWvXB4rV/PuhDO0A8lyiWNidJPZulprAxOAfs50UBX8Jl
8ju0C2QP3HnHgCNnOjIdDHfALWdCmBO67+Mmgo3n+GT4576BGyjFoLsGmeju/ud4
8bgXEz0IHo6EacWZa4nNXTVeEB+zMBboKA071ZgBH+PjYz3iRGMlK6ivDklrieB9
hmTziBsl+YQ6RaK1UkNtiW5ugCZHtlFHo+fOv+sqGDMG9DcPanBPXG7ARxkdeb5H
ahHaTaFSgBuYpCKkBtaeGcfG74h5kJgDBq/AliVC/sohtr+TTW79V2qLEF5iJv8P
MrX3Hh9WaesYEz7iQgVukSIxEtpXYky+QbeI3xmQemqXBad2daJlAuaukhKIb4p5
0SfSS3xS9f/q8Rg7Fp6U3xlxj3RKPs9nirmt3VpCF0HHVqE55yWHX30X/UodGOzT
OFmFXiwDw3KUojqXck0dHZRiRSgipkf1un+dleBNcStiwjoc6uQlkjp6IstJ3Qxu
ceoYUst7iAOUM833bGzKJqJ33euFakSRBddLuCW4gswwsHn3ZVCTrC4q6Mvqwbav
VwzoA9oilllWeNojvFpb5H4oAJgO6OVuaze8yuabDEVZBXI3kleDn7BXrGZCusw7
Xgiod28MqWVxPGoQBuhdVu1JLaC5VkLi6jFYfilii+tLCfWeouYpssJfGJh4Vw8X
E5W0IR8VDl0qRVy3ZMsV2m8yQfilSnxnjVsrHKgugWF6HbvJr1RZb5DerwsTfg/x
vu7xhOWhfBVHbS1YWF0IgPircgjS5XY5/GrCswIg7xcEAq6m4/UiPD+ghcSl41u4
+c/GU+IpbMoTl4SujTadXkAy2mzAD9CBMCv5+TWcWv9SvSnZUmwxLqO216zsyyrQ
tIzUvYHbgRvaiUGuxuenw56qcv0x3LQ4Y31+CbXTl6oMnPbiBv3q/+b8gDuKRfT/
W+KfOL4GpoWpoSYwPDWStP/6GMrkrSCXDI4OJTyxs0zboogMVgM++ZYNkiU8wKJ0
ZwszDILzyZldd2WtOIDdLnk2sTIh/0LGuh8Z/CevYojcuJHibQk8AHgkIRmsQ0xf
reHLJ1c4piVUfkFWhTBuJLuPe0TCLBDm75TVBg1KklIr0BUItYQnffonGyYBuoqF
Qb6joUU8c5qH+2bQPqcXFyTh2uz6qJwfw5BQSsGh822azZvfA1wgTJk0HPgX93Cy
5bxhWHMOEALQq/Cx3N4/ktza1mlvzUbAkQXfd0i48x2q0WvwbgIwJpOj2aafDWtA
p9XZvNAFaiLq2n05HHu4kTv2feYXacImSB3+Itj+GsQtE9QRaYXbwtEy3J4ObP2A
nvPhkoz4EqXSujfjfiOgJFfjSL61JgjzebinaxYjP27g4CnIrkYgnx+qWPGcz5qh
IGcNsI8gPABI+yrlRygEM1UB8i1GRMWYmjIaXiWrVXd0YlCJxtOOZO8w6hytm7om
RTPj98ThtlGlu5NjpxV5C4ejrNDEoH1xg3oiAmCoME89jpIYhmP6SnfrT+7vlY2h
wc+RGeWuzFC0Yu78xwbAB7ziMfxofYDFmCPfg6JrdTZaz527RTm/ckanvRE9Tt0K
UBXhXveZPz0HF3haSd6jDMtaXiZ0Rn/u0UKeYb3Gu9MrHj+nVynHRt5noB4eAEOJ
2FsSui3gQcJ/e1tIh3czCotAJUFpH8Mzn5m/tK0fJ0AakeZGXaE0WJy4yagKPK4a
tWriLf6Iy8r/l9jW8eA2HDuwWdHiBX+R9A3nceNlZ0lrNbTSTMv9FH/EYB//YVqy
IvgMEzqkSYVkkuyT0ImKGRfbfHS5oRGdO8XdXHzRMIMyDGPxgXmYbvfWUpi0h4+C
zx4M1I0YCf+1p3tVUM6z854a0TmxZI6sR4mfqE6rnXQRnAgK5fcyQuMqBE3VQBhH
Qdy3JJrwit1e3+wbR2CccYWC6cg/CZ/LVmlEAIwjfzs/6lS3mOhessAK6wKAmaaf
+vPJWRJXNjGgLGMTBUmmHa2wFeASlALQKoAmGNC2abcWcSIOr5FWFs8ny1nkFzuA
QEWx6zrx3GhLclfPQx9zsxnMTYHdVJuLS3mxCBMUgHDUw4mt/U0G67TgcNs80GTp
C9UiRK06/awQkvRY2xNPYccy8izfVQzMC2ZWl6vCSYIFYJR412zU1d3hgkGR4Y9j
So3/DPdlSrbwmrdlhm72KfLLLlbFj1cvwmgNEPklz7Wz6mfwl2936ddMN2XEHm4w
hRwlbMXitW5X7jF4gtLnlPMVJiSNmuwCvlxthag0Rj5DuzvPZT1bmX2U5XT7Bty4
QJ6dFM2RAuq3sgoeiWKAA2pQ23vEJMy1QFrecO5E/oXaWIa5Y6qhu4G7UeNhbLlt
P4uvpW+/eqqm1nxeldZJcAwuTyiM9nxIsHVimT7NBg2hUOEuvJgNEXL9qNKKTWie
Wcix5HawjX3kzN51ABVWExTSj6+cE71j9RfgJiLi1kuMpHPZSTdtC4NomfzTtcXr
Xkjp2jAtYKvSmSiM8EnB4PC5wtk6lAYMbCI415uGxG979bmpTqf1qoYestb+/J5A
bv6RClH1j7RMBBm5cuJ+OuBiovRIfoLbehH8ru38IUsCC9DSgkfPmvCjdadRERLu
7qtjsNa6j+HjmzNczIGjDVotnT33VUJS7JRff4s2WbdSpkhuawky6tdMQAT3jXth
R8OuXkqLqgACqOf12gpW+1a42gcFRs2CwY4q5K3pWJdUvsNAPZI6zQAFTbrq1z+r
+eozqcfbuxnUYLEeLiTeF9kFvuIRuwGNt+SsYztQg0I5OXkitjK//lKSiELTbAxT
4JirCKvG7SC8OXuvf44AnngmoKOLcxtb6FO6viF7rtTnSTmwC7mW3p5PiVW5lxef
tLtJn/EkgPUlCIbC5rP35SKRKQ9xCM9nnYUxEgodbBcxIT9O89JW1ypJ5m1cihnP
ghFMagksThxDC5D21k2lgLbEPJ6DUxnMsNQWf5/urP8FS657xdjR9pDGvAYAQTF0
tpXIYdn8z2btN3ERY4dEqxsH7WybhfMAYSvUrUiHJ8kIiiFfyyyQTdSwfXSIURKG
vkq/Vr8xUnMT2HRNZP52xzhZScfmDR3qhVRs6fLHQoMmQ1XtRo9a5FsXAVgUY/kF
GecHbPZLadXHBeZ9kNrML0yUrxagnAIEJbPexN6MrCJCOq/UnSBWyuyPB2UofqX/
YqUH6TKmiWKFMv3c83xbAUDni1USBy5cUk/reUIkuFeFaxM6BRuVL01+27MModlI
+OCehTrzqDO8x1anyqkUJEUulgTS5gFmQqivPea7oONjtShgYI1lS0NBbTjDXAst
x9FTRAfXqOVsIdnacuD3ehAOVcJq2i5NRpzvfQqhDMW+m/HUvH3ah+xyitWF5Cgt
PXHlt9fCBy0669tEANG2FukAmsDOd//fm06vLaVpZQCueey6cd3cBakNoN83FAZp
BrpC1RRX5B6qU+5quBajsks1SMxwU9Z+ZhfBnd46DchwBZ35XYfTUXJLly/71GwX
PO531ItU6ClQuFhhRQ3SS+42gxjdI/4CHCVPcv3aPj+RS73qwowjzUaFMV3j2h/O
6vvuAzTAUOIYuxrq6bFtnwIUGfhcfmGEeCdYfmJNmMbEmwdbol9mArzg04+8CESx
07ZTYhRD8KFIrKMkNhUe+rfGMwKCmfLYExdfSXWcOk4+DzGB2VmwqiNG/F3V1xOj
jdC7jXeuCnAm0qjQqeDDxHB66sSWoJaXl/yMmJqPEcUr99RnRpKH8c8OhsPmxf7n
ZafxpjAGs1M/PioXkf9kPGRwmMp/XotbdN1vX5Q0pKgVPIPBe6Qc5FOSvNLIE8U6
4uGd/0k1sQlt+Y5suy23uVHPUoLxcxBRnSKwaKOwoEC4REjZYXDLIq3iTHttQMYC
w0z8/DWz2Trb1r0ixSbAHZSPa88xxFtx+btmrhdNzdYOOw0hItSrTkhhfUhfyk96
n/vmR6ouuebtYO5Iln1h7QKam0z0bccPKtBw+znQdzXLRVHQB8P4q81jIYeHAYwz
/yv6J7NkDu37+MWj4qNdImp2m0iOWUX+WDXxU4AYCtJUHAyPfSq5hTg0r0nGBi+4
dzTExpEZclQErltsTYcwQmbFaDdU0fPkdynFNOSA7kxmmEN5Z+O6MPTZE4uPIk5F
j/JzuRnRiN6u+7cnsZt7MPQrwVjl4/IPJpDUmIHZNcBZnwEYlSICyMPcBVCEiFCO
6wNpUcr0CpgcuXfn77CTasB64rZcDvDW69qWOGr6Aibgs3x721sAttNtzlxYAyok
NHcACuiB0IMvpRdXZidU7hoHj6jEtRS2xEJQ8I3ui1lmcBCxchqcxVIsv5h+NV8u
/6G2HthGt4W1F/KCX5lYPHQAfgWAH1GjPihXx+jgt6xCduVVucgeitpV3aorKwpb
rd6yf+vYkL5UGhg/Yqhj6ReIJaF2XLkVrNjBVm4bnrD+DGY8UydVIwI/C/DzcRqn
cSTKVA06Y6WNqctpg1gxpeHeOw3KzByQBLgemWdKP8eqc7k8V+XipC5X6koI8HQu
3rh6nR3c5CaTlwQrfY5AQnDMuML7b+v4eRrCMZWkRztL+jNUgUqd6kR7xdDM3ch2
gCuhQwumTm+gQj2cGH//bLUpGl/M42uHLObHFu3L+TYs0t2dyE7nYUnZuQ1M1XsJ
qTyS29SKZsl2sWc+Mm3+ze5vRGs8KUw4nr19o9qfsvnOAvZR4FhuC2+23JUED6q7
nZig7sxKJmN6QVCKRxi+D7l+G9NRWXOkTac675lUxm3d+k0c0zPb9epZP9v6Yv2x
riLGEl7RzRxjRP9svcYl6fOmPK9YgA5LBaCb9prANnJDjwwcr/sXoEuxXJ7RLHK7
mkLEtPmqUjc0HZt+3Xw+Db1cyfbPSWi2Eh7ql5LM8KwZ0wbWLS62TnUfaFBBSLfr
iU8b4PXVmVqRLW8pcqYYOn2/nIpghLB0NLzcJlp+P0y2wfEkO8M+m5o8m9psWWP6
74XwJByp2/Irr731VT+SPN2a1gu/DTOFFDsXpLZGLo27QiNUUvY2bluSF2Tz/NoC
gjbLMvwanEC6xoUptz8f7pRJRrUEf4JoYuro+aJgTjHRnqyNb/8yxyONbfGx44tA
/7qoXJE9+hP8Ix1y8hqhQu4EikSvB/gJpigzlTMIbl9zu+xbEYw00DQ5tZtkO6Ua
4tP8+kk9vMPg/nzaOH7wQzpAeTOYUIN83CfzbQY9ZdPeaJb87uVfTmljvKqP8m3U
4/4KuPg4Kjp3bIbn3DRAXP4lcHkWVM3H3sL9YSfiQOH9IcoYSDs+q7P+X8sTzDBP
w7jbyWTAZUMLjm0GxZ37UKADfbrBaJypqzbikKSsna9wh9HVZ0pJS8u9QLiT/Usy
9m6kMyUgZ7Q95K9T0wvHWEosX1gMy1FBA78S38HQR/w/DGk+W0EaKOUPrXtpCdbs
f06Y642Omf3QWhtV1wPuMguJVoTK5rMxVj+dGTX4J/pRwLIXHvCoW061wmCphKPV
L/mqnsxhPfMfrSIcUTTVVCZGFtLlVGn6H8ceQAtNkrtQJLfp630G0vZuTO4ehFGV
qwIDs5vWqideFivMThL2GTKAvZ/iPvH57J5JdNzDg46qhPm0pJDKyovSW2cjnLNY
3WQj5IygB1ImV0VqJYYSHLwFKh9bmiQF9nf14JEzkBXkcRj9IrfcPl5vMGVkDp8L
//EiCvjJxM4zS5y/MFdgNrwwEr03F0C77uy04M5wy00Nki7t3oWuybebD2i/Hunk
/Qjc8RyAuhIqXljWyOh7m0EBhLbWEwZapegLGTZSgJaWLW7GkOc5a6xYzWXatQkR
7rmMusnqgiPVrSQF4CJFlmRnFIaFeV3ma8wr5zpjUxZYlxczwASKCEW33l/wGxmD
o0a4uKxRjn6YpLDCnwSexOF5qJAq8NyMf/w31mcQxT34PTOsIJe5ejIv/Cl+L0hT
BC62aXeegPNl6l+MfFuThlMIhRnMxkg+nG8ptlApT6sTpoR8LwZ3YlqidtrRx917
GZz+4vdQtB6bZTX2KjuqepfwWIR1covMQf0p5Ln9vI6pn8yMjjuHM3//oOmrrGyV
IRrHTMxcDwbXIHFFSrpAQbJspJ+K8R1WlfNJSO7IPJ55JohoPxUtAg9cTE2P67Wi
OsW0l2GFjP7i2+xAqADIbXHCW/lj0jtwczHvJOmfCFxXesAh6c0HZbM3uWH3O2JF
baq55cCsld3neXjvvWVe+MXQj0SU/vhPHhQkeQ30jsoC6rXKnftdwssemuPGcgXh
LfVUUjUpXewK4fzsvEWGglf4XbEYuAwSiNq85Ybw5q8W3xkRywLFUZBzqjdaWfXl
Weofd6UEhJsSR+bRoIfe/+sBoQkwVyvc86g9XSdnLNxwcahGPbixgqb/qMNld4/+
lHNTy9ELGOossUPZRpV/g/1NNM+WRR6RwMJJuCscGmGHmRfuyGgJ0jyX3SL6Gf2M
gSV2S5BtDX7JibD0dF2nw1a/1ruXKLMFkPNC8pYZPkk0d6sdbEqpId8/vDkOvFiU
CQ8JWEd1A4MpZV0YD4V8cblOCqAF1zSdE5JpLagdoG1fOfa9WvZ9cH1/m+dLy57S
LdqFAtUHEWpqUKKZbJJhGKzpMvHQX77IKKM1I6Jq9iGTVqbBfNc8+I9qZ7d0KTYC
xxRaRjGx4Bu/y19lMdFrNiqMchgOnCDom7lnZGEORw/DiV71GXGcSPfXNt63xDlW
I6idum8k8+1b737qJMp6Q9PFj57WrKIjmBEW3XS37XWFm7PKkRiJzNifZkueYY34
xcIj8j7gfLr/VocXugclRWTWo5/+LiiqBtUBFEDFRGDW6TwxVfYSo3Fp7sCmGmpT
KMcXu1RdUcJ4yHzO2vbjDmyp+fIlI1EgBuIQAsicCkz83SwPcADin6ByxwyzW6+D
JTHwGB1ElQsKJ7GQGu6llVYUvGHh+6fQsRxx1nVDhWRGJ+AkpReSQy0NUKlSXDGi
m17jx8cAJAdpkmEWUPmeXU3Fq2X6NHch2TQmib7zXCx4rb4kgD89/g0f7BAUIjGr
2dEEx+nsu2+tAbTUV0PLNQ1lZoi0E1xqFvpNERujbpXaX6NoNPv8J0Bc9ao6iQf3
P9zYoxXJRT6aFc+RdZtdR42Gp/8ka2K9OBofKJmN89vjEyRIPx4pUZ5/5jplKEv/
jM/2TBS7PUrMAR+K66W64Fs50nCrXN6QNp0prYpRF8m85P9yqcRXl2firvonACTP
WrQ9ZnvoD9qVW8JtqEzrY0kWyiHhFBGacD14qU1Cm4KsliQxPw4TIa0pCF1rgNas
ZrnzCnin7ldqaLP111htlTxoaVrqI/o04zezPn5QFUM5hRaEEEYZMXHc+tNhsTli
Drz4en928EVwD+blZZLz/ZDZY7pj48p8FIsOuOpQY/FjhRkUTLb8BdKrxLQx9NY+
ejrWfnEMArDtDTNgfeCb2IT47dGiib6fvSWlZwfHvN+Y114d+IQF/qbsAyLx7d3b
7RfUgd7SKA+kF7ifSbbOd1pUfpfjzgZGMRfSdzzJBCPlVArVMiOJOTAfuq7l9r1F
EDr7PXjpo/zAbbZqntJYi8u7f3tHf0vP6ghD+xYPUJGIsObHnO0nfAZc1ROhJ3A6
eGSvMmBlSj0jtHfnRsNtZt9rJ3vrvaDsBfFD1otoWcKfBxHiJO56JO6+da2F0ECv
0dCsdxBwo905Pnb5jG+VHlq6hEQiknLwXL6mOLA4sJU9z/7NpMBdUYrKROBdm466
UyLx850FdzM0mqsnCS4Ulq7AR5T0ulL0mEzRQr1qD3cq6/rhwwLrOYrAZ4iHdLl/
y+PmB52kb2pKH6HeRSBr/zHMq4ROePM40ZAVFFtl60lIiT2T+utehPrtVL09i9MR
uEGSlEnrjyBjPt8PyStLYTtnAm2qqkcAC9O5b3IfKUOsKEUYlQYsxI6lZ/5mCMhj
rQIFCFrwSI/oY3qFOSr9/IYW5TsxZhPZwAwG85ut5WR5uvYHh2o35L3z0jXzeTM1
v3EHijRjNwPUS9ghJexHJzdVuaorwDVmv4QhIYZFLpi08V6zR6F87rM7Y9IN5tUv
/fyqR0pkHt5AGvpFtg1zwT3OPYyQ92DYAHBMVdjiuk7bMsKq6wi7QNtJ/WoNq9B8
W1wYaPm9TiG8pNkNvm1Yza1pqPOpPmZb6nNPTpke1eL4nRW6QuZ9nf4N9LUMuupJ
Z/6VEUPFmVNWgA6u15XWhdib9Tf+/sVH1N1TYooLeWfmLrAreMQetAlJZxTSy4Xy
D/05MV0jakcG3AqtEGaYOgQUK2BafPH70eDnnuG0z7DmTtjudsmIsclZmoAV2BtG
42qEmkuW4idEA3SCqebOkB7N64nggI/gx8LOUM2rSEyJXlA+uD/qsi0rYyyVPsUg
m2HXdPO3ND71DYs1oVYKv/wSGGxdAWqE2Rd6BfY2QLj+spFlGA+GIVeHlRZ8te90
BGs8SIM1E+TaJVUyI5gCqcHqv67017yRodvX4rB/r77Sx1hoidUn2D0jZJShU6Sx
J+xYEM7lNVR1S+Brrq4FnbMlN+6MD2dzawlASLISKL4vn4R+AAJat6abZJ9Ta5FB
zxNNgQ8eRu0lal8LyGcI2HvYalx7kXDwwza9jGT5bX/Pf3N3dixHEH8GOF1cCFB7
KW2HQX19wPJH0XGY1OfLeh0Z3As4g1k/0NfBlzywPP8DZ0Ho49lXg3hi57vbxIXA
7Gi6LTNGAGgI5ojZP61prCgITAuB7TdhPu0rAlQoenMKwEUf/LaIGA9Y6j7jUgRA
iNO/aRQQXiZIlBH+8oeLmWLSN6ds93rvQ7lcN/+lCQXd7JZ4K+6zJ7UhyzOdvR7n
mDAUUh52Ti6+PWaurh2PC5H0adPdOkXM4gKXBnVybHtcFBB93+zO0O3pc67Loy1h
k1MkoNgs6HNz5Ed1S8TZ0h8A+dpDlkO2hOa1DC2bG3PQPCCOci+WB8DEcQ9Ixq8e
/vFO92NDz1x++e4cFOHwu73OapSfuhJXeaAQO7E3kxsN4ZJv1oK/YC++BZyRn45P
9pDjcCbtVaGcjUZRn40mqors+YjpVfUGWxWqUNn7M0g+ceTHnxNEnNozY5jdplMX
kTnvCYceyLPCo5HXG5HvWmMsHiFeNpQNaXtluDN+azIvVKYHmtzttLS7V4110p4h
TViu50HAQPfXGpzHMQRUyLNHsnz5w/cksSCrNSrBs7rv1Tjo1haSuZgB2gDbhXCT
G7KgJAVdYf0VjrOd8x1Vi3ll5gxrSMzoDMLFb1JwSc/GsoUPJpdWPjl0sbNVgSPi
0W34601wlO+7gdY9O0qDTOrJuGMBIZBO8F1C7daddl7nzHooPZV/A2WUH+HPMolR
siUievDn2HcA1M/Lkbsx4B7gJx6Zkt1JKl2JQejXNdsAlhw+tK8MyAwwCwA4S6kk
GIHBdITd/kvNqDV7MZ7Ib1vAh8xqaOrDA3fqRT3dYn3ksvRRo2hnaEpnSYczRaCD
pK+NRD/PPtnNH/ZcLEHVZZDd3pylBypiP9Q/dbHpA7ILEiK/7133UXXg58piSZ9t
u6CMgubkwFYMuBO8t8zAhR7fHTcm5sQgqxOaFjgTEC7Ok+w74UVnl/C2r1QPe4/U
IKDolehcnBR4ZrMBDHL8PevK7nMakwCNaMop6wNqdzurep+MDJW5F7T1sj6f99nM
m6Q+ctaJPXhFIoujDrcssDCtuNfQBANCSuahtPrtRgSuBwf2xpxCc5W6qsyqahSj
ElNO4nAz5dBSshTwEe7r03WOTg1xT1g6HuR4VRuUYH0YbNvORRoTbS7KXzaYJ6Aa
6mO3JCfB6uoseI1xQvvgV74RxJwcGHmQQaAHtkk/y2CIBKTTb2PbElp2hZzM7PON
/JlXWwm0rrzdxnK0a2e8KwaHzSc2phevchVfSXtgaQFwpNC2vXdijXgU/n4aMkAc
pdxmRbgErMTGgQFQBJVulSzKVrLHaiXpRNChUaQrahRjnKyH9lE4IXXwAWHAD6n/
DCmLcdHEimY+GSdSY6o2Dp06Q3tw0hqDU8UUscF6O0j8wgUlIeE4BlaUQw4pfPPP
WBoh15nsq+TJ4FmNnPS55gcH7qqzA0kucL4RoxMpmEbstYZjzixf36l2Py9zROFG
7uMm+0+Y0GTq015hV7I+6zIryVsZc28yxUacQyCTBL48dnidRPnu9WRNPQp4JNzc
ejOoPdWv5h38pAX2whoKUW1IDcZvgGTbgBy4kema5nJvWLO8sHhN67kCYbExl6rd
Mi4paw1Kas8l5R/8LXlb7GogwstOwArSA2uomZLoDqpt0biJR8LrC7j5p6VNwuxn
D6ecO9A1m1IngC00idYvsRSkvdKx24dpgFhwxqZjHGgV2zv8+S7cdf4qXV9uNDYT
xHiNu0qR/XbY3+MiPo7PejtAKJvwf57QIKszmz02ZQiWC1IQwRHSqZNrLQwpVrA/
UG8va3KVIysXQL7hji7/VxlTm5RvbLStRCoTTgl5HINLT+bq2dwCcY39ukc/58Fm
FgzYhy62QHS6K/gEZ8hYruBvtQYwPpsm1oYpCFhabdrz7AuRPXS7/l+F9f0h8zlh
1Zz/N6P7N8N1AeLz+0oRvXNpJtY5/WjVp83/GWwGSwXOzvuHAOBQUAhs5c3weBj9
tOAZK6Baa8OhIHN5HIFbDijP1n1yg0SO2qOVuuGFKqirOLt5dVW3+KhS6mImRkNG
2F71okvjvvSGddw4m4WzeAbqy1EH9ZH1ap2FetKxzMd8QHnz8WS4SRTcD3Uryp5+
eQi/abpY2isAqSIaTF2Q8hTFbXgKXkrTHRrJqYltkC9bLp0/isO5PMvFlPhe4Jrp
G6nvqW8Mt6j/RGjodSJ4zcwJwQqG1/6yhGUD5s3IC1Q4diVzwkWBp2yzFM4cS2mr
TDCUlzIWFZMY6SfoTTynxhRJKfGewUE7UDLypQtuv6g0prymW/8VqiHSvibSCTZ9
7RtCRsThwXq6h9c1YlFnU6EJMSAv4lLRAwQNWmldmeQqLCACYYXf5ICD6k1z3nCz
ly29NIBZeUCYLl1zxAHR11jM62feeiADWgsNxArkEGtaeg0pz2ErW8846N3cgMWR
9VIpdDQ7iRlhixF9Q0IrnM9e6YsBQq4A1mwH8/GGGhoiopVMbRdFrAeitzBlokiG
3aAuptF73MPmR/jYLi9NSwiMQWgFJ4MHuT38v4Pf0JbJIS/8ToYOSZsaPyKDFkD9
ZU/p7TgZbyw2uB/QQS9NgQYa+QoGMEqys5gnv9Jd5bZhOhLjqiapIJwQwMv5mOgd
R++Kd3frATVZBm2XCavg1WrCqVncjWLLVqeFnAlR92ZaZPp/OqSrv4BDwlgaa5Yf
eot+Fpy/t6hh2OShcH6TY/LxzCCo8ik8CZpsy0gI3swplpZX/WtnLgFhzTUiNS0Q
oOruS7tOsuu9WK8mR/P/AUVDfh4bx0xASgpZPko/fhIkjOccidKvyfXJkgCNGpSL
aAzdeWj4J7nElKJAq0KmdCqzmc5uYMSglpCVdGDOwgF26Q0Crsn3cCds/T+xN9AR
t3+N45GN0ZKljB/NxtG4h0e1bIitxcCw+g+z5HQ5McF1E9CVstq2x1k3ka8axTac
yBc2mxJ2Q31XDD+J3kMw4TFwlx0gur1US8tX78hNkD0Ylc3V9bhvxjAfSwyObVdD
txNvx52JEsJ87/dUb2GB6/bWy+6J1MMXQXz+p5dJUzOs5KlMk4y17pr9b1Muygxl
Q3XZSknK47RWUXKUhmFD64KqXpGV3mIDUXI85wSHlvJ6HVwfNpvBN9ErwZyvf55c
1QER0dbOkKioMnFovv+dOdnPBiWSVUc3YykvV/WDBUAA0SNx6ixTubWPxF166MJ6
skabLwVToJ70ZzostKbwcdyIXiPN+PgIvQlAZKzK5buw6g10yU04YZapAG8ZhjG/
VSFXitcr+yb/ltbWxcODo5HFgbdXxz7D9H67J0dM77ao528x4RK3eaONM6qT5nMm
cYlI+xyBZJRwxnA7bj8xVYHNPsce3kJACdWyiRkNSMy3uxbpVr4RFvjd7dsZHg0A
Vw9O5WE6xtCBuH0UWYcaI6wP4PvQXMkuBElHdD65CH2U8UlRnAr+kFWdNyFSUAt4
E7tL4OFqrDNu8MYAWo5qjK8HnhcxoeFMxyjEGXfo5+tywXc+DX6dJbKFlINFp2CY
r9FaFfiLD8plzpa4M9zHEVF8bDZTTyTxR5ykUlV9P1AYB7kDliO/d16BcQGoPyGk
fJ19RVDBqoxgpFARcGf0p4eyfEd9PmvZy7d7c7ZW8xoaTmM2Zy/lGHjooYd9mlVV
qfUMdGJUKx9deWIgUR2XnjNLAQ3PuAMcBrCz9+39l11lEo2t1K4ghlQJv1orUUj0
Ea4zgxjzUytzkR15YUasAw72G75FaJLLJrVjYkXz2ee4MzMM5rlBMzImytBMspIr
cJyUOjTdiaxYp5WPtvz57tCVdnNN711y2UV6wB1w8Jk+DWujTpp4l1d3kI7hk1Pi
rJfse3zWeHYLZH1YWXK6PFtN/wkuXVGHZFeMW0QTtiJee5cyR8e5b2BxR6jItHxR
jzN5t4xvOT+DheCcry57HSnHDAD8S0elbZSvBCZAm+/VBmb8Ytv/AgnkSEMPHoyD
RF5uDO2lUj0MHj92DoVYB+cmuVX9fk29Y5wSW61F6x1Qi3IY6WZRdR9e+6IIXxK4
Pd3FcWO6lOV7aOdLx3+YKpWe++hrZ0cv8AATHA7NIz4c+jMiikUKF6o9Lb/539kD
l9ksA9ojKwLbTDlzbRSPFWOGiw5vEUKCHQrXLkYPLXPjM7bhPCtrsgoyxvlI+pk1
yUnXUc5YkH2HXGADMwstB6b50/nxP61wZcBHjq2DGVqfG/AdI073v2yHrFLw71B4
wwJG5zyvuRHZsNG6surkssftJKRJpDOkmch58J5dJFgrm1Sk8i1PNVRnCJr+oGof
947c5oeJ/6+MCnMGiTGdOdzCxtdYULamD90sEJOvtUjHnhtJkVGzSghzVzvyAP+s
S/PwNb+GKF+fthU5daccQ/yDarZ6H3/T1mCcYo9gx2vfJS/k7FbiWcrPvRz/wl5O
bVmZ5cR0art/PpFu4W9UHKwl2s6Oeo2K0IBPP6rjjgLZHacn53c/KtT08JO1xsSj
donKnzCdUdLKPNq+rw9s8DQP8+dYgDJbA2cqnYCsEAPhCqqNQhh3YxAO/b/4os+D
fV3zGArr01ZmA2PWkbaR0Vlv2xeN2BrpdLQPjwVJQgY0SL/fGJHRnlPvloqOFkF4
Iq7MHDdblk/0HqK7wBtOXyj7Ow8J7R91CbES6dfo9FqobMlIbhNvHrLhSSBPoCPf
3EFIxP8rTrPjWODk1r+hHdlZP05ge/pnTeFR8VYHYa+f2rOYX0CYyh3FciK21RiP
ERNm8z9gT/dGjqeV3H5ZeA5qJa0Dx6UF/z/6CjVZqPMR2Nls4c9B5Jrwt1DV6Ngo
KaPbJr3RKuC0Od5F3aqgp+iAyAw65EZerUsHNbpo9rQhIk3rTh2IxNQBSOuxfkUv
0YmTWlF2alHiPD39v5QM3wXQKrFLnoK8F/RQDArzJW4ENLKMjxMXFhoXjzQPJqXk
rnu3kaqPlTPV3ilzv+zfWxGORhgOjs6FlBpWA4edwkgTlJ0ocFy0IQlNrAJV9n+A
5aEBwp5V1QpV9OxpynSiUVOOBMnPTxtBOz9a9NEBAZXlRvSuoXLzRrLprK7iDkDV
eMP7uVC0+qEkitFuA5Mxn/EX7W+4/MpXxOrSZHJRQC+NchMVwF6rmaP8j3NUDlvG
5tuhNKl140rtTZaXHfj3RkR6tTLPncxIdyDETtXPqb3EOJACzwb8Wwi6jLH+65SD
lIPDRa16jBhqLAIFO5TmUocCXXo+hZaQrTSZ6hPPLKyDd/H/DWg9p5tRrBoTBNUR
kQvQ3JYNIT7L1tv8UEQXGyjL2kOQabDt1mfL4YIo5Q/Ze49MjVmhuRknkUGEDXZG
xgXqVFyCivEVv3JVbE/SZBKbQJBv/bgE4JBqtCDVGWN32jGUv1Eiu5kmQG7yDd6o
93loH4+MNXNg1Qxl7UCcTfJeNlTre6MhFFchi4paVqDDI/6thFDb5pgpXM21XFLp
3B5yj4fhmJyJWPxfCflQ+AcEcvhDj9n9tad3hmN4CWffF8z9Pu37jWD6Vum8pMOz
rzNq9MIPvBff01MAchlgJlqZhSeen608pkxuaB2IpX6C5PvAbK+ockrqx5PYHcw9
KZURGoghnx1PkseXsS9P0o2WlCgm7Yko0dU+9iYVzzc5e6XS9FcO20hxWeldUxGh
W4huHUnl6tC+Ozws9FHYHITmN6GAhaRvrq5Na4QBvkwKWYC8HwwBERXWpzqzn8IA
x3d7NLQ1nPdiIKFQmDeFiy1EAMlPUUJWCIbqGZeUnbLlcg5lrO0Wa4JnxfmK/pxS
VEOtfowGj/+R+PFQWf1KmGGWMksGCjouF8X1e+HKZbBnbrNwzx6MgJ6o3y3JLsJL
qKWz4mEEFLzIsbjqjTqTFICNAr8iPMeMGflAh1YodV0ND9JHRjpuAB60lp5y1WY4
JB7I5+G9vy1X6dr9qq/QMIsrQPGtQ+Ywvprj8jtyTxYEeIsTqBRca8gwza0tAM30
6kpMjre8vws+A5/9SXf4Qz0wTHJiTEpoVZOFY5D2c/69XzeskzOh5+qQfAnZqT1v
ihVFbzL0N77w7R0GE9FoBw7e+kZZTmOVAA4FyS58PFxmrTCJZ2OV+sTey4qfC2i5
lbes7477nOnaKtaz2uTv1nR0dYbjciTNf7CCdERqjsO2rHwwcQCRgDiEOn6IBZKi
R0+Pb5FIK2Fo/iC1gnlS0cWNFgktWp4IBOgtmxdRUh6hy3amu6UB1v7GDooSwmm+
hQzBiL5pxINinuj8vpToCq+eYqwEx1yWyUjUbIHCv6k05X4vpwNhMM74SqD+0kho
QW895y5DSDlna08tDAp7z8M9+94MPrGtGz7WU801tOgad2nC1/+4yQ5VASzX3PRr
CU/b7Kie0CospW7n9ZAYnTmdrqumKI5YR+RI3mx/FKUn0ZcNj6EnSOJTz9B0Eglf
DcGGjzR9hYnRU/47F4B+mofSTISmWkDH2FB2B1sVi03A/D2lhjYdDOiLlHMCd2N9
LEgxe3ycp4VNg3zCCpWKeV5GLS62SHH/yHFMoCRBFF8PGV2krwRWNpPe0kFr1KMe
qmqFccRG7NXWBQkeWUBmZdqii5P3cSIAeyzYwxJicTz4KVkjZUTcOiAl4CFEv5K2
8R79cgrYTtsCab1gZ74ltlBdN5+5jH1H7l9EnZfgHL066780Zohf8kaCgfpzcWhw
Fb+wKp0pPmuuri5pIYwb17WMCxbefsLBjC2177vuNG+tc+xV/PDh9t3n3gWG6FjC
ct92fMa1qv0pMFO6doflWAPL2o0LlQDlmfISk4i6VGRpnu8+CKmrcKIm79yInMtz
lQsVEQ0FDCarcfkFEGA6FI1rtJk4zEvPORxrM+jiPX7wNPVaUgTX8jvkN2B5BPAz
suacg7pSfhZk0wYps62B6Yx7SDhW8jyqCV+eOakTcLzfez6II4j4xbks8+TyoEtS
KXsp/zHXAmLsU1bjh2Z/xOlRM60LBS7ko5EFzPwtV01XRzRd6U4VSFoesTTkWBUz
Ttm3oQAzQNsXMb5Iz/PahTSkQXpfFsWRnDr9ghVrby9T6PtH9jSirfbgjeqBC1pM
qpU1Yyqgof8prnrR9fZ1Y7NJSn1uedzUckIFtUUEKQD7xrXQapUPNWZifl6SrzAI
Ey4YHkVST415RJGZl42whoPg1BBHWXqG9nWwFAQN8uHnTrUCrnFd78vC98PDn3+z
tmeWWvbnLI7NLFFNU5BByhLTQHE1lBcFJRIH2suI1AWszYFk/jI8mfktMMnbYe31
qB6L1hIVKqugQvlaxyWwyI3bqBFvPcEN3SlzOGAbIDXU5RofcizM2srzgdF2sXoc
TrMU1i2rJnzbOhboaNNTeissSapNS3705A0xHHzVAfSuPywDS1Sk0GY5MCnvxUH4
IA+6EPPJjwIRlx9V+hAB4w6sMFq3qwRIAmiEx7OqP7XSTah6Q3pqxFUso73tCyTH
LqPvt93bXb0xoZ6hYRcOzovQYzamTP22YSk4ONC1zdHCI12q01+FNH85e1zSqb81
HZ2ByZyEr61KJ4xwR0Hijco2KF+qnc4aoYv/IfYfXKr0A7GOKhb1kjXHQ7UTQR3b
XjoVCDXQ8s3EDNqnDIPJJMzziJ2VEmf+fjBcBNnXQE+OFCjtMePp12D0LviJliL/
bxWDcRHapLMipSLNE7vCsOkZqZheWy+jIT+ux28h4ffmeKladkU2BoT+02eJA1Jq
z/VHr69RgeFPE85UI3fA/pjydXAfatfWEC8fkSKJ31T0d5ktDWKfLWlw5jSUE0ME
GK0DY2YzwoRZAF6cO4p0WgYMzF6l23DXVYEYKB/9I4Rkp8qVhtwOUdZbxVVvmGJB
GzNCq4vZCDTbnLzGVZoD23+g6ttRWYhhntk3Hl9aPxJMLRSKXGlfOJxMfuMbRsEk
7ogKo3MOX2J5UIz7IdtmYIcpR18WzeZn1y1Y4Jwsl6wEQvjOAoEUcY8S2qOhSDDj
BoBWC/XiDwX/FPshtzPnMWk2RzCAQKDL/FQcHg/EEuTpSF0UzpzTOP+QwblEDHb3
no39LsTwxqF/B3LXX4v6Fmn9yLuVdAhebiW4EfQZQyqTNk2a5xblzH9jNWREo7Wx
aWKKf1Ho20NKrOS7dsKOsZ3bzwJLUkrhvODiuKxxQgfyTeYqAbOnmWy3MZemrfHr
QDYGk2oNB8LgQ0jazwHESDwVWbJQmt4k2RlQ/av3tIpKTvExoO272335qW3Hpypi
Ftf8V3Nn21RRg9FXnGMakzmQ9NasioWWdlKTCC+Agv6jtQJaQgUUB8ttPiLzyI/M
3R6RdHTkiI1CTD+7hKq61A9tKQIk/B1Bu4DEHbhfp/14YYuRdxAolb6j2wTOnDiS
66KfYRVyA+B5WdakFgbNiFKhxvAmI5aBclQccThvzmeYztRvyDhzOEywToojobE+
t7LizkAUjS77Aq/8dRH3sWKZlSBgFN2lP4jYVwAmsfj1ZTLU38BUfxcWNHH95UWv
wsKxYCRgTgLm06je4q9YrmXIC9LBbPMipaSJWGbBZHQ321kPMprdFO2Jda5130AJ
GJiL9SISKy5+SubQKeBOMYk8uQF9TI+DPutSpcTnTivUu6+O6VnosR7qLvu0ljYx
DSRN0yCyX4tHZidWJ94Ek9mw9UWgiKjpFVE+N3aLOKwlJuTJLOC6FwE//ktxgXr+
TMs6zmrOY5QIdqIIhlleOOy3LJZFj2gaABPck/tLlNiTKq2UJ9oy5ocCKa2Fvouq
3VNMlfz9ucV3a/TXDXj6zN/gf0lMYuHcnJF4RBzXhn+KTjcf2PHv5wGWGw6SQnNT
6RdYxpJt/vF50zlqk3fAf5GOz8l35LFw74vGl45iQVM/5W9oLv537UxNiSIsPZDB
OH2JKYlYfbZvE4JQh/ExYeltWhR49rPyEU5my+cs2UmGnOw52DfC57MrwU9m3SiG
yDSRZDfKDaC0kVt8ezoL9DpmIiWqmOCMRhQLyttafZxKj50UO6a1Baz73Xx3tF/A
dN85WBn9XxAnV0OdQ48nzvlNCpYXt7QWAo9N1CWoI8w3zr3/UcCqB8xkFD4L27rw
EMFqQutU+KFzCth18z8SVmpFVVeREIYsNFklD/INVNLaB0WdJkYvB1PIrEUE7sC2
ldrZ/I6Si8zkDavNcPrrvBff8KhYONSAahyC5vWn/2Hn97Sz6IqeGpuFC+xbx1Jw
5TGzKgkPGgtYMr8dRs+4OUMKlAs3vKVm8M1JdbRBaL6Qx+5Wch/gfJ3xJbaWPJkh
Op9uqAxwvtBhz2sVyeg9SKEqukCCmTlark2CqX9vkSIhMIWBT2t6HgN0xOHiGzOB
Lyt6AuYrZSLy8asetfE0F8eO3rAphDnVFkNE7aS41iMGpuCMo65uioSuagvG4+fR
CmXdcHclKJRDzFM18zm5p1wpZfSbdjJfOhcHZiRI7pHy2KWoU2sbgaXGHdPfPRYY
vl36uSZR+y5Vu5/ZiHN6sl3WUTd+ptlCYmv/9aeMPGUyx086oHbs5GHR1QK+9bwx
Ie7Tof4AY29T1qmD0RBqcpdJXG5Du5945e3I1bTw8Y8yOF92348fQN69otVzFV0q
kcobDItxyTT7t2XZob+pmL6lMCGlqbyq9t5MB2Ga0btqdLH8NPmBrfYZ27T5Plcw
nDrDABNIMyfoHogNW0eFDc+W/tQM1g5fMwts4Rgb6SFj1NNqWoH5S0kJmPwOebia
MExc+4vWWmfbjd8PuRRRqf1KV7UepD9pKJ/ICVPQLfgNZxWybylwmvkEluVReYCc
eLSqcw+z0fF7h0tOz02v3s56r2XNT2HJsibAYPUQ1sFXQv3QeDcZx0FFX+sVd5sV
qb3WOZWhS2yWPoCxUs26OD0S0UUzGlbO+EAfoF6Nu8Xvw8F1+hZ5u5PRBjDrIOBS
vJdBciU8j4GBFCjf0tA2crqLxBdeCR4qY97LYZp6x3/zzWMTJ7aAdb0BWAKf2uvM
05cOez4n12d7315zXCo5+AsSVawX1VRr3+7EVsvyYTInW0ouiDxsdYx9egp63nvC
OP08Z5Hyv0ZuMuG7oGrZIFVjEqLojJRewhux0gPeE1kCsQ3FEJwx4jFEvaMkJR1w
CqEumWX6uW4s+coWw8jfT+iC0X1LyUmS5XCaxUQlnqjSdD12PHUN05419jldoLCE
90IMwrXej2vstaspb6DbLLrc62dby09UV5zWG6ADS/zZQB/UYdn4UJx33joFIjDd
Tm+Uonl6z5auz/NY8qKMlNhABF6og5xokI4jn2u/kQd/oQmjzg8nP0iG7ef/l66P
LdbQamR7ng6YDRYmmIGcjXSLNMvCX0UyL1b4AnPMdZasOcCn8xdHi5g26BirTgc2
GZx5mVLxyxxuD+bR6ayguehZHQ3c6CiIX2k4sKY02PpZA6kIsDSYTxLQPz2dOclL
9n65avIu7sws7okZe/N2vPx87/S9KfS3yjDEXP6z4D0OsqlzTgdJ5Wz/FyNd4VNg
zlPCbNB4qHSRPLw41NqrVOGa7v6t7HPsYe8j6EGSavnjDBpmX84AFVqLb7I3f5ki
/OwGvZEe4afTqIoWCoYqzv3RAv69lY5qjX9j3zsmCChP6c7jbsso0MkIceCxXqyf
GPtjro0zILzEQe4t6Wg9YhQdbPGvP1k7dBpCZAk3wePMOYf02Ax/WOFthK8jTHvq
aHm3nwnxaRZ5Usan63bc8yyAkWK8n/DRaP7hqH797oee3/tgkDT3L18qglyuOttV
5wLqD2LXKphJtWdEmyZTkvhSmVSCX98yJLWY4ACequJsFy5BNoyv/AnS6SZrMSdq
5uD55KXUY2Kc/kkfAPdt2Dyfdq6YNpLbGag3sUEq0aRKApLDE27gWnNXkVIhr5F2
Ge/62Q7UIaqBwhesf+1asN07PAh4q0IzgrdXQQY7A1V4smrozioLF8QHjnNEDW0F
036Ocgt7GRb9lxYBMRQESvMrefy5QjxLSUeZhc4wvVD96yRHXCqUL/zyimd/TB6m
SaenN/GN5mYWaR6HnTMJhBpZibCVEvMSdd6dMXmV8v3jj6BhQIwX1Y72TOrqjmIW
bXq6EhqZa2gy0TNgscb0p1oJotNuwtFeg0Wf9Wqab7wFKONpPLkk0hSiJAJuSHe3
Ji5SqZU8DyyabfqoIaAUvpGgib1r90Y42+JhjxyR8yt794YRzM6pY8NTTMyWysOL
ZGhdEC/TwYtCORvHv8ju/RaA5pRQ6+fn4MOtxWq/kc2APbDGB9zhVlrDatxEpqVR
xpr6Ua+zQAH/axiXZfLpLj+GPeX3YjZ2G4XCmhDlN56iFcKzd1srUCI9R6v9YwlV
wm5iz7GrsfFIIRSxE0ZZtnpHSmPqBMtXSUmE9n27O9iUxHlgytTSjd9xfqAI1E8U
/XCy3Xem+v/KZ4KXx5UrLFqxD9tfVw/3/AJvNHhTf3+LPDB1JBntMRsTJznfbEdY
r2LTjaH+VpqlaqMD3JELID0DynFvR3+S6k++JrhGv7R4UxFqtG7mVUAkEk0A3MS+
Xt9BvPEa4DYhGQEAQSkm2jd/CN42rxv3sVWOiYfbPqbtQdFkCgDp4PVkvDhDqkSU
fc+PRqh/86sl4Ut7SzYsn8Ji97b2cIXTHaYSBsvgNEoEBNCEeG786rHZbGw/oi5c
RTTtYcc384pLo4DeJSnPrFVKRzi9ZMfNDFv96Y0tVPV4CBZ7j3Wd8MHJDIq88Z1q
TF97TgnuT2Vqhl3cLjZOZMQT3kMfzYxVcMSuf2tJBWizj4P89YaxHEhpT3jCSxN2
Cq+ywOX2pc7jHp4XkB4PzZrPtENvO8NeMZVkbpThlX0nTX8y7Av2AAhCuNb6nB0L
vrBjNzUARFRsiz3ZyiyFXRTx86f7DbUPut1zHwjQf4o55udDrZ0FbmpI58twbJIJ
n17HlXUkb2EtHCDdy1Ii8B0FYM9wYHVUMRHqOXlNAnv4ik4/0YAHpj+JyFbYYzh5
CRasAFnyWEGrM0o6flu9HaD2kb1VfEqvYWS+u2i+tDPZtj7wu80FHdHFOweAFxK4
TS0QJFKTXjCFKQ2fT5M30vf56ZeEaNasURRMeVsLd7e1f604VIy8ci3LLqHGasfS
RLpUHCUCYj7wQBD8up0Letel+0HbaHGnXU3YxdVBszsDQXNTlDspS0mWmdfRAjUw
PP9l1YxWIsSbGR+Ow/7ucNfl8NqwW8uz03CyAOodlAd2apnfmOknfhsSp80HXwqe
ezIu2cL/fdmepryvgs5TBXkvzZh/YgKDECJIlrtMQTCOpI/vFs+NzYizvqNyXoro
HCGpXWesstJFYJV+OGfSpSwrHYi4VYu2JH03lOE4S1uYRnN9JZuMC8X162EiS/zS
hEVtQFBuCbUABAiBJ5HbMBtXMjrbNpDuVp0yRMgpS3dm+J0giW5SFVTPlLCo8v9D
hcMu4gQ/MFRwQx5nOe5sVOP1z7fW5vkzYj2AaIg5H/rHLA34NbjSqkI8uy+nebm7
+Ej1cn1a0JYIkuZyMcgtwrZoAyFzhswXCTQxOg40CPFIaJgOUW4s15Tfr2kTzXIj
tePeBnCadjnvJRmzNhNsx3AQ624UV/pvapzKxi7Vskg7f8P9gmIpO35VybRMkFy9
F5L25QzrmJGGNmyaWdbR4o3FOor+vIA+VMHBzMMZqn8JbAopCbGU6MPk8Z05cw01
5xxyur8H9hSLsT3oeVzECzWrn1iXNOaHwtvhdgfHVvKK3XJPm8nQS2+F8Z+RpWmd
RfOtWluXLrh8HR6oKuQIs2RNEGIpkLR2pvFVnUanbwOK4AJBf4eiplqY8C5DfxoP
7kUgQQY6COEl5hFYMFAc2pcwFSS4x4nmGOkKRiuUxn+Yfcv8eppOOgWGGsx8NCHu
Yg15kba1b/udMv64+UGnR34TbVlyJ+n8ZtmXOANkoL6qYFJbetUZFSEJsPrrzVST
b4RFr307RgeIqAfYjgbE8UaCzDdU426MIVOUK2Obi6uXhc8dDYVCNThY1iLWpZcg
cAW7kh/82AgK/Oqm9ZhZdiHacytqoSGfYaIDllrl9zMJHZx1FVp8R5mjssbeutLi
EivvmRdL7RdRvXSlk77DOq8ZJfcINqL/7wasl9V28vESHtMwtkQ7xxj/qxN2bMDy
gBbA6s5pj9G6DZklFIPVLhwCXPaufqe4k7GotQwnis7Lf8x3F7R3b498rhKO0Vab
8/s1jIQ3/BlL0BurR8q4/iE+0GHR8ejtY9eyE0K6NS4xQSZ1/VXRmRS+WyUUPr+G
UPr3vYCVpfk9jm4iOkXYm2jHrMuD5cYm4bWV0u+vW0BkW8MbdVGFyHfIdjuOciQg
z+Unl0YN/UwvijymbDZ7pm7AuX+uCidCCcsEdjHLD1r1rpyEl22qN56lQzHt0FXS
N2WBMjnoLYDmdWrZjoOTqhToBl3qIcblelcOI1ydhWxKL6DiKESfq8FYWrgo2JOy
1VO8QmjwyhGN/l46jlsN77DwFws2LqCO45cnZxLUooyXRzaz/1PclOoB+0Domzyu
z1q4hELEnOim25OQUeLiiW+D72fnApZLTujLNQI6YsfQjDiGpDd/RGQmsBQ1xwGA
DhR6WsgTjeC/53CLXQRFlgK0y93zup0ZICTrftEKAg3cFmSsydokcu4survPV/Lc
/sP2KlpCdQiGhQN2x1E+EJHbP7vnHl9RzijR/X+7fWiCpkX1f/uTDq7s2VMgwMYE
7wbbI+eOtB34tc0rYZgN6VnAFGKkKaIoy6jb/F+srEh5yyOHd4NDfzcGg3VjEtlm
MHjoxiG5nnz+UQl+0AygTUUh4ZPmJhpzfLzaacJc7nDORVZV2A2kzVDlp17RXAXC
TGXrpHG/pSYGGdTKAm+kHZSrbjDtSZS60owKI5XOT+0UKrzg0haREBqhDua+Ks9c
5n/8796bxi3fcdU/6M8hFyTgqCqVQU6vk2sedI9rfP/xjmH1QqXaDDEeUvNsBjaR
9ZiNomo6fdFYdayTEAs8L/plMoQPAYA3ijNJYrUBnGvmoe9KsngA0ff2NPvze+Q7
elgXjGTpF0lxYGUB6WQN2aJZKdoZ6u/8cAIBDdMStuzWGwxg5hBDKyKW3ztOVTLg
mAiP+JBmQkYPRjvm72gyeB4QiqkK+/k2o3imk/F9+pAbcZOp1CWNhikXw8AGXN8B
t2QyNkfK7eFBBUdk3dTcVtOAL32jAyYG1ryACYap3oWzHXX2kC40YnaOepTJ8NsC
tDGkzCoy16pNmn9M1uJlFGMFx7bnCI2oTXb9TX0X+LiLMEERUP5IaJJJOp6HcYvN
qx9KjQj4tqjHkLB2MCU7fhISeafPv/62wzv5Zre59g4lbFd5dSpXJLb4/C5AVaZb
OKVU5csk96S4pRU/ut71DEv60j3DMiziRqRp5My71XFXGsPIOpfBJvTNe5Jmhb35
fBJlWMrWYrnwiULQKsQOGcWnE6aVOVSqrKhOfrgMA7UBeuhuCPHATkccNH5ZTAm6
bVhzCuviiPUiPEQpKr+cQmEhCJLsPUZBjLgn2MocRh9M+327h4hI8XOuYl/LmlpP
Vuyj8Rg8LJjq/rLSg89qnD3mrOcHWhl6cLXTWIvYduE5lXA/JWgLgEVAzix03DZC
u6MhJafIpM0tYH7QU3t3/vQ+Mu85lAeTE6Fq7skCEH1hgQGNKwmYxGxx8rV6p+yX
6ysuC/kdhgrekcz77E8g95GAO4THPzlgrTjAh2oIFGCIMtCkkB4sbF39z/SJOSaZ
w3iLZX2IZW0Fftf2fL8R8YSm1E804j1K0cv5Ok5s0tAxR2CrbWgo0lGMrNd4K6kH
3/7bTUCTFwmoNBaWjfpBOatkL/kVmNhNoRtsVzzhweEx+CzwSJV7Q2hDSx6jfS5C
zCzvmztRYOjoM16cwT4OUTHCS7pMqbqxOpoacwmRW2iPSf7i43yHHeFrvI+1Nq2j
ZPQVVSNvxh914e0L+Jy+C6f6oap6OT3H3p37DgVcMws=
`pragma protect end_protected
