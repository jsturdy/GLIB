// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pY/vqTMlXEhLsiHtKW3Dw8oZ+PX3HWSCCGrs1UIFLxBN/RKqqkbF+2Fw8FaEQNqv
1WKIrR6Xx+sl/OUIBcnOZvc/2m3bAoIMGHYvdpmVIVGICw3DuIM3nB02Vp7hIu38
XbKdx6Yz58eDD8p6h9YrkaYdtFQ3Z+A/54qegLzlh9o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23040)
ftX+LqXk5qOEqpzv6rFMjp7H55mborkcPcGSbi2sAtm2FDhndZsJr3fnZthklxIM
iyqBN87SMkIMs93n/NZXcJgp5SSImngQtgV2iUOrkv6SQeTSKjYGkrCt9JmE3Qjq
RonOJUaPwiHtQRFnMc5uClfk9vPQg5Nxj9NoTqsgWrRStT+47R9Tfg/OwrcyjCaI
mbX74z/kqOHq4r69BQ4/RV6E0ZsDxWIOHylGK70WTwabmsa0xSg7kkZJBxI03hmh
afyL4WMMewBFhwi3TOccFc8IbBDvGS2qIoHitu+wB6O6MfRdc2wyyLcKBA3n5U0+
fYWfISI5ACy4cU40pmQtsPau5HRwWEX2lurhr7MuliT8bbYu+3X4/0J3PgQ/TCsX
k/Rmvg83E1aMSLCP0cSIi7Wc4GJXH1SGAY3YnzyDGNffNvM2VanuJlX5YvBlIMML
uBN0/Yf687npNtMd7y58+jUsFtUhP11+ZBSGLzseIckoS8zWefjR5AUinhuHErxt
frt5Xg+wlNvcZ0pAzhExyCsJoYJC7tizTes1hQ+5FMq1PJfFbduQncogALdP2ikH
bVk+NrGn/Lt410PHLrKlwLRhJ+dGfm3qO0NqOUYPZ0yxIZkHPFI5Dz3dQpnRxqd2
imxh2pvNI++tkSdp7SHyJ6GPEpOtFD12ExVtHhedUWgBs30LjtpeQKZ+iejkFImw
MUyfx8YjsqeQcvzmToyE/3sWVWWPJsGJHkrdFBXPW+Qha9q/gDvk76ugcx3kYREY
7pBzHsMqBdJw64D1EhPHPpG5rwzGggyqQK0KF5N5N/MAx60coyYoskwuFQIinKCw
2dj1Jgux+1kvuvKXpePwH7kO/JF5Ikfh/oXDgqG+ZIvrffB6wjlkbyVVrsuzfcGt
Q3DZ7lYMgiw0UeUWZVQTO24EOZ6aKT8eM7pgzFcvXfGDJ+7P+e4m2DNWyKyE6EGj
Vyx0allv5Etur6TNAfjoVe6FzcE/5IlzUmWPlr3ziBLAg4ExHFJWA2+9mTgiG6KS
oAHM1pHQBWCJRrBpdBfcL+BtVJEG0wCav95QfOm42vUHdY1CfAuhvuUh/A+LJDAD
dkiQkMHYlMB8UHvvhf4DfQZXkOo+THqfwJgt28kbwUgMbpSxBbqgQY1doNjo+M1v
sv3oRk1XO/pnzw+I1YnOV3oZNMGejz1viaU/vnZ2Vn3P2WWbIxrwvI2hH8zwunA5
Lo71G8TDy9KVJ8ftZzG6+m7wPgbXkk4ha7SxwaeAJrh+0S8/06sDbRvmUqrNkSFn
JBGwv9qu8HvAro1f0Tp5AqBkyPJblQ/bo3djmLZ262rv63Wm6i187lEJ1M4URRzW
t5hVdmj0lXng9QB6pfteYC4wkzKhfngxuuRAb0Rs1XlwQV1K1N3u6DMC7Vj2rq1R
baRtmxwkocyOZgfvvyFr8mlYfZ/satTXTspUpoqRZL8nECgmRBvUlBWuyWgiFyv9
wZWXDTWMN1AgAkY+ySR6/m8LnkboIW9fQGR+hHD3B5gJbDu6DvLiXACFeL6w4GKH
l9XwjSiPA4q2JOye7lVvjo6qED44lvgqI2BGUIlzPnQXFAMaLT1oE+KAbsHpYc7R
uQKlrrpVOcqohVYhLTAYBAyWxR7HUgZ5YCxTMTWmF4zARJ3ibPFSlQcwgL2FJ+Zx
9xRQDHSIsh/zf8S4ymakEs4asrMbg0AvaMKhnfdn9A60j6LfrNdaRudOkLlUu8dM
kmpRAx8VsZqvRcalmeVnql26zRLfXkQqiSoVwudtcIq7+TJquZobuiNQn+kKKD/M
/7g0LZngjIVW5Y0SuRxT0qgGBxJ2a+3cgIqwO7sI48IinuhnaWzUS0NwNZcOTZmt
Pcw9o0Rh8TkxH+BV/vSB6N3C3jJDqjF8XDM6Eyw2Ov64v8oCUecASvyU2CAivonY
u/OQfKcBHSKEo35rs15H/r1/6ZmLS8rRA6MyjwjAHhp8NgE6XCbIDkC4dVc1TWPI
0d0c+HT9G96qQK8P4WD2W/tWqtZJ/sgzvkQ0ID2u0nQtUG+YXrDSA7g8g/D6fvoX
NB6BKqidRuS9qjevg9Zow0+ntHLE2xNP24DQJdn0Fw8LKbPLAUwkXAqCKShzMlM/
p9jJTUmWP+qVc7JAwWOim/E/R/Fp8/3jDLL9GkSnZR5ncWwVKfm6bPGuP8K1SMVT
8I+22X21Zo/wI3y2Ljj+Pzxbjq7w5BryCh1ey4cb196KZRuJ0ljAuG6xXF34ga1/
fjMXmBujKGCSjAqxbOSsTqheeDcJNjym7Ju9EwTNAipaUNQBEnNHDac+z2Nb38lg
0BlyL7PaBgpBJBseIBuG8NNpa0Ss+h3SfJrerniK9HGgdC3wStrwPo4kPpzPcZ1P
0cGoYShnYCfWabA8IKbPG3GuBU9NLHY494oSfUgakgvxBocLk9R5EFAyVlkSODwa
WKb4DsdAW1c2wOk/XHAyFISEEFCOooNIT8OmxkCIs6yXmIi4yLVNaqD/kiu3JW1T
6m+PHEx3N1JGLzobtLB2/w8C7m0no38BAI+duNM5skcqui+SRd/5SGm00TRJNxxh
XFIPdLxkmy1lbIIVUkCz9uEwu7zrgAtwPkmXFiMP9X9PMqDZBtBLm1smogNuyB+P
s6bGBufaXTIzCDMoC3sLEt2tD8ibN8612XAjtwrMyXZvQNBYuewAwrn+9VGEmE78
37YIDhBR5aqCm4UYpS43WLojDPX5kTS8+b7s8DwTkbea4EgsDJe5g+FvIOIC+AHx
X6fLNZHvZs+9nP31QYto3kGt+I36xq67CIGXVvFeCkqsqyDUYHtyMm3xNMUKW1+F
XVZziMqriy/6AyEG88fsKxmr2z3qv/ZRMnoDzwJBIzLxEspO1CYnDHTs2ykhdZg5
xkLUmO6xY2itda6c1ax0/fsho7MGnC4B2fs7SgUd8T1vLFf+A/lh8lCWHkumWVKe
TOesOw3U4KSbQtOIyNoK8WBMdPG0NUsfIkitdaQsT31g1l9cQpOAfolnR/haXGxm
Qpc7R/s2WWZYydSHNMlUpif3eDJNzMtq93hUcEHWbCXw3k5Cji0xp52vE3q7GCWR
m0rcGX1liLFLa9KKwJEhn1rhhz7V7nZo1DptDHw8FW+Jyne6iRr5vAXsveu3hPEo
bDn21Avre8ZZtozRTvB87vihVCzyTdpZ6k3pfpvhyu1q0CN8IsLc48BIX0TZezjK
aWTay7Cy3r2TmID8xjSQBHGs9UrFHG+3rQPuKpYvY+dqdkozG6S5nC9tdpJTCazg
xMYDSVYBmTAWZDruPQ/ZiIc4fRXBlIrhrH12M2bMNydielIHSN40f9VmhngOeY6S
3Kaoo9TRVQ2EtbDBMFHOsyo7flx3KTzegrFjt2IhVJvn3ggMxpxxGI9JyHzICVhC
ubXFs0AZV36pUbTcF1O0HJ6Ncs+geC8RQYAI3+E+2cHQODXVdLvQ6Qq10fGPIbLq
cR/gf7v+jTulJmE95aZs5InqZsWDnJQVuTI3S8HGtibYxAfwwBYqEMR2pu81kBOr
pTsLgBfYqDfCFz9pjcOHaoRNttag6uVB6VkP97jwJMqt1VZIuGlgLhYkUFAZiTUn
rsMtHNZeihZwFhgP00kHYDC7PRJc3laIaVmkDUumMZjbbhVuciqqYjMlpXdokVJN
/g3N+Fzz/NE4D8smaMPkycCKdv65jV67UqKNFEF4HWTfNF8ea+hMViEFJaurm+Wn
NHLOOoZ/xQbUc3K+Z229f7T/aJ4gmVeLSgSxnvZcGNi8+gwN/ozNdzoibyGjr55N
sj9sD0VeiA3z6vRogfISzjNRLa/b3EzHzLVOY5+8hlqmVSAPTeqiNdQ5TRqxhxyL
JFfN2yT7q3UwSB6sFUqnvax7pkCnf/K85pzjn4zh6ILJfrQf8ql3TxWW2dpFTBPj
DDRsRwymeSsT8899cC4ntA6OsyvGvqqGBggHQUCGVNEZ9FIKLvVoc95MpZbn4dRK
ZGHDJ4CF6NQ3r6ZwtcOC8mPYwFz6fVMoZKpXPK4VNTa/3U0RqJph4kSMVxwFzgq2
Njn3s0cpwKeOdgI2DIaiLWp+nVM/Nt4vRBvwYSXykJUo1l3dCam5keFdzvHBtgjA
h0A8MsHvsI3JlQ745l6nwczgjeyLSfNDmr2rpPNPE74sEjSOa41MK8gtUTY7dgm7
oWzHkEOTJ5mSVJtt7X+93ykSirOE6eH9zj+pmRbu+Wsopqg7v/cPtrwD5xfnYjr5
ZGyEdHTZ768UqJy02+lE9ErIdyRRgz3InZOrn1zYzpNGbgiEoKxv9ZVummacKJf9
x5lQVIYGhOAjoxBcsWfwl09wDQBEqVONqZy4NKPND92aCHG89p50HThD8qyY1ZnP
Fk17LYFy8qvLCLD6SiYbBrXmqgK4UnE7JGNbMijcz/RpHF9EYlID2spK8C4Cg1gE
ghjJLJvWI3wscB/zM6XweNvXQ+wrbTBbpkCOK5D0CPbNawffUtDNNOchFO6tARtn
n87Sx4sqmzRoKDnaEIOqNb5/weQn9hpwgZKkSb/S83IaCBjWKaLotbZ4yFC7bcOH
vSjX4wt1HK6ddJKgUWW25a2F8R7FQy5pZ1W4eTyLk5nZB//V7Rc8ejXFSF2CkQTW
PXhcmIWMGt9t+M4lzK3NimbzLTVVW0Kv70RQERJyi/bJ+CCmdKGgjXvt+X4Y0Pfu
lOgxgUMeI+OI1JuyLz4u/mLhaJfTwaHPMMIVZghsWVXxe8XFpCmamrzqrH7vScS6
PJGtkkLTEox3xlVy3lV2Wlpq0afWYHLtsZMmW3S2Q/Yy2OVEbtKYmHxo5sRZ4WHd
fxUpTnfNATAwxedtc5Kk1hsRVKFWEp8l4gnAlaKIZLRiRFRVr8Wt+PSjteEADNLn
1NtI12yID3UQR6hDoWduB6/JtzQuVKS4MFy1+B0jB/gr/5C2K6zOxMuphvjtlRHC
bVsmqGGV1VGUZdg7eZoM/Y3njM7EPjb1JTebUX1ChQBLkGZCMaKNPeBgKTqRp8Tw
hIfRGCDN91+CB7eDyXV7CJ3KMfK9ukEyNW7B1x+y4cARS8JgoB0NHl/Dmysc2sAo
qfTWGYeUMebMYsL+jFbz9kytQJuCRF9/pOO1t6HM0UC2uvvRjRL19gp059zC27K1
8FVSPUFjp8NF88WBxZK7C3MXIP5QY/80Ovad67w+yPk5VwwKj/VAJm2xyvyVraz4
WN9QW4OgQqJVnL8Dd7piNrsBWXfgvZfkJnTXfapQSmzkmpbp2cEa2gfEVtbWsyjk
rGb0HtALM2CWZPndpUt95/NM4NLXyqJIGF4logJYqNX72whlF/VJDhzj8b7mkSz6
56Rs4WPuwVdFF5RgVlIQ/WhCXxyo8P/qSTXLArzyaHhMuX/HpIsEVk4S1CMB7deO
TNYtNLw2CI1OPSYHniWva9JSDm8K+sv5cL1UwtQ7ZSGM3pYxgttlHGoti+bZgbdm
WhPUV64EvcxXKC8J6t0lTqLI/m04Yxqwgt/3KXkpE4yOhScWP+OS23voV4mYmL3W
GfM8lkWFZl6tUMmbzfLdHpDHLVhyskyXrLpRUloOWTAvfRB0YCdCwbslhBMRMcXH
Xiq+BexShwS0Q8bLeFXPgr8ufNYj+jipNyAG5JmALBMle7wOBo7uiJQ3R5uhsid9
vU8uuPC6uOd3/e491nADLPCBji7asETaPiEScozF3OHYc/QkMSTRGzr75+Fyj8C/
S02vLX+OUscce/kCLBpiRxzrWtF7xAkn63s2uO4dlsJahq4O+p4i0QTv8uly+c98
D3cNimgUNy5vqWlec6BC7JW3231d3ueUcEAV6URU7u4zsCJn1JXBe2u4KuKGxbmq
nDP7IO0fE/QOuO1vjaeN1bLArmo6zYqgGrT9IK2qLZnOEM8VokyXCzCpgWpj61rv
JBszo0ozRdo77a8xMaW5obF3jUz826wodmPJ2dDgj40tNKY+avup4kmPOl+OqiHT
WanMmeL4jFy0jljDkIcqPgyG6Rp3QW5CGHFkCf6elX+HQya/YH3XNkd7amBozPgI
8ysADPS7cb/H9Gkv2lPXO7pWG4sOCcoiIlVW07dO7ZoRWOytai6Cuak7ncoMOt3F
qjWaxWzxr8ZCew6dmB2pcdAYpMa5RThN1DmWXU11+eNG5aUOoFLVrwdX40h9PSpk
ECzg2Q2d9L6UKwvK4wi+0yyzBpTuytbZr71hgmkUNdmZw1jiAuwdqkLkj2DAVOHL
r4tZXhzMc5AoxcaeuauII1gStc/SPFzeyDAOECGxbjPn8W8sjqZA3Tk/H7tz2Bgy
4nJnc9E004FPvN/5gysXxw/el7rJjerC29JCFx2KphsYPb72QBHrHCCcSPQ1TASo
fiA5SS1H/5nn/MWoS4pjHXg8cd5B6dMnmDFj9dMXmdEba5NqXzbb1z71DaS8aA5E
IQPSqvIPZ+TYYCBR0S3+DuT0Yz5w6v5AydXZjeMGuszuHr6fdShLBfHa5Ui6Q9hF
YjSPjrhzFRmlyFnu/lYwRVO11N1bVksI88b9TaCSVDUUX1GNyy8lYVzg/7rf8kda
C+9DJ/GL3ZJuZJnpz+dfU8F7MzpIMJRgb2Fnp7EcN4ts+c7zkJ2wVuinpPbvvzt5
T5Z+7aiGseeeu5fK+XlzVINznY5AWxRJE55zKphp4oYiqe1BZn6VIj3wGaLlQPZc
PlICpiNsV3xbzRvl8J/C0/qy1wWn7se4o9OgBuB1ixBYJBGxStTZ6VuK72Tp0/rh
3pmB0iCyaOO64bMXDJtn1EMbfIdaE+5WQR65bKJ03UNP3UMmqesAZW43q6/HnJeZ
drFSppYeH/0bLtN3Z3H0dZ9CMSYJDSYnbbiGIX0Ct1lNb4L49IZP+tXKCCWSW/Bf
0CaFXy4VvQx2b13vhiVplbqAzgW3HbDt+cPNic/R3SpPHzBFwPxxVnzl4tIz0ubr
cmEyO0Bml/6stU8k04rU0JALQP0jVqr1kUO5a7QkLiBEg+kOgvfxv4yR4AG+15eL
VKU81K4aUFD0QWimBt/35p6JpNNYO4kE//efUCHmarRklZc47lMzkSQRhHuOCPwr
mQIZEts9ZJUyB6qFFwPhSwZV7eOPqzV+frOY0V1agTetnDM8a6DXnvRMKGtLy597
K8LiVXzP8QVlZJ8ZpZJNc5S4jK+rIHgNBn0V9j+gsf8gdTKRFvQmYMg//Uhj7aec
fPxjj+pnqFy6i7AjYMqAbaW7l5B4NHktejPUzkgQDttSOmi/VV5+U7MvQisMYPMF
pQY4lk2PmnMJztZPkBTsNm/NVuzTuoBO6y/nvaAxr1QnYnnnlvE/TpS7CdRcHhh3
ZzMPe1tYX2vyjLsB1HKzrodBE7BezibRTEaBNv0Y/Tx3zeQfO4ZPdOdD/UWUsFUh
9SjOXXFXAUJvKn04zFgiCrCQ1lSRUj6pOVbT1g4J6vc4/ayX8G6FBFZ4SiP6/MyU
Mk98CRTCpnm7mHYUC0QMdU/JTNX0ti1j5rMUz9+UqR1SW7JEP1R7syt9PGGDJs9V
zPTB25VCbuUmkI89I92a4X4Bw1yJ5bNOnN59K1vO/NWNbXe7o6VvL81V3dM+sLxd
RL9Q57kaqCy3b8MYIwZ2QoxyPXxl+8YDpL3GIRCeUKHXOIO6V7NArDSYEJgsCXvD
uPsJy6yo6FnF5Ieih2yInU43CEfC41fxE4AF5TzoaIBDDBtA6noVUJhQ2kkCmocf
nLlfsslAuRrUnYxIqhOzixC7iPvueNkEbim4ZlsSOIRfyBZGTIdxpcn0LeAc+Y+8
LuzwTswRahNmvrOQc2xikcJ+oJiTtBDyOrtnVhBNALo2/SUCrXQb27hSwD4m3gfX
pt6EymnsM/tKF82LqFVT1L3rE3uSavW29ZDtHckWXjQ6DQN0yyayujn74KUlI2tr
mUeZgHJagRFvwyE4NFydsSdbAUp193bnq/wExQaUvgO0vuIn0ocN8crK0bbWleej
Mn8qXo6mS8/69OfyqlCsMrXwAP/k14W+eqKykts4XZZwbGtWkTPx/1/zQna5wuEb
qFmbcB/8p9dM/Xi+iXOqPxVsUEthCkgdbPjSMD2pvLu9F8Otuxip3lh4q6K8jhS9
xOlMzME0mv+nLHQxkxA2BP/ykn99Ss0CCmz6EkXKiJ3WIaHoD/2AB/x+RggLpTbL
guIwN4JNFovYxuWda4zsskc3vRbFayHtZ0I3LSkLTcgVo3m7cv5g6VxPIdl2F372
JdV0ZGt4wEj9KyDdIBzPypKjxBunS9xO+5B7ipuwlofl5hx22DCYOfettOhE/pzY
1NzxLYSsF3t4XQH/noYC9vHUXcQLEgTlfcZQ7eQhuzU88sT5x0Ue2o4mt24YZHK7
zNl4T8uEmRryexmJJeOV120j63CIm06p9aqTcBJ4nuv74ayhVba9o8JAmflCDHUy
55Xi5Aamn0aeX5+2H5JhozxSDb2jorV3kOSrfhmh66r7G5Ayqrrq5KXg7l/fouQU
HgvQv1kXA7ojGFgN2O1WedBSNg1sH11fd6VTJN+g+EpKDGKMMGFi6yj3DFbrtY2k
XCGKrYWRA83orCkD9/TY43XKGvD2+w4uwQPmjkm5fuACw4lD2XbECdObjqw/1bTH
C21GcW80aI0DBhrY+kMYtsoHBet2NzJjWhelFuVkYXOZ64n8V5I9/KUG6dbCdmNi
unBhcLl/BI0MCcoAMPEwsGsJeiSyQa8N2YzuZghaQ3wjzVZ8hfELxm44xIbJbZDt
aC3kHZ3hKiPv4cg9DICW6HO/QWXwcaNZIlgCQZi7W8KMi2xLIs3lz36mmZ7LBkGJ
ptD06grZxl295J9q4WdR1w4/hlxO8FLvDCuA1wFT4TfSfKw8enaDpBsBNekY0U3Y
JW9pSSEYhtzb07nnWWU7tyWIQpgAyMEvMYeFoUI58J/tAkMiQVpkApMK2c/gUBl7
B2N9k/AEL2uxYPw3e/ykqzUkz3tt/7yP8P7YqIQiIj1bGky+Cl3mbIOIrML48RdL
HkiBvcPt23PZ+dADVviUrtNGZCU3o18wjFXN79s4RE7z8EQIh+7J+q7c8qedFri3
jzx30nleZRJWsEnG9OatmJslQsL7YUXL4oUIrZRkGov1zBLuDEkNNIFLLUUUPs+F
nKJu0ZwD0KJgs/XhRholnIUlfprWz8xH2EPF278i2zMAFsCi65B4cxWUnzmrXh3W
Bzi0S5rtLqgKlVHEOegxtTPG9E24KCQk1Jihyyf+r4j3ikVQ8WSBwEy/BWfLDf9a
bXqccWjt+o1MRDhykmeNjItgZPeA53q9i/B1hlPGcM9RZI4pMGrJGC7DgpuVTk8F
l/0XIMUcOMqr4iCFfkZavTs37u24/XpZqFPgdu/W0GnF8o3cjlxKBjiJvKaLwuBR
7AUKbvpYHvSYrmTOpAbt7JFYYKbRWI+GgJ+kcCfvC/g7Ax7CKIShUP95aCTNFhYZ
NMDIo3f3jNqs5bDgOQXiYIXMUmzSypVQ2tKj8IXcfsIF04rnOWtSdIinL7Lywri+
A8B49/V9QTylRu0WLCnEDzrQ4TTxXtb5X8xLAEx0dH4Q2X52RTAd8FV7kzHJQvsQ
rvrttqRaNKT758JG3uez9MRqELlxlM7oq9JZY7PPvWtNTAMS0IhO6lsrDHsyO/NF
fJQQugANn20oQfNfbSQ88GSSKB20cXagAHhXT9Dgz0cPDt52rlZ7RW5NBfb+5ZCL
AxzlhFaWEfVrRHbmpd7V6PxeRbvVfJ6qNcXI1cNZzIpy0dqr/NMr4W/7YCT76X6t
o1IeNcwUEeOblgCFLK2L35BRS0R2KPKu5FvGGWw52q/WiTin6DPMJ8KFckO3dbCe
fWEF8PD/vt2fzKiYiI0pSzVGl05FJhRkuUQgulJnEGhT2O5aKNMgEa8FBJl8Rp7I
4lI3QEI/wRoDlXxacuGfLHOw7CQZ2BK0rqqG7z/QgunHxPLOWmB+8A5xFr4Oj1JB
C6aSBy/77y8ZH7BBTZPWv2Nj+UwzkX3Jc9LPHHmcEBs0w3MW8PLPtc0cKyofp1si
OggCYVB9cZ/VHbWk9aB2vgQIpLFTHO86nSIT9Mcbe5ju2EOtPDzXlxynMNmF1KUH
82N66thv63mqsELS9bq2Ltd0/2V4dCt2Y7HZIt6whl2WQos7guhGXngWsNyDrDdi
s9+aqihQkm4O/HTJAKgWwoi14bU9C8kg5UxgQM/Lnp7Rq44oK2uWCtcRiaTh6uDC
bVcVqS7+7XEFeKP76BQauHMkbWgNFytGuZF+KWs0KEiBInL8u0tXS8I/+iJnMWNb
mctxXoNMjpzG/fraLFc98nhx20udW/Hs8YR2MlsGb5oRMwvYirkQNbhF+g0DTuUD
R6uHymJF7CMYvcy0jdGQDaPtEgzYKUizgd7twlm+mcFsIjx+9O0l+wKoWuHgUx7x
MRULoz7pHHFVs097ysrVM48mzAciWZVbJxIVel4sxdzga01XjWsJTP9behj7xNjb
1Oqte4T6WcleGOe3rjtqMX6HIICWFPdhU6SnY5nm4EYBnthki/4YSO+iAXAaQRfW
QnZX1lOsjLP4Pc92QwfTRjtuBwTp2K6mN6yklbL/67/BOkezKrGUaEbsmue/tFx6
BauXkcsiDgMeQ8cNnRUA17mhfD8gzaf9sjTt2e4CCuSi4N7nZ+GzkkEeo38ZKcPX
DlmH4xZ5g0KvSt3XKkYknhRLHSkRsGFjoLfAK8FJntuOokXbjZVgq01hd9vvUQrT
XTSORdHcG4SdbMAobxPKdCeUM6dV+gxqE2zxhlsezugyzDR2YI/iFq0tVwDMHCY8
w1CCDal6p9NrIfQS20gMV1mIFUemJnHYKJEaJeqcl1RjI1iGxr+Ynq9IsVIQvV9A
U+c5CHHUrHAUoY2bGo169hmhzIusj40cOAobDcVwadQm3EF4XvQoO8LZbr3conIh
AzdLaaH+i9cFyvuqT6JKy+KHZ20R+O79Xl7gjlctsStwT/oXURwMNRcJsEfhQDMV
d4uzhZV1do/82RuMYbVjU+uHexlrroU9KrqrAY0vsujsVF2owjL5+MBBvEV2Yb6O
7o1XTbzFyCYdPzvkrnt599Cd7tORU9ohltQyK2/dYdeRdhIzKapkg/mB/SGD3Kom
5Oh8FvuSnHkXW46/TOAGOymzpddxkiGA5PyswB7ZqJRCyZXic21y3Up+JMffdmJf
WTi+6OsQQkonnwTAEd7XpXvOSRJRY5Qn0ArNxTcPJqbUTiGanFRmX4hIsFR1xoMB
rz6QAMkBprIdzcEG1ETqHZRWV5jD3BH6dZUHY4G/cdJc2JfW71D427RM0bsrkHCn
e6wKB8NNDWu6F8l0ZHVA9N0AS2oq/yl+Q1lrCrZ8U8cKr5DKi9gqodH6D9WWEU2+
0iAmfNANn2cC7ai6ybqbfiIiF/ZqSmSTZOUdguy/+6G1JoMHWfeakGBrM0schaWC
cjjRJQOPJ/yARhgGuq4x5zV+d8D4+7QHcu1FeSuFMlmXc1ACzynBv9loOJtr+IWK
QddwuXGyD5lUNztqLCswCRMEfGxFMN4LavZareNrG/pBrAncKdDHseti/9URjqZZ
esjIuq9vZWp5fHjugh9aSVT2huLg4040TrnhwyirT/yNkiStK2ZOIquiolvKUqP5
D4X7W7ZW0gnjD+eSJcpE9oJL10+/ndi2tsV15AdRZ/QnWZcz6Rfl0WQyfo7WyaIt
6Y1ySKdo2U3LQPf4YMdHXw1YlxRoIpGAz/5wUNjvGZluTssUVk3RccvGAqjWdPlW
SOUnmeAqwuvtKL4IYn+qb10tTdETbrIvnanMcKoFUjk7+65GB6OlzwSbpoxYpCnR
Eg9HoHSPCsKbtKs9a9swdvUpCsO3aaZs6czJZoSRK6i/sd956dEAiIPz8QjZMSwi
sY+6LOST1BLpChBQK2xOAk98dYDwVCBtC1/tAbPq96vnsNCj8yu5+dIv3XAF7JlL
45AQJ5MiBwMDmDuCoJ6bVWwmQmWhY8SsMF2tyQaFZV1igr8zOHUnEkV/9g3opbrO
FFOUY0ZtPmS5tZeHIDH4bZPtBibrbrgBQMX9VllwPletKwefLSUYkG8sLkxkfrkh
KLdVaYblfRc95xYu4VIh1jizP3GB9UILwT4Z7sfdMXo0cT8PzY4TFZTx2xRmRyLh
AjahfO6fgvR8fRvOdUVAsmw+cIDJvSKNqddakySHh+FdHzDzMnVzzSPapzB5sdwB
IQKqAEesKFG1/SJ53DrwzPsWINgb7hSzOe3uMCkrjEqQbFnWNwoeUaZ6FmsK0HOA
kkoQix6WPUQj5ajoPeXkWCX4vqKQG4BUZ3Lceurzz0TqTISFf95ukVMRgti7SdNo
mL/n3njWtkZYim/zsDDJQSWxgUqh/OrYex2REB8zKXKii5QBoiThnBRKabbkJPKf
kQ6w43dnZ2mZPWjEou+w9u6hH1SeDe+JxKmC5Q2YxRcbnqn7Rlqz7fEoCJXyENOk
ib7aYfV+C/HfkMJNsCXpqUTkVQ+xqwEcHFB6v4njKc1oFu6Zlmt5CWcPKC4cB740
s6ji3IQVSuAwmA07+Klfh3uZvrBe5DB/AgtW4tpaQZepZIPbYKLevXfN6k31fL6a
GfDkuNztZCF3UVo9vZch6pDWV4nFZgHLTulTqrySkqd+imt2QZLj7KOXtFZo5+dQ
or3oxajmIrodhqDtSrtIJGhYTCROHG0xMgX/SK58k789lQ0/5RN8fkb/18Ax9zJg
JOyF74ExNVGkWmwOWQTxv0aUHZDysmOW9q9lb49avsvF8IzXqr80WFM84J5iyDrW
NLn85+pPeLs4HjGQXwm9hS4ze9MruPfMvzxcA0LxA0J1HQcZpwp0pMahS+2FJEy9
A2QzGZD1iri0uG/KkHaF3SFjr8ObRC1oz51Ad62kmbMjf+rPK5pD/50zGNWoC/3A
xujxZTmPMOr8XEwec5vW2HECLxj2oAp80YgFpqnI9+pEyI2JTw+Rb9dmUCP96vXT
+NDJx49jBbiOaii9UV0V3Fxgr1NIst/5boh1rYs8fEUd3SNZ2np6EDFuTeD/FTza
i7yzuNLm38YTKkxmGoJOlnZ3eCzDp2tkmm2FmC2Z7BwsKzeQOnzO+2I7T8afJElZ
rFhkJGWpyrwHteDEaQai2PIZuMyghKfnMkm1d8Wted5dEveFYHLijS3qUV8077hd
x3xT48H0TMaGsd0/jPFi3zQwPSqOnuCuJR0IiywQA/rw+TxG8NqoO+THiSybzJ5c
LG0lapx8jIlzU6EqCjlQb37R1TI2UBAVgbejmDzyWLJrCRhzYzQPmbPcI0SnLCdf
zga2tnQ57rwFQWlYNzQ4zUIPE2KsoZrimqSV7BbRRsvHyTdHMcnotcmOngmsvq4g
4oHqx4FGCpfN4IHG6Hm6qAl4SpydjOnXUktxUAH8/V1TKVtuCd9wcriBgGWBOXpa
8djqvC1ED+Ix7CyiTSEesBNlW3WRB3Sy/FJYtewUwWxxpB0oMfSB5teotfNm+/5p
QHQShHAbXi1eHVdJvzZ9s0pDg+eVZceo6Hn6IdgFfb66wEyDS8QVPcVjfpXn7CYn
cS7UxrlxC9H4/pcPln/2z05jT0BgTBXTjqq0SUVfT91HpNYnQdRU152UzUnAVVO4
AU3EGtrce9KxVR0abxo/ex+uBf4ca/wwyMOZr2M6upCNZytEH91b6zJFf9rwIwPS
5MexSyYQcJKrPdh+NTi84XD63dfq+x2zyQ04PQTtWepHrYy4etDSem1uuDUP+CRC
Tt7tJISIaWlzQIrAr81VYEdU04xBBXLqomLbY2FlzrqxX6ygVicvfcoPtqpI7JkL
yU4tnEesccYNoHjjW6/alXenO9Hbslx0MTLZVtB6nAhdYf+K9r/v3Qy/KIxCbLzY
YlZF8OdhQ7cuyX6Q8xy1/0UnIQO2jQb4vIoEi3XbB8zunjxjTYoqX8/oCxyBFm5O
JitG9eWh7+OepxOwrNcYvoAIEynDKYtEm/N/deYUukbp9Ao4ufDjotyAymFGJryz
RflepjiiHY6655mvfTPyVNhGqv4wiZXUJ92vmtY/9S0nN1k3GD7z7ooPOmK0bbV9
ApOwM8svChrmP8SJovrUh6isePKRlFD3aDfTdU/9DV7K2FCGSJjrtQS1aJUXA6DA
PWrM5Ft62hKFdKdXJf66gS0zFRTeoTO24bjuvc9d1xNOeTEWBsBUasmTDwjied4b
t1ZxQkOpd/u94OnV6Ksh0v0hIG7Jjggs9Jxc6lahe5aBZ0DkFMKfaNZ9RCWhLB30
HPpGw5VgcXWX444/e8cgsAJ9RcpOxozNg3qCnmqmDsEm/2PrUCVTL+7BahPj8TYv
vTEBMapKrLokK2Y9yFZXXLleKgc6HVxhCVfe6dYrZJghS5g8dXonSiK1/MtV/jsK
F18wlGhiHqnBf2hGePWZ9Nuad8JG3UnYw0NjGc8xBX7BGGaeu8ySlILypyXUjWcY
kp7mY5h6vTymVWCiTkhpbdxA8RRRR1G0GFismcjIABrEI24mvkQyrchritZliuvt
lrQqeCdn53lEi/wbntLi12yQjHf6bTY+W1N1SwQFBSDi9QuOz7b9YOOkxv3c6o02
zA4PKM4sbgKrWJPFHrjcdbGPkSXLmLnvblqxoYQzoI920sZUWZStFeKIO8yf1Iyk
iUt1kGB2qDbRo2LbtFeTWWlKbHGeGhYY2XoUL6EZriv7UIQ4CIzmyVLBuU7gsKoT
FnDsUC0GJuVo7x6LQJ4bK4lO9Ycz9nWPDUuxcwIAMEqVIi0qF9NOI3Ru01Enqe+w
pK6VTwxl0uFh9DrSpeBGzFh2Bd8JILftBFmFNaPbeskTOf69NyQQj1ycXh5nru6u
Tf/CritWAjh0Xkrxlh8frSs7a8dlFPmuJmISbz4t4+gAwE9Pue4vhrmEf93fPPR8
cZb+VRAv0MBDdKR7sc9YPKEALWyYuwDnpZo4zrVdkuOg2AFqbp6wj3mcudiTZkCO
fEvEHxe2Y5FsUop90gkf6XJuUmiQqEOrYhDvJZp2qU7y/iM9v2Gvef9L+GdaB6uk
nFEVL3HWDrzaNnqYCpnbDdS6EvURQ6wL7c4XJ6nIuwoRUZpmPoTEH76QX2PVyshg
Vo3GSQVSI5Ib583EF1HraiU3F3vea1CxSp686baDkHWFJ4/yc7piPRUZP9Vnfv6O
qV7xdfDCIy3iQalB8cnWWATCPMdrbQW7tMINO7EtNf+sLWfOUovSq0Ly4AG4XKO0
0Bi/oNiAGbPW4tAecsiWnd+E9mBr/m4HwS+rKz0np0D+WI9uYPLbAM4MmSSzHEul
aDNeUxHZKrgMf2rIXk8D7v9TaprcG/vXXlwmhUHbUge27VZtnDxbfgOENcXs+7kK
EerGMKFIHJgCK9/HfSjd8KH//hn5I/VGNo5FQrY8UgenajPcL/RA1dzF29FtPul0
0mfMx/5v74P4fZ/FLXDJyg9xPDoQ3XVJGZDb6DRrbTeuNbj0mtktAIHDWoHM+hCV
uhdCGJ/WKJq6Iz99e+TFeLzyLf4SDBMHgf9i8aaS9iQc6m7j4VJuMN5F4LJTcZM7
sKTFBxkaTUwwSzW34o3gSCwJvgPkiUc4GJZkTYg8IQ6hGE8HFh/bObbA1ctCk0HS
GBIuvceqnnJHyd0wYAgoDBz7P4GX4taZDvqTBgeKL1+EwI9Do77u/9Jd33GUu4hU
c1U4oZkWpwWGkTowZ9kYrkCl0gOcM4KGacIDC9UmtS4u9G0slCmSRahc4sf++9mI
tSJZAiNukLh5WrI01sDB/BPsc27ZgPNqdLhKWJImmDPhTxY7XI1g9smBURWhoStl
HzXhtXvLdfJT1vKS+k6o196SpI15oSSeSXZqox7ppKGfdDTgE0PPo7aCHTElecJg
TCcZd8g0yMSOZVeeZ4sd4hRdKngRLGpQRygvMb98UcoRYYBjqm9MemzxkaBTm/7o
U7ayDJEvoyJqnSxYcyCgnSbvZGkKAJQxHK3NdsfXK2JT4VggFmefOwu0heUlkgHv
Xj2sqAw9dV8n/DX9UrENyHGfo9nH4Rt8xqobRYcnm1m9zoPKTsNiVlhb28V8M9A4
uUXVxyCg3QHvrYZQGEcEdSoLbPtrVdr6y9kHo79uhQqeM0LYuqS6ZDxDSW8NxON+
DsipAZyVv2H07lgrPsDZ2uXBGAOHP92bz1mzG5Bv6pQGVslsQzCwiQSLNZTbAdfC
xaTlXwZpf7t/k+wF3opotD2tEeF1vaxrHHJXDZLGziEME5jwnHIgm4jeGdJakfom
d3CLuV2t5sh/81LxzLCsSXkmhbFx1rM++7uvMjrmlc2tPXG3+Kfi9fR0pcNbMfMT
NAMQWuTFl2s7iZ4vN4xHszVLL/abis/8jtAAWZYoJr/IKwUBK6rn4W9cVErglIF6
tdFhMOiRVjoZWt3AS6NG3fFr4F3MrRAAR3ung2/xNmepjcwWjbX+/EQeE/1vELCa
m/I8CKKjrYUwUqvYohdnSBId8Ca1P4B4ybA7CoSzyPbPAGlqSMIQaYUuorkFPjIp
HyyuZBAr4iic9695+eiuVv5iKK63db6SdgJ50SGWLAbcYiZJqA9H533fdaef0rQX
ydeq5xsNhBswvHgBVPOpp0/KGC/ZhLfbu8aaOadyO8rgyeXwCXn0NMzZOilc+Qkb
uTTjLEGn2/j11WA/FbCA8o+T+ELZT+EbGKAbi5wCL4nz26abM2alqGgSIQat8IUX
bTX1vXiVaJe+3tSnCQ2Q0pimZbTKVmaNqvt2JaPKwt63VEKJ2AwvGhrTEjcwLm5c
BWk5QXFR3aaFn8TtOc8V5N4KOcHH4KkCrCyGz8OyhZ/rl0ESq5YjBIzvnI/gLnY9
7Y07/to9rbaDh2cddmF1iqhf0gZwIg6VV4ounjqIsziVGdkoJLV51uyh1ijI+zpj
Ax8fMxozpAHmrlIcGjE7han0jxeIhUOHi3o/vmYOFst1fNnmJGzpBZXpB0zOcKLn
PQxZZcgRsi3qp+n3eeFunFjkEXcHYydyxujL2/WJtvguX3L3oOz3AXW13bWLRavy
bCXFYpGgufEKaYV0BwbcYAeNujyEmd/kv8Lke7gCleM2GVj7LhIrnY3cXmzqxaha
qjMffV9iM2q+DA/NsgScWOAQlJ/2MSm2gdb24Va+lGPcXHXUlL1coKZ46SrvvMHD
hBzTsCS53w+figPWvG1cHZoOe0e7tsSH2XfyoaOdlY2wid2nSzjX/ig5piPr5mfz
zn5tcGzCp2A6tOtHTa1uUUO2+cWeRJADZ2qIZoVUU7JGQD8C7HkZubuQd+kHQw8T
cLkbcNGJAvxODGe98YyreCrDT4bbUGp841JA8ktJwJjoecTv1AnS7h8iffY6jYqW
EfB4Bca48cmjV82RtpnvxVlrD00c+NFtW8mgRhb7/U75aFywX8V7GdTrPPo3Ab59
IVVCK8Mn+vqNzI6yf8uvDRdQbQFG66xyzzDYFc+j4oiA+FGR6j7ch7B/Kul76MNP
BvtXIBmCVpavuFClxwnobNKazGp/LBUmHUXDRqlXNFlrnCmkkV2j1SJX8czN8GW+
kdKuFF78pMKD5moBau1OzUnMMyAEHwqbdjrTttTzko4oOlfMZ5BFeP6iwl+azfnX
DiOgYFW4nvo+u/beB1HzaSMPxWKzmo+lWWpopqrSGjKpad3dPMT3j5KPpm8dnpGN
VfRORK9ncpsLmfxh4zvKT4aIagiLArzAXb331Atngl6UKcBi9Vxww4qGhxusFUpK
2aKDzYUYbxEKLPSC4oWsTwPcO2ffJJieWtQf5n3ormTNLJgKTRiIO4c5y467VTLk
/+gL3AHN9+qvX0k8a8xpS78Gp+wWPEgcwuAvheMP/3/al+uqU1LVIKGvyAjQPaDR
gIk6yG69umbWbw5fpGSkxJy2EcdV+S/l35s1io9ga6R0ArG5oY3d3kvr0eNYswo6
hOORQ5luGlZSra1xLQoH4knh7IWKZiL0UlPCcuPgzTd97pfPL1zEHTZb8RwR6T39
nRPmSZ2+wXI2XuctexB4PrR2vTP6Yvn14Qn5MThm6WBNHLXAaJ57vJjGtWeIVv4i
HvqX3enarXfcyZrFGz4EgUuZ4viTBrOWNDgjFPSyzwgPK/SbIw0a9U7HoiJlcGD9
kzCcisLVlozdhFTv7A5pgNt04omC6QLF7IIZPTdhBMqRNdZYBQGVLWQLOZuJhCGk
z35StVe+skEHXxm2eko1cVLVKQDUmAUG/0jL5xujo+NPdoM3PK2/F5DbV6R67udX
cIi1MQ6R7EfrHgwvAld0Y1bMHcnZZtYwp3owZiTi28YR1E2n+xqtjzBo+tdD1Gb7
Oj/KUv8pTyAJ6bWzfdNWuTfA1GszSyQ8aUwxPj3jyizOiWrrgIGo0d3hmfx1AreF
Tq9/Lp+7Hy+6UVaimNEaCDxRcdU8fufrGF0Eupbp1x4KYQXZHFiA/2h/KoabXWYU
MgP2wQz++PVGwGWBC5aIADF7F8rLrjKfmB+jK+Ej/JGC6O7PVJ1IscovQ4GSXEes
mciOmEKYrMIBqUJ0r0Zm6HUHG/sdg2itc3rq9aIRoDxA5mztf/+chO89mAWO2FUn
ogQBL7PJYaJ+kHSjWQaomQjHssK1WVkvIfxrJiG8VcKMbaEpdUeg9Y1jhcaG7MM6
G6u76exFGgbxUcu7Da4naPPcMxvdr7tqPDBZPr4sESJ7Psj2u3hR5gWvgDlOVi8R
fl6xQ6SDDCojlKNeIh27BS0RAAWgrq87yyMkt3ViVlH/m6AfphBk7gI7MkUw0Zhe
1oqQT4rPzfax28oMKN7Mz6WOVV4ij5nz4YgBjRnhtmXq3FDgcmlZfHrMVhgC6EzW
B5d5tyC3Q11GljINjLjb15+7sijgRu4yVEuRi98hSQII4llmaIshqGXsZEKXxb47
NoLpXwkE+dybC2+IdNwwDN9SVULsMED9Nan0FaWbFTRuEXMP4nLX5K10fx2bDazG
t3XUhFifbkImMpBrUyZFYt5U3DjJqBbwaon0Q/YAzWuR8sqfDPqtWc+56N+gvwtS
dHBzLaecMX3bw2e9/hPsxe6IridvsTHKYOj0tmClYgESon9bcOiNuKgojVbrsF4/
n+ajhtAEqqTBDpkf5l6LyyIzSglGeLxxYwLA/cC5AI39fgNYVxtVaY8mNypl6+j2
Xz25F8ZeiRgnFsOvGp+6hIGW7uufkeC51BwAs2nQT1LJYU8tWLYXR1k2sgHQj6i2
OQeMwAMkBh4zM/spav+qgIAj1+V11RVKbHksAQ+hQxai8h2aY133KPFR0H85E3tA
cUpW1pSSs4Tige/PIhxiGp6ecCd9VIcQBKGhkFGtH6SVW5abZv6dQ+ZrDKnGKXYc
jDLS1fb0PCVJa/ArlnLlKrDlMxBUMw0iK1/8m9Z3O39BsTATobjmWWh1anqXUbDF
0QMvKf+uYMAeoIEv8UN2Gx44lfFFjVWFw+H+UrNRMaoU3pFkvQU0gD5ZaMx9Qw1R
UwBmXN9d3hBP418HQpHq3tqyUQ+CYdW8h7FNicafJESZXvEUrzqJZlTwdsJhIHaD
HatK6yrfbKQxYoEndV047/y9lSNjsQxvRlXI0Zh8zS0rd/VcR0VoSYr/yThTvzwp
mnq1eVZ3TT1ko2c7aslGIE1rO8TguV1pOO2RlYZpzXyphgGFFg1ykLo+5nL//leK
wdGU83HBktcW3jZbBD3Z8OtxXyZ+EUyVSW4rpCHN6uFcU+oyjb8qNSB7UBI0TH2u
SP49ZVyEuDyFiZ7lmKgzA+OZ/zP3QiFvKY5OS5sQ88lwB7WrjAUPsAMnlMTc92L9
x1JYmfhUWZdEFeO72t/LAc5vvi5AmuEJceSbATQNH4XC3G/HPZRPShbzenuj29OC
h/ZcAe0fQ7xe2bctKO5v7eRp5uOpYKBJSo1q5olv//GptfVCBklCY/usgj/cDZjM
9BAbBd0XJ+BmuL2D3aRyevytEe3PhpYbjJBf1bwTlM+pIFlyYT+UeSA1Z8RSzuaf
zJyK+zBOJX35IruF8fjgn/k0/YmXnaAsGd+p03tXn1n972K1XexdaFUjF1DqvSlz
QyDzUAb0wfv1+Oa21f741UlhVvoEmZta+HYvDIgy3iN7wKAJiswtB3QV1w8oq679
K06oZFafKah77WnWvXLAbsUBc8uIh5KA5f4F6n6+TMnV70nkrqxwDq0LVPHAXJbK
IYE3Fz71Pb+PJsBvc/c7KG1n6ySKhj1HgOdyxq95WUgfDcPzIxbTM4EMUE9rNSvS
OijTD+V/2kvSacamC8YFpS7PC7yycP3Xx64ejp59plc2fCV9HjpbcJc1r5Zvthik
XCsBYjFuNr3An6o9ZTUmIk83ngWtnZ+S3Z6jjmjK/4fj9LOjbtapq9DYlZwF+Y7J
Hns6Dr/VsxPMddDxgBS0wzwEHzney01M2Jl2tkzeGSyMNEgLWay6u6/ifUlyyXfB
SS580SoiAdJpsag4VVsoVyLzfhEPgOV8lcYa31eBD9Nw6Q4YfBhQOVv77ONDiVWL
/aOJvsNYFFLci8MO1LK7li5h7n8S+9e/Zj1okRYtHDP4zaJ7+2oqaWGUH+ypa+VE
n2lqunp4Joag3M8WTPUE0g4LBE/qmf+hVMQRGSxOM7iLXn1Mw4TKK4xcrg89Yd7z
WtwGhcLBG0bjSGp2+IZ2KzKVF4/IstnN9S6gwRaPB7OwD3MR2tUXARaYAnlcdexO
pQlNjmzgR7nnIRRnTWmK3//HzSQusu4iwX0V6SACh8CFIkmLgLudna01IZOQWiPc
EXl4PBfDtISdmVptAGxAYwg1LK6bdpmDN2/wqhR+bSIClBYNv2xQGefDXQp2XIA6
16yP4fo6Rk5h2Yp+fpBlwl462bQYQ0yCbEE9HRIT26sFI78UhLB0wWH+v67J7Oyn
C3nx8LbhFozZcgCE7++bazMCzLelcYN9pnr6qFcWBK9RNS+Pdc4KbRufceezu4jT
vzp8D2ORnfXmbr44Xn2/LizgLFtslz6QPwSa8ydDM7nD3CXDZH7E8jckwoaQ9kcF
wAfoyOBGiVjtAmjKXdZoD1xvbeDK4u14Cznlu7+Fvoop3MD7G51hXnXJaP3XY/hi
ANwfyZGJbgWP9JPTGOwY4M+kxTs1t4GmJ3azSbu/xVnaMWFjCuvRV1gF6mCF1+hH
iO2D68hzxbwPK6J6dbMmdue24/b3alhslbIQ7SSv/4d5qqrDWa1AWJ/A+/JaYuYB
+7EQlo2AO+RslqJJnRlCwRNhdDkX71u4cVUuwTRlTugKj/YJI8w6bosz6q2sHu70
hXAU5GtdfvzpHcFwTQKoQNgcbJoZ7i7hMpHGwisQHxrqWFfOmzzRFrY06F6JdWAX
TrioewXoSUgOkxRxFN+0XjOoJ9pYfLRqmn9d1sVp3B674C2HnKhKs6vXr5vN1mol
yvc13/diW7KehxC0hSjpguUxWzZOEHwad+d6GGp3uOF0rPLbVcHG0/z5m8Cg31I5
F/HjZB4xVZQ8TmIQ9xuUl1ErVOz+k6JC+Zm7w+JFrjnHDh2Gfdlfmq4Ks+1vBrJe
ImX9ukUsQSeKQjNLMHLXkhl1xfo1ANtKwGPuXfbBy645dLw5xFur4CTuyGxyf9ej
S3QIlqzCPhSJLtR159yXvGXgwNl4jcH/LjOmWhSmnq9jiqxWFof6huxCH3BJGeEr
F65g1+SqXWoA6xHQtXDCvAwd90ZPSeRIl84TWNFaNXROCMbfrdrs9Bi4gLD331y9
jau4vWwh2k9DrnNwh/2Bk7LF6039StzoywgkVv7Hx7qcO/4ElPpVyfeQPZeBkBRc
oB+NT88nuOEFfpl+4Tw20VhPnGqFhNlTU3TYR8qj8UFsvobUIcW9OR7FZ/ffKMKj
Xql8ycq3wA3CS4hY0wS/UxkoNJivU+qnaAlW9k9btzfbgW+aUEExZIJVKyMUkcA/
GXYGr234p1KxRz7HTuwvIp/JzPNPaxE7Fpoef5QdHSG4jKd52+u3nvYMcf3nG5SY
wqC/GM+iNEJy4tJlPkQTL4X8vbc0fgHPq1sl4uQdfCn5BEMUDtK//csxP1KUsw4I
JOH3+Y9waG73LiiG8XUMFqf7HiKstbthc6E7b2RL43dqu6YuGN9pzrPXkvNlaNOB
o0IxwMg+YdQi3IH10RNRvs+cymM84MNVKkKOxPwy8LGx+iRcZSAAKZJuPP8juyzc
7fps1Yrwz+b2u04wlGDUm5wpJYjg6eg6m/ZyQMf42IlP2kUhVOdex4b3tSMo1wdx
wAmnqS+8XClpD+uSWRJ1xRyUcqiALRau8T/9070Dtv3tBLZdK+2R7fun1z6gbAcp
/kdFiW3qbvj7VECe/2o8kIROUnvWNbAkhxt3yr0hB682CPnQ2dBGzWjcELPQiEkf
YRq+y+l0Rz7Et+Anl9GcC10x4YnzgVtja5Lf0cLEzjj9Rw5kQm+urn6SaZYej2n/
3u0rYQMAsz6KUURcAqlg2jNw3I6EmpcI4KTEbCEmp4zz9kFgmsDKnw1FxnT6FJYi
6cl83lzt70teB4Kf9pi3Hj8P6Gf9WnsmbfyFts1tx9zXEPTToQsAF9x6o9rOmnkw
7hGiiqWlFiVRQzDMn7fQE0wxZQ5z7UR46pmmUcsm73eZEa8oXwCwxpaXBq04xhXG
Siq5EnMr2GKkQ7Nw+OPrv9I5+Gu1odFg2XcmC8QjwqhI0yGbXEIi8rvET5HI8N5N
jG/aYkKnicUU5NycOmXFAA4qEXok8bwoFgpz4evqtq8M64sJ1JlX7jDeZNfBQW85
ob9jA+1OOe8Bb4UAAGDvnc0GU1IPAFn02Y0DCJD3wus+kwLwZdVSLOmOKoRSEeAz
OTfS92ItDWKiOlXJU9QPiMT/qvx9EI6sndVUa5hpWoP1GdQETtEjRDUk5fhSPZvO
mbsa7bOpYiQSPYEAaLr3IOyMj8AKizd/hRWBbLiR1d35+fknWtRFm2z9fAWIUYZy
EG3v/6zR2iDLODeRLQ3XY6RMaCwwuOestQnF8cWszWSDvYHhGug7zyWlZOtBSzWP
k/XKz0s/L6tsBXBI+zSfrvP0/qCFSfnKVY42cno8mOjGXEVu2BHLJ5REGsR0qSWL
Isrogn387EmHtyPgA5SoAbVf0VG3DZf/ig6bdJ8vGAVoNcmzYpffebShcymP6jxw
pyCpXL+9DR9ZfEN1tfmyYvgBcb2KcuuPLj8TQaBbjfFKLYIo0jOG9oq71uOPjop5
vKMvYdTcvAFmDxjC4qEk7CLVUYY+w2fvAPm3FlRxKuOn/yzShiq6EA4C1SGFQggo
Jb2M7xLSuyour2bIw4PRi/fF5EV4+Bt1sI3y/q2bK6IIm6wrgPfuoHGueIQQwN1r
7wGI4CoFAh3+IespRaLWMHjUsrjqffjY6zfwjC3zaDum2So7yK0E8fyODaI73nUE
CdmSkFU15LXKK8NwpXzr2Om4uBNwPks2fcS6o8s424SZJJ6DSBDzbGp7cumBpMWj
/Fnsy9SSsGYs5Ljz6Ht4AVXygplG2ggLdxBHAJSywHAEVvz+YXOiUOkCd83uQ58p
V1XTXlZV33yM5J8as4b3/nJvkBU9VCBST/+nXBxDb5n/cZyO+CS8xccTJJnaDc7b
kYz9CrlCvwFIos/JQQ9hqclfqeokFcF4emLDPQFvFBvEjSg2kW+ENJk15tY3sZXI
RT4StTiI+FvZZPkeBM0VE3L8BzaHCsSzhIFcfXlOpKOY2n5502slkWD4scUGh0Vc
k5MZ3eXnA1Qyk1z7qlKl+UcKTmxrS9W5GyKuIpOtaDUm+foMgJkle5qTX9A7ZN5g
NGAyXs+hIIC7ofeIpSgCte787uIX4whWn4PlOZ4UnHoTqtS0WA8ApU2E0iTp1pSq
F54X/EmoOmudqSSr/gEcvGS9Cx/22UHn5etvn7grVD3ZTmTnVoV0LHGE1/j5rBOc
z+/1BREQWNMUl+49PvqyCitKAm0ADWdT6hlma8bdMaEETpz1NTu8hUDz9RljqeaU
epYKyg/GU4G2GCxfntqu6ExVngIwGaQuawmstpqDi0STP1PKeWLRNgGdZmyAu/Yh
2DMWXCPY6CQb5Mi7m+OWCfI2RAxtoUpGlgN+63bgQkNopi2k9cfdT0H2SpFEP/zE
iSt4udCA20TYsMee2krHLRmxQ6ez91SMNNxCsb4F4ACmQsIFTmPjsP1LlOTcDfgY
xRHWNbkpWGVN2X3m4Nl9FV+uTZD7tyfSCFhpxS/YVGnGndvRhbi3EbPDsfrIBcxx
sGuzGJeaZnPc4c5CEke7Q8Z4fNDWU4oT20PjtCqN7gyWLp4UIZ3AtYhiOBMJ3l7U
+o9BFbE8SQqCsY1nh3YNuNJtyXax9Bpy6rDFdmBXHJAffTrlWbl59gPOW6OZSOIJ
lwQ6OHko4duICB7N8bp2AAjsGIZ0Yqf/XoW7hfwSJrx4x+BwilF6d3LhJxI7i3M4
ti0uES3UhIkaoO3GY0QR4rDYEsFfuch8+8SVxfkHJGnktARbbNVbx7bHCRuOKWYQ
TPxVqKKS3mLRX3nIEE1WL2RZoQnjzkSaeF21/Pz5x2UvGwcQ+m9WMBuEJ4NtorCJ
A82n1Ks5knS/aJ6XdJ0otqCESyA8sGGxZp6pJQRw+zscztJ1BnhzDRFMIVdU2egI
q7aFdNVkWt3mQ63tw1fTwVP66W2c33v2sNMmVuIO9l3y3mRcp2vgxNjdS4LrQLRK
OctD3qSKlEia03nU84Y2vQFohL5DT0OIIrSQ/CQC5qO8jAHFMYYlh9trFDThuDCj
2sbfPcRPgELS1AvQt65Z0UHtu543+Xhi3IG2V+NHL1ZkjWiMS03gtiTcsbAPN1wv
OpSfFl/49nm16NHqgZA9A55uT478Zoni6ZIbDBaLEgFzqhdOB91NMRZ95lHB8igE
nqhy7HRgrQgW+Px2QH5+XvLFXiWUnsIfVNOqZz/uoW34yjYlTuXcsM9Tag7od+Ox
DiCipHQ1AEbDfnL+hCM0bd54L9wj8xPjOyzlWtAmuZ9bQp4Y4C2d42+TP5xAg0jh
auCBmuRlhrs5Jc2zC14cYM+HJ9AU+RBdrx3qaQAVVuvI0asMNKPgs6dxADK1jjQB
Km3bn40gSlfVgjIyOWtLrJu7G1bpnVEf1TWE3Sm8lozRqfEY274QpC5g354buiuj
+nInnFNJQBq2l61uXp9919eaCo+Loaoou4X9BPygiXNNYRFcdQFDx7N5COP0SAmu
IPujrbCRtBznBzJBJTdwPxI5fwfzS8BUHZN1ATMxCrbxYPOG1IIR6+prjWBhD8du
59onV8GJVrdMD3JNtTXeJ1zxEu+y5Qo3UUTNOV9B9GHasPvuqnSifMqfMyrx34Ia
oY8GHbdT6iyTtBFMx9Xt1sWsku4w8MM6OC1mivUdqc6IvXrDmw466GWDEwLu8HWG
LZHaRkeHQ5qm1GxchqaP7RBhnM6DsBPWh162UJPccgSCxwPRlCK/O8vgQFFExVuf
ZQ4sLL4NqABf5BBfYUMtfzaOuSuMpdbiqfQPPuFUpnCzbLDVHy6w3IwfAgbE+YMb
whus6Xymy/ZoQfm1IH8HhKr0KuKDIqhMkgfwyemMM+sZR6uhg3Pn96sGrV+jjXVl
9p9ClP8/mdt66k7GAXtvmSPIO1mXPoM5TCxDWabDZpeAkOWwRFZxzhEmJ49Fa30n
W8AwRKMxxm8l8xduHFjyBlYFhWlXjs0CQjN2uPsQ6UB4efXTX+8VY6yJ6OdMq0NP
KfcNZM2UPfYMa8v2nNkDJfLbhMJf7lxqjSTAUeJ87GyhuerrjRPQh8NGcLGJSK9b
dQqp/Qkoq6tmR8tPVQ1xxNNtwRi1WKNNFBNmxa6we0a6W61e1zjDiNPOm+gGWsBR
99aYCuetc3n7oM8Ms9ZwN9lJ5jXrzGkTVkpxK/lZ79kfdIToBXt7USXJhc30XnLr
+AgNr880iJNKgVZVtFFqLoLIOdODoMj130vlYiAWkIbHxkJ8zUxY+rsqoPWOkBxm
hR8DNXwvDip5OciJneSbVjKU/7bsVr0u+QCLRQtf1CzDpGe49N+B3fVGfEUgIuXo
YChZetNiSdLRcM75aobFtF+ncOpHUO/uNJxtae0U2oBtY43e4Ze0UFuqzw75vhKH
oWpxzLTGP8PidHRS9PnlGgM5WggjBCEJHZiRI5PlNaxMAWjEkwLXNArAhfB+oGa/
GT3gch1vt9Bgmv8pa54sCxt0B1wHvvl242He7CXFBp8fmCBuepLWaH1QezP3t/eu
lu7FD2Ud5nmesfOzswFIwveyKxW8Yi9cjgxVgazlDkCUC27L6CnAVqqpNkyo071c
NFohXLFPuzvXHU54W8vbDQjLd8/PXg/0/aJCPWkYuUe4nlS7df9TxrzoirvMBL97
kQoWIlPnJFlYEB91bLksLwtSrQ62/w+6Q+En2BCkmWBcO9a1UiTbCexVV9MRpImb
rZRucooGr011JjICM0LGjcblZHItQVgVBC0ul23OaGiFFRnfSeSm9VbYt1cTnJK1
F5kl34PHGCEaluV2peq8nCxvGGeGftIC9/lILDWPRcCvZ03cBL6BO3rTvF6n4Icn
xnz8UNZ0NmsxJeNnibgbuoXzGNoau81pTtePUSLrpFVzcaWfg5EEUgP/kAlt+3XR
gwn1Rkbl89nUgfMMvTcpKNng+Rieesluc2XIY/PD8VQQLdm/x+DyLcqtcdWW6l1k
fUJkILWA3xXOf1Wy34R1o09F0kUNQii6tnTFkSW8HGBikjKY08cyYd/eiTkZ3vEY
o+iDcokUNNuOFOqiPZyI3lMDYFAm/NPej1iljU/8bXVdRhN+blkc2YDjoPjflhWg
XIKkDXAPdSn8PATO12mXE5EE2OyYFHkTBQpSVF4ms8pRTB25t2A3yh25iUHCRhhd
FuvYnSA7t8nzUJmWJhawaL9D5+nUsd+rIHt5jxZuw9UcgKhe+RhdPwvh+Wk/WWA8
vCzaogyJ28Pov/k67m6q9BK+AizmiY3eUMwDCPyZlt9mw8bZEIV9iOY5PlBZ0ESZ
f9MdAXG0j0pU/lMVewJaCELzchwkaJHQveAlpfON13xx/dXHk7t7xQRSqSofE6WV
un46v7qiPmuoz5mmHehouE9qCPczRkN5lz4H4kqg2l0WTNmw8TLX0R8DRWEWu2Wu
I0caL7sbN/aEEGQrtoXK+F4u1fmaNNyjhfexvo+mJQZmuwVOWKeRUTurhRp5PeBR
0YvSoWAFL0EXRgXiN11IyzhxtUbBxmdFuE8yVY4FgqriUb3XeLmkBqloagAfcfUH
FEoUmy/HhbBhk2QY1Hn+pkNy2dV8LzVBp0bfmc+TEya4O9SQVT+FZJ3M+3eKaNjn
gWCcpY3lvIZd7TV3LjRluZFYfNP1GO0isKHeMKL067NdC3ix86vYyzIBfqnMCswu
DUqEKCwUvECTfdfJQ9gP8Np2irtqrfbUP10b0IzyD2v96qOHWJGAoVG0KQPNKX++
8cVGSBgkxp69tpGl3R6y/vgMusOCliQqjJ0Y5ftNqxo8J1DdexgCshfoSWZcR0Sh
wPBgAjkFGCD8MVlODIEdx03P/VNyDK+u4UwM1+gOVEeq0GrdMK/Cfo366JDo5ryk
WeQguMk7Zc4zlq82Cbz7nVR1EwrGlFaVs0Vgje6d0lWlGMZcNAQcJHzwHvx74jwH
ktFMt6dXv+WlJwg83IMSf1tHCZWT5dndPmdazvIQg8rs6paQq1ImWmfHs45v6GI8
qVS1JIIHCMD0ki3bVkxhxNXd/rXOXn9rif2ao6OyS8P42NmK0uKJfDFxzlVdebfh
kGs/DXwaAX3oFgEPRO3ODLRT3jQDa4UcVm142ho/Fr652wd+jjF/i7TgwhyHCodl
7OV2JF9CQIofGx6fWfrSfVvRcp2wWdnFpvVazwtAWqEZkizTy5ZCKQqmikKdLgXb
stWkFLJUuD6XGrrUpVS0TntvaTI1FfHmVp0YoiXl4Jw6aOsKAPjLjd8Q/d8Oiwcz
mIr80O1xe4DTJjrkjgKPlRXG2OScWVPOPNU5QHbtwUN7b8ado+RAVlPGoCDc6fxM
dl1EH65+u+655jjP2gLzyIW2LutS0mw7DcOKSMqb6AcjeNQPS3WOgOsmxfyNYJgW
Vm8ygXzGXHlHDzDNN+lQiZUZkaCIp6rAVehddcnnn1lpjlPM57jkUNd+C4NdpClB
I89YBym9mi/VDt1yXUfLgBxzeVkrxwtJlS87Pn7MI5ocDD6KVuKMLjywIZVRabaT
AottI9r6gKcNeqRtkmHr85ht5AIZEhAKhK+BdqkOTMcly3+KbgCsYwRQXe6tWss0
v2ArmjF10oYUZ9PUwQLCZc8cvCloyWImum15dKO70DsWddERsic4qXJbjg11Id2w
rlfPE3MY8iANX6upJpdGNaV8EjjS9bJrJl/2LvNEYqSb989v58XtekOz6xr61EJR
cJ2LC1JhYAhyFIGR3xFzHiwznxdgk0ZHoOwqr/WlLiy7nzoD+zrDzDCTANj68yXK
K2OwApoouNvA6I1D4ZPqHFd4HHgDQNeo/zbpccQfO/fj7mbk6Rm2wtduax2aJVxA
2LWTXZecAdDa6DFpLeGkk6ZXjecg0XQ2ob/8tyYVJsQ4ym41eSbHLhIB4mnGGP9l
SWFFOKWZMaHz7IHbjVVtclugee+QgN3x/Uk3qAgD2+i98WOyL2zsv0nz0EaJA+I/
8AFjAwnmTo84q3Jt3qVq/2tJbDEcofaj5JpsgBW1ymSW4voquXNUdr4xf5av2n+6
H1sylbt1yUzUY0kRnMBComIabc3kI09JNlyHR27p6DXoaiGtlwRXgQBmM6kKZyOJ
LQl9HivzEjS+Zy3OL8FB7A5FkhFRl1yLKCa3DVTjph/BEC6i8fHvGkLwEx0JpL2y
Rf87Fly4tZOb0PpvW3pTaNH+hqALSV7IXr5MIWBNVQes5cNPzIUOiczA9QZ/dD7t
Rs+WVbWoLxR45vE9TEZHYuUnVDuVtMPLVJTOHHx01CD/zpQYyq8Zc7pxzQCLiC9V
GS4b2zWHLp05tz2Lx9bZtyd0dxtbW5OLlQN6kqYt7PIh5LkZaqVDC93AwSfK3R9t
lhyxEy5NcbbGC4wJMwCCYRw2zC6SM+SBXHzIpAS/K7vikC7EPajCGx1a1VPLRbzn
2KSCEaY6vO5yOV+9aM+uWzTjL5WAqQnq9GE3GI60oo91OimIyFl1WVSmg6nAyNBR
q/fJKGhsNuQoPkRLm8c76n0w/ZTh/9URh1a2jgVLOFlPSW5lPh3xrVCskLmbgvae
3QVsvtCR+e5g15NQaClEzLi+Ve/bp6Q389sFKFAYyccvosfhttlYc0IRWRNi7+v6
oCx4MgvUDSkGh4qlZ0xodYNmEQlY6RK1tzUSNDv37S9VhE3Ho9K0rDJl69vy71Jn
PmXRu4lHAhuRXvQ1ueKEqMK93yxfIFZPW17JD16wcChAfKog1VqAZ5R/qtje49hZ
0FuYJO6Hf9IZgcUhlaII0ehEAd8w6adapuoFKoCN8QxJIAUVnyEBNLmRPc+p7t5K
HXJQz53/UwyA5qOJh5+9CIUBZQXV0scniaXgc1NBp4JaW3pq70YhRs+t8nRuSDc6
9cGX5fR7iSs9ERMRW/3m+JLlBhSvA7+vssiJJ5Vb549u0em5IhrGwtw5o+ezZvdH
ZwM3S/B8rSi7WY1FNhuOhW3LSkzUBVIQS3tJd0nLyYJGOVpEsgIjIPx7eQHn9llu
8Sm2VJUzSN/58wUYM7HNNcQ0Z+yBBlYPym/8kRt02iYhCPOjTqWLRbyhgGg+uWQr
JQ0uNF6GKIfULKSGPN/410fuz9opcwSW/1MQg1TyLnAylgA91RTKoA3TYO95eXSJ
Rn/IvKoqkftOd/6wnnt6Or5PBdSeuCOep7wgIEkAitfQSB+r/A2YUuTf7Hx33vCG
7juhJA6FmLbxDJBu0itd9PZqC65uHH1TV1b2w7iRBsq48tAk0VoLIk4T+nLQ4cDp
5zYQg8zd1h8h3FGuRbaDlzBFHlFfytUxY3DH/KH1Y8winnydP4JQecI3g5TqrUJ5
qMgSnkpxsi4/DS9lGQ1Gup9UZ0yh8bfIwcorJ0t1HvJJ4TdQCxLIbpAfI97iKp3b
f/aJvVc1KR1dowClcv3aYjjX/oVa7czCRfUcr9MoJNGyZspDDC6hjDQwldsCEJC2
4goNtOXZAy3dOfgqhSo/SxPb+vkPqYbntCHUAqAbohGHXlnOq7hoKJQekBvZ8WjP
dKvQ924yOk6IQwupvjPqIDLLQOuViNwFhAX9QCz9g5rlbpGkep6An6PuHclrpYUl
UFDgiRYg6fH9Xeq/D2u1NY0p33+8ck0LJJdRgU+4d67J5YjCVzT0FWarL91eodSm
hT9TUz8+L2JsOAI/zv8WFmCDSDp9Rtq28g+iAprUG7Jj6ZPkLg9PYa6guxd69gtn
06x2h/cSGLaKAzw1GuGCxUVkfNf0SDkj2nHN9lDPxr6m+7+LUUaiyw/JCQPDpZog
zrifPTFRBH96hwESzkaj3gutz/8uVac0oE4rxeRErEu+BA0z/dCIKIYLAj+4GHXv
e/Fx3GwpFJEjbAy/hv7icpbPn/vT2bkoxsLtWnKtOk1WaPwaASahh2yaVLfelllb
yDwV/K/Z+3FqpuI3aRKOisOI77mH+2nA5zp1TQO87GyKQI3gN0fhtE+7Zhp7CL0x
pX8CtQlIWBoNWOZgkVBUxy9Z5kydTx6dydch6x7X0qgpHlXEszw9K6u8BA+mFHzD
9N0aBdlgNITeRgP7we9S0ajKupxgJfT6eut/yrqC7YycLn+b8fAkdEBRwrpag4d/
prBJi2MsLSTyhJv0fHmXldaQP3qgsnbnjlEtLM1PBMHo7p9CE54jyG3iZ6IF1VUD
`pragma protect end_protected
