alt_sv_issp_gbtBank2_inst : alt_sv_issp_gbtBank2 PORT MAP (
		probe	 => probe_sig,
		source_clk	 => source_clk_sig,
		source_ena	 => source_ena_sig,
		source	 => source_sig
	);
