// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nc29QoQiJxGYyK1/DKh/TMoWekj9u5PMo6QSM/8atOalvIK6dhfEZsebixlUXKnA
fIjcrpb93XTyHipH/X1L2UmwDqTbGX6rYYM2YQB0dqxPDNnB6/k8fCKvwR1wkTt/
wO6xNkW7M6Hr8D1pZYnymTSn7JZztJFSC058a09cEEA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8816)
Lshiz8CL9wS58DH977zaUeDnxjMNePCKEJWUDcIdQrSXI8FooXpJC8QQcV1ldpmP
JHDza6i+dW5JM6lwYetkjTOr5r63W9B+p/SpTrmwWveockwHiOY9jxQtRbf+qqOM
oS8naE8ylHdVODrMFjbf8AIdfA+ii29FEMWTwxhZ+jw1NitlNGxZpLLV86Y1Uq/6
6dodaMRkz2Er9wMu8tUHuogf9s+QzGi5U9vnknr2a4sQUkCE9qrKL4clL9Yjcl5+
5Ac98siJrzZReDrg4AQayoyiW5oDU0lsNdyJAA71SsfjBfjRm3DAxv/12JSF2q2J
bPpezxbskgqq5ArQabWeb0BM9fJJlX6PtAmlniFMPWOdX2xMdf6jtks0W7/1FqlK
lNJygALQAf9mp+4s/DYOeFI9988g4TOyUbhuAD6bEnV9WN+BO6BIdoT9Fatu5tyc
xJePqJVDjgPJrT1iUvORJx78be2jdK8Z1mTsYKoGCOkekgKxVyyQVuq4E2ly+wtB
T3bEtbwrLDG6qGj/hjf0zAroEA9xhYXUFZLdAUJVFd6/2dg8zHVc9/TbEv0mLdP+
R6YOubPmtdLWpOQQjRf+GVA9ongPGD3miSAprGof6YcoO64QJEMykjA7N6AS71Uc
EOA9IIYKzp73qJCpXpAOQptey5YK0gPW2A4G9ONyZ//TM0QF/Iruah0Jy0s/ERDv
BP3ArSP+8plJlFG7Bhqi9BAVNrQ5eORVZohIyR96CW1r7rQIvXHdBx1VnXC+YSO4
NAZdYC8ZaBH62cmmSBNmIPNlSCobKcvkARHxiyIn7tyMrco8jsup7obWsUAaib30
ilbQqCcjCzlxLxU13pIwtoAHKofQjGbfLnaSeVh42DLo1icVtCVvnQKAIBot4Ys2
9l9i0l9nShyJ3QPEYOk+JS3/0rFrxLFTDIHufR+f0U4WYcMUytyd5E642xZXDv7q
oUGBWUvrC6ftXrZeCO7MvL7AKji9ZVZ4U/y5ZwDdF9IzCkqf+JW+bUlWRKXgbJ8P
2hx9blXVGyotmrbl6fZCAF5pRT4VAqLDTG0+43XWdh8DeGX4dBr5bFJMnNDXX+vu
FU5HH1j6HkWAOi1XIXbUq/UkWPKllCi7jrfirx/zLJIY/IPKdHue4Mj/YVtL/+Tz
Xdkdbmn3O7+Jk3cDCCDK/162chx9bl6Ztj2KOGrJ3Od4OxqnPEp0A/HI7lnsB8ci
0f19RZFc9T84skvgZ/4Nkl4Pd14FdmG6cl7F6weaZpDtCdxJrf+G+YmU1u9Vi5xE
ph/WOdRjJZrGowoGUoqJooll926Pf53dn8ZkLpnYf/ksq+J7wJeEGHgKlOF6Ra5h
+2qkSW/+xWFwTXnfjA1NyrlCPLdMo7kWG+W/LedHbZl9HoZI52rbEaDCvTqdVXcp
qxPYdb78VqcuugZ1YGSXVAX4oXRMspfJhQKBL7+FSIjmpYRwXw9avST6SH5Xw7SR
+aSDYiICXRTWz0LM7xtaPWxbVPzwmuy95+xGDF9MdYjnFyhoRGD1+vYgXM8BkJHC
R3F+Im+RaDPnrR9i8kADIA/9vpQbvuq6yLtccNrDZ9WDXQ+9erLC/dVviBpap84u
XFiNwa5LrHuI2eMzP6iQbghEeM6oYGIdbJ6UIJYb69n+CkGHcQDc+kPqNZ+kueVP
JK8HGCQL6Q+TvK1qgYAd2sZDxqLWfuK8F/gXod7SltHD+Yv867r356Mg69Po12lt
BV7c6qJ52cC4XTnikdmw5iDgGL8Mq8uI+Fzrkw8TqchkqRZvLAnKlOiOJS28msaz
SIZXpm6xu2fY6KP5Qie7VZ0Ntq9ALxuJ/GsA/murt2Tkm+vWhG3KbxcmU4YEljMX
Pw0uw3QJpv4sOtP2GFs4+DJa/J+JAoQVqZ2tJnD3HMlwB2GyWvDijc8FyXvj5pmA
sV2AkCI9D7fUbHdQqXIup7ouz2jhtNRI2ykekPBSM/aH9HO7MdYPBsw7dqY/Xzf8
KUhSencF3oIQ8jruY2rqMndf+E7vYK6Rd7/LCTzeW3WI7SmWAjYod2E8U34ALdrZ
eX8ex7/PYK5fhFZhDt127KhN4c4t93MoNL6Umne5WVwABIkUPws6s5jJ+GxhLHiv
p93QkNmyXThYtFuD0avBZFXzY4ZHDrfdhyCrpE4qMnNXUgjIG1YUt/p6GhzNslKL
7TRG1bVDqxYjeVWHkW7inNqITZ0f4XeVqrP0jcQRV5uH8cqgyrUxgsXzZcuImVOe
rW4KVk1yXeGX7WdvoHZJaJI1aWON099NW/RMLclMwEYypEbFCf8kRNN+Gc83p5Mw
RRI51sHMwdOyPGBu0MPss1qNqqaDXSYFD8jSIig6nayuCK3zUZluWB43O1IBAsN9
01orA/I2RbORUYzmkF1DgimEXa7g/rc0e5fJBphjPa6Xhd8jG6TBHGEDPxlQg79B
k9eGK8xT78UcaR/PirJjJ0dRywJr6b56PfR59NhlivCJ9DH7TRT2YgfDetRr7e7W
PZw+/GKdbsM4MVvUsXXaFNLmtgvmI+Zzeefkva3eZRge3lWL/sFd5jITwuNrDXqB
zhzGwxtbie/B4QNX6cw7ccjvhCv9+7Jv3awgfiYFq57MS2lZQetBs18i3o9jR0r4
QbAZZHPKpL7MMGt4mMtorDe5m2Q+fqaYaeXBxua/q4/4CpRBcLNGTFa2Za32wUie
uLyqr7ZHJJXztiW2g39sYiGtLF2lD7uOkHw9aAnrJWv0iAKvUfMU5lybLSbcCQmI
LuzqeRXI/a5LALVQm74KKFyz011A50RKI06LmeiGBYvXc2BkH3RLBspPzQZEjt0V
Bd04VEMsU819hICKtsiKay3GZH1S4yp5IoBw8oAaclU60OrQg384yTAkSmvVkadu
Z5d5FiM7jPIbbYGqCvWBEylDXaIMGGlQVMtuBIsU5TrxK6iti/9fDJTxHqs5Fckd
lsu4H4Nh3/HYMNEGCV0QhHHMOUEHoBd7QScfbQ9QuP/zns614AWdjphFf2CezXeY
CVGae3f6AxEg3zs4cOvAv6IfCYc+PaBwBcsQrfKWdXRFgoSDhqnzCveLntElsBJV
+BFBL12TuAniUAxyx4yYuqiu63c6jpA87DAj1M0hbCE1biLpLaeLpqgBZFQ5YjPP
ZFFXrsdOsNChY+uNTwQFjRc3VJFJAz0m5umgd3FQtPCQwib9+XTAaWzs0GpZ/47N
jrpWUnzIWddJtIaWspFNKHXdaGHGEOKPVLPkrhs7jsmfqkPCGrHZRZ4q2FWKe81n
xqaB1zQC/4ZEHCAc36xlEHt0aGisaQW+2oo3zGtkZ8zpXoHDsAmnJRfIq/pfhcu5
+B/ZDkozFCyL42mmvrvwQv0dp1cGlxZ2qSfT1koa7I1e/Qh+yLC8iAbxFBRhECdL
rafey7qSti08J3ddc7hFnqggn1R2JOLgjdCjeu3T1/WIKyghkIo+q1J0BEP8Sf/n
vBo7txyjujjPNghNOHmue7Xfx+qIAZT3BBUNeKDbjuugcHSWu2dwyzT3Wk7wOFAQ
66S0HEo1H1+oya2J1Mxazl44HeXYL2qdg55+Ya2e6MhJcqIkoY0+WZPyoAeTXf/v
12TBt3XOzUuCyFYJ1TSkfHwNzBjAbMRnY7ovgCxfFRKOATTCP8NveHf3Wt3E9rgU
hjX7tuyAD3x234SBaru3OpfOQ8iYRBMo2pN1LM+on4XGISVSBpiQYszqx8SZjef8
v8y41BgieZB6OHOpRlQkFjX3tg3LFA2Ocp+VX852kpeLOxB6V7dv3+kQdjR9BSW9
xFUp3UX+0Ubo2JWuNImG2vMTEMcY740I9wAra2hImFAlQgTO603zvpp30+VLFmMi
mV4PoEpxxmeVZKb1745KoEKCDv/p+mCpXduwo20pEintgkPmDTG8dSMdidNTT/Gg
XMHzo1kXm/0i/N+SHxTCuoTeYF5qeOQjxNRD1iE8oaBSi8iUZlN01C2bmkYmj6ej
L9pBxbfobrIK9qA4mIvhtd9YOjgXPDq0jWpSKyAIkTvtb8Tv3B5OI2I1HPXYCyRM
z5UzUugjpIYcPd/0BuaVKwncwtkllfy0tZ3K8t+dIpyVIlpc6vu2BeHjXiI7ZIJ3
NAn6N7eV9XFDderhWVZcszsX7cxQjkepgt3vyK/UvikluyRkEE5moffeuoiWAjHD
QTB9L/6lW278i1YizEl/CI2t7IdmPxOp66poY25tWP/ezx8KcQHJWCKQj3XK4zpP
SpczhBokOTJnmwHUtg7qkBZrzWicufP0YVUTIlrMrha+usYzLupsHrLBVOmAyAUi
YCbJOQ2GZAHqokszuIpnh5HsvDlJbe4eHnTQ2m3nN//21ySCy1Km0yWZ9NWHaGLA
LxuA3a3YjoGdwSNmz/A0/D9stuR4TCQfwliPUwP62rl60ecnNGh6CwSicSHG1DHn
EB2BbrmkBU8Uf/GhAJWN2tgpFxhUKZR/qchNy0/ve+WSjt+YlHSwaH8SYN5fat3d
E0TUJMg9GQYgSAOB1UwjJc37v5TDETy2ZMJAuBrf02QR1AtkKncdTUqeGkgJfb/v
LYS9lprpELWafH3lB3wZlYVL/JaCmOLxnswcrrZJijF0AFhlTe5G2aXDhWsgKH2V
xuPhvNsppklvlbVSAqDLc86kfQrVQdChN2OW7ZDHtjl8YT1dXkE8lnypfsX++g0A
Km3Y0jLEQvRVZgalvCxTe5OUtL9Jv1bcUHPUeRD5AqiccC1KrIBmafRoUyMNGm4T
p2oeOQp0oquCd9R8D5Sh3t29vH0pQAQIupwjfnIVEFpuni1xo3tjW0S7K5HeSngn
t61U2STbvcuLdWsakz/5eDAQJyoNR9xnCDDl1RsuhwKoi7xmmtb2FPP2Mf+tNo0a
JxPZsKkteirZtFYxC8b/gMnGJ66suhfnm3DXe+V34FDxXxUHivklMZcUEImkScB4
wNr0VXh2709hmZoXkql4jLFN1Kg0Q2g7XCVchA6QZu7opeC1/9vvVveYNzQ5eL1Q
cPmo2RZzgMHpgDRE2yE1A9CZBjMqOfQjLPWUL0IW/1N/WKr/lF4DlWv2HWi46iBd
xRUBj4SGbpb4vqNQEb4WholkN6C0GITrxgtywG5bPMKDnMclHHSTmJ7B098b+G4N
KUY+Qa8fJBRnyTYp63aVFlMUiPHmPGUTb5gfYOY6cAOR8efgUSsa7dv7Pp7HQo6S
pOsuMuwGUokS6iKiQ76A8TYAqT8KT/VwlfD22KKqvaMDWrWv06ORWdP5u+sf+JYZ
LwCBkI0HYrUEmcUGG1jFf4iaJJFQLtlM7L/EbQ2oefoFHkTkEz3t3muceYejSolf
07qnU3RvRE59LoJAfyuIuWH/99p0qOPV3mXiDmeD3+6sX0rkUynGqz/SWQM1Epx5
Y1LhYfK82FzlMsND9NYUt3LAh9VuDrvHdadrV3j6P7sM/i4vmsAv2BNhDXqeh5pV
+4VOXQUSC++2lIPh/hl2ee9rq3GLq83sytSyBU2uCNgpHlNrCiMaMOzhJIppmpE3
zOyHxrMrW7IwN8aQeavLGLvLmUnwEJHuzJZ6iWs5ZY0IruPmlh+aT4RZr9bSyBtG
x1beshlvKtL5f5cqV9DDQKSsr820wJdYbp3kqPGSbbREa5C7tx2aKi0WeVPilKtW
RcIdECVUZxUtsEV6eqgh7OOjCVkRd9YrYh+5uifrI4a5jcdfZYvJ/+F2z5To7oHc
LmmSHghjNUIWzKR7K1ypvGQKkuUik0S/tFV8O2IM4USLccvmnaC8UdElrs6P/qsS
ovOI1d4jRZ/cSLt0vlUA5tr1Oq46HbDgld0gGLeJ4fAqmuXMSOOdeZZt7M0/oYuk
nMfwhgUgadfDegdyW/4p4TAzEiJxc/0gQSBESxfckBTJlJ7nYR/orHQcZ8tHkoIw
Ptja9LvLbSXaeax1bs4iNrf2fzxpdVqNLwc3v19HG/arvQEn8nXbJYbDti9bD7qc
cHM/bQ8bMmNjZKy+Qn72T1IZPUdlt+Sm+OWkpLyyi4LewhXbSW30mz5EVkNA/kHL
Sf0E33BZL3TIQJpwKZNp1l41DaVyiu8cuZekz8UnOVrEqWHWNRQaadZsbfoA+kuF
maf10hdcbi7BWARltzby22ICQgbUx5DL3NC+rPBwQRXdOx6wYjlF2V/cjWAC7v5o
E6c1BVru7BxmNAwNOzoGGDuf7O43sxbS5W0DwLLAY9vihCE/HpwrhhZfSEZIvoqU
rwoarrNdeirRmtPs5F2V+VZOZyLChDM5jsNE3UH0xtPYuM9igTwYXKD6tTRnEEVX
lV1eyWuATTUe3hueXqBmPtE96I2Vw3GKrObuB4XceurojiN9aU4OnOEmK961gTJ8
PHerSwleUmdzi4HJza7Rq7MWkbxN9iKeOsdVwaGkIuCW5q1fKA5vFYNMAujzyrk1
jcUfc67X2swGo6gP+DvSg9CEve2oUGP2nrQ6qxCwwQ3MO5xk9Z0wpZ0pUi5Z00Hr
rGCNP72Nh69TbVGj/gSr82xSRHqAlllzO4f4nD8pVIKQbVfzsa5PIf6QGHCiGr0d
chGPXb/17SnI2re4FX8b0mU7YH6v2STbYsjgjo48D2s6bjnOv5whX+3bVpsP92go
uwb0rJKTGTrCiO1rC17WMO/t4forBZVVLan6KcsPL/wvY8vCI4X7hjiJ1BPwmjBA
SCDEVdFPD1j1HmnKAx70L26x7QBYq+52/OAGwCmqxQ2GjANCXmzFGXY//cFytS+i
JpJsX/5dwC8lDQwveFQdD9ocr/Yq7YsNmQZpPgaWAViLnoJte3Eg7hccMlKTqo6a
ZNqMB591iUQBPm4lOlEBGSK+i01HGvc3pfmOLa4xi3BR69Q6mNMVfQFjn8D8wxxc
peA6puCdgCMj+YAQH/GoqYAaZCmuv2ubONsaphQlN0lJYe+07hkCLmgUm9iTQJvg
QaJkYDyTHZJPJH/Bs50mitJMNdQb97QIP0M0yRuYVL7zfFOJdYll7es6RIl4yfOh
XJrFUX75Erm0sZfGXKiRw9ppWCgJlXVjw7ucBAnFljMn2H0ZdlWEKT5Zb1ublTWX
UiQIf77gKRUkuV7oMqZjFGSgk6M5K21JWu1SCq42oARLqVRSIP7s6vzceDIW6XV0
a1Pd4ZBKBWcoU5Ubum8VyFpD09cZt6iJuiUXgYTkAPFaOyJbB9PD3TRmSu07IMP8
LgCtpQCLS6EFtJCRyFSjCKd8Bjmp38yfszJvI6uaI5I5ruoTqGzy3NeVZcDfVIoC
miqFzkxVTrUNJqr06xZIazESMaIeXlcEqp4I5V7BuskWFSa50e8Hm+TfaEi+HwJO
yu8tbQADukQr6Ff40bLVMOZYCWQHzf6ILb0jKhiK9pimfsuy4dyFFWg7rD6wohw2
Dpx+wKYjry9BkHsO5pNrwpE6x85qyKIQoO1CHGxb9AwRnqbqIVJY5OH/HNBXQjc9
i1gqgsfyzMY3kVNnvMtJ0ZrvHchUgiVAiKJYoVQ1fhihFjHKkRAbaUFpb0DUIM/x
1+EYfbYWK62Cvi2h9plfGqiItCeo4ynhMtXay8q4Um1hpvXWvS7oFEVDV8p723Rs
o3tix5ZGUl8/itYP9J7+BhkmOJVK/h3KsKMUdrvc8lZliKA/zPIfmwUBuY5XXqvc
Jog74hjKHlEYWwbXlOSFsrUTvQ/p8sHxkyRvtXG51cZBfsHTf3OBB0p6kB37BiUU
BpHvdBMYyU+XwvIDzO1SvW1ckZXiIYZ7fXYmB6D7Eux4ZK/gt4gw7BaWsrKpUoxC
sTmly49BmNyOAR0Y2D3NHDH8U4HLKJb/1rBUSTehW/BbRUCtU01E4tA1n8BQCwXu
sbqecGVb/zTBG53GBURi6GV0dksREcvgjsJqhYExyZKy7GZnz7zrXW/rqcO+ULnv
C+yCjeMrlIyhveePAOXFJiHq+d/icAJBq3MW2Rg8G+uJgaOLn0ORO2GmUGeMGtKx
qXi+tHCqXtcNDXmQwOGV9UaSdhhc5yY/MRVu3DAo2lVADm69YHEqq1zmMnZHq8Fr
B9zyLkJWcdvZYREbaup+GG3CP1gUbuYWCwHdOnNTnbp0Ov/LzpSklvWVY7j80fRm
VnSTQEZ1V6SPz5kBReGLIh3dgvKdNK+wVPbnSgqJLHEc/kQAw6TgzxX3MjFQUTYX
2+UBCepzG5EitVVHun/OZiTfu8Rsnc8gatBrFs6gWWLrBwPvoaph1dgIZ3aNIhE9
+Gq1zPhojBfREs2HwR9ML5Fdg4psC6WhLnfRuLrQcnHmouwr1dgVM3CA0AhEaaWJ
cCvRyvdZkMcyjlj8jRyynbyfDTp5Xgu1xes+tpdK3TfcGkj8mQlzHvWPjVRbdtzD
kaLunayRwRNHg9Ik3g8u/1va84gPq3rCDAAEdcXC5PpBbdRrFDEJCOJZdd6ks0dP
OP4O8TZ8g8m27erYZQHlXw9AWvlj04olvJVSsTsX4a6+O/bmjufCc4ffaxpSCiK4
yj5OqPNdfd6MVe6PTK3YgNNtIXqsDxMwDed7jXm7GbEyJGwtfGij4zG+6df4NxKm
ZgmeUAROKe0iYjAA61fyZuMG9rAqg1yI/deOlBEaErnWo4ok7WREidXPgzzZ5uJJ
zK+NAcw7Rg0GyVo8os7f9yjPbQG38IjIixIcQmL3Q/1RDn/ctV7E5w29DqChS+9J
zdIPuy7pjmQ9CDWOjXiOkVcQKbUKH4PniQCYPRO85TXdkqsBXg6889Bu7LgrAo0P
I5mEXnBQcXQZNTRk1SnMR9CDVcEArESaZLb8Ehj0tj1iURGzvBJ9b/e7hTWLW4EL
hJbPyFMkYermSSU6lCR6VNVykJoCK0uMvoNHedYdHv3Tlbr8LHyjByyh5ve0EOq/
3QE4ScHd+7KkNGZtucn+CAa4kHVUdsmP8QDDnSbP6gVq8fny1QClSNC2F46S7u9I
G2ThrQjnanZZ2c13u5KjDvAEN274GNPoN/suCIXUTOQUAyEiQxvMCMCXuUdMkjRX
DV2svC4ZB4Whna8hARDzPZFJFI57BICwQBISjs6Bu+gBAK4aSaw3S2YIRSbtlCGG
07wblcFiUk5Q15AFjZxdqqjYCS6sV6FNAAjOOHMY2J8BBof1FYkQYTK6h6EoGwuP
szM/jZRALEzbiOlFzlTRtz04YbpyH8JJrkqxsVDWbrSWyiSIl4cryaISwqKX6xgD
nsnRE5jEIBsT2spKdVNA1wz3za+drSH7zDoFmgAXEws8e97tOWRX954Ld4iiJn9L
deYLwd+FVA4wly4gabZcpvpFLmhgbe4tcz66YgeXtVoKsGL0l3IoluDxb+0M25ff
KXclUkVHRP8vB/ppo+JNONnRdy95Y3znPzl5myNaVO3Nk+tSMo3aNQGaXu3HVIHe
auABl9dvXGJEdAMHLjG2NUE29YRWlk/W5okqhdRBTfDJoM1czIz3mbVsiYFCZAPK
E+XnetHS7/jUN7uk83hA7v7TcEwqilDQANfQgNqbYyGCfn2unMsdqgYwarQghfbP
V661keEAl6O3qiFzDMs7i/Q815j5sZXLwYsgxNuWDoaMOAdGSQ1l3Bx+HOTnVYU/
1OKy/qm5zUCh541kejB3lQ875mtvTQQF6w/wqxhNdLdNEdWQ6/DTkFYNavktaZtn
283el73Z9YS4uS+kC4WbKcn50xalj+4FSN6pKS7boW6t++eCgLMfFEas6lAbSsP7
igLvmMFCjBoZK/5ajTxQ7Bn5pJrBESwURN5gjnzaD3rhvYiunlM+6S3EVNN6bwgX
NRtYYb69T7Rp9H7JRydXjslj9pzaUZU/9iKQqofHPA7/NtVtyWol//ni1qDEjqXz
UeQZXGwVhszu3TcR6zLYamkjnW9Hpddf7vVWp7l+5V3gE8o56/Whq1fiBaRD252j
lGpsi1/z4xr2/O6T/IaxB+U0H+eSDJfsox6GObKyH+OWlbuAxhxV2I7K9y9+rXSR
/EmMx7D3kC/UDF4zjgcsN8DX2IVNoe7cqvtnQJuL4Mjud3D9Wg3kOrTr8YrKJ/Uc
bpT6FFhSLjXS4B4EwZMwCoBKexOpH4O1nGm3wCj2ZFjtOMSk0ZmGRQ6sCqO+gy/l
yo7eNqn1f4u4S2OsSP0OUCnEcLQyLJdyxCh4DcTwX3R7rtE3jS5RF1uGNIalWkvQ
Qmvmy84LkChFvD9GtwF+RvkyPF401OvPc1++6C0k98XZlFUVCEKJ3bzsOgc+qmIu
1o7elhCBcTJE72Hmc6GUu96DzQbC4rueqZ5yaBRGZaLS28MBwbC0iJn0SFQzHjdC
w8x0GgFN6uEhp948qngozQK0ABktPPgtFaoRwS6DBoEpXnnkbWv7O00I4nbV2oQ1
IDSC8Qnn+00yCCb7r+hFwrdwqMA4L4lj9PR4a6SfVfSC1NM99NBKM3jHjxeNOs9C
4GZZezvsuljXfwDeQ618foXmShxvH+S0NGgHX1y8wDdsq5D3UUzbpNBOIY+L82rU
gfsTGi8K1UaIQzlivkTIPtWEFWDhLsYyUsu43ipMGUXVd3CRtcj20KBWJlmTKrmN
rlUUQW6XfbujdXCAiKDTNI8ob77Rtyo1iEhvAwSUUKk2E0vwI5qNjmXpAW3ivy1+
HdRV2qAIjCAw351pNRaowIsHLezZ6tGdFIJHqp4o/O+JO9bsEpphtlDWHAmVYk+7
W49hB1xrthyLrt8J8tOfeoQ3w4DTSHsc8/2zYKB1IkfgQPw/sMLoTWO/6KW7ADa8
xbqQpAQ/tuLojJaRmVla8i9s+TU+k399zXg4Hsq3NUW4Tpo3B+va0VUeuFiZmT7Q
cjvFZ37WXdrDSonxV4Ire9cgu/lSdamp+aIox+FnvzXGUEhElTogJZoDsZuGRmfB
gJ3fYrcXDFRwuBvEmd3qZArY8tK3YAeF3fkSEa1QrxlvLJwBel8o5sm4uq0bJNDy
cCpwZEjCTklfydni3B+E5crtQcXaW4imv8q1U7JE3clKurYpSzM4mKfaFZTrCRYE
I2PPYCxZPHhE6Af62BOBJrna3PdGFHON7gdxm2h2ITlGDyumaIsG6QdfKPPBPe0W
CGvE1EnDJvamBFh9WUDnKqI0/Gogc90IFzGK7vRV5P9I66hCnR8PI21kZ4sU/BXh
mrvDDOFpv5FXy9SU+Pjj8GlImO5kXpkoVF5jdl9hfHPjRgXuo7DtCY+qBtFtAudd
TRNi1HOBb0Zl7Du+EN2XBkQIoeQQmviY+8LU8kO1vih4HkT8t28sbXnbsonqA2l1
wQPcWFnjgsszamRJIrce4Pt2gDI6gkYlVvld8wNtwan0hiKEnkFx9hcLMD6fUjEn
I9SpEXSuhpHUqreZpqVoS1t5SLAEaTLflirEPJuwRzz4MeDcPDbd/wtBn3h+v2pi
qEJa7cD+2HPrZStmikO7SyoZUqz2x8AinQ2wr3f0FKI7zj0fal72diE9PcYfCjiB
BK+s8/O6xMdSzFiCkwTD343nWoeNmH8qb5BkFUtdmEahTw7eJWMA9T71ohc2geM1
u2Mq6FGQeSMPpyyCukFKBLfAjbLL/r02Sjwao+Tylp5o+7u7zRPqQoTpzocnkYap
HvcBx4uBROM13jvgThm8GP433Q4Q0ssQUCmdAeh6vJFUjbgWtHV4X3qJzFZf++oy
jD+iU3YGDGZouJShhTA7jnsAIVZkV2P6W6RH1Ri0ZggOo/wcOkQ4Uw40K8duQmSG
HhJyVboMvufO4DnZD1qCEJuQ98UFgqVZ8XzVYpPigYrED73H+xDF5jnXIOOi8OWz
JWnwDJoDx69Vg9vRWJrLcDuYWnklXW0FUookwqs2NXU=
`pragma protect end_protected
