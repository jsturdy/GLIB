// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qK58Dkx7CVNyUDg/Tz6uUMsF4UU94KM72RfcAPolWY1dSCChl356bLV0/YeJTp1P
LrH5OdNHS2Zq4Tny9N/r4XoRBwWnoGbAaTDfGRazN5HLdKwj60VR1CRdsoqwMhqs
3nCvZJLjX/PI0gvUtQAJ08uSsMHAFXTIUub/dHbid4o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18800)
zKpZa6SfnAbnuS1UJxQ/VAZQBdlOmmSBoRpE35P9LnP1YjjlbwvSmwBYj5eOOCol
7B8wPz8P1OvNj6V05K99iip6NpQEcxU+6S4TFQK8OuWVp/cdpPEAtQLww31oxBKB
s2mM8xrblKliCAGof4Yy3e/DNj9vo4lIeJUyYESmb9t5Y7M2/vJiQ5sJOgF9HkyN
/AJ0q7RJTbcpUpWi+J9lSaX1L3LeB5uQMwk+NORPDcCScKyIak70Zqbdw9rI28mQ
Nkgp4bD0F0ANW+Ug0Uc99AHoQWufYaf0gQVxfpeElwm5c+27wZAc/o0IQ7jRYzof
NqA8QvVMlg+sr2G1xPhk5bnk8ZZvWyUYz9ennZOEIxuOQoN3ufxUG4Bw2iOrpfI+
iM7luc0hsQHIrcx0xoIAlIQk+CGFwvdZrIzWF/8lf1dwOHsebSJ2EoHtdfifZg51
c3npcil4ZsYEhig5lnxzJ4d+q6LZslMA8RolWys4FMCizVxg1/NDBYKDt95c+0SO
5Pg++zP7tyBYHT/1UZkBKo0fWraJEJRSq6E03TBJEwT/A/HnyVdgH+lgA5707Gk0
BmNqg1elum8UfRBqFLIuGn54oj8xOVp4nGxVzzwjyNkxUjX14cKTJF8ZvuwYAODl
9ma3nYLtxNe7FOWpMKXll0ayOfLgDZI15njN8IREq6L59Wr0d3umYbzmc213hmhv
ijDDrb+GLpnpYCckcV+N+if7Tv2cwpf0vf8yY0JJkgWczXt0Kcr7knaCfXoWd3Il
Q24ETL8jAkoReYY6uLngnyPwm72ypwX7yjJJaomyrH0UG5JtVNvtqhNnOclCXker
FGmzD/G6hOHJqaD6R4ZcbTXKsosICMvXKknelj8g7oAEKExBxMT5DyxqB9ZYIZ05
H4T3VdfC3t76MVPdowp8H6g34wQZBC6GQIQu69ZbvBb2uQRPREJJdr8MD5Mpxdht
A2dLLays+dXUTnxumCYImnChK3R65X267Cjp3t8QVtnB5kJynDVpzeiOdqEOk7Ie
MHNPvfyRwwz1Z3ze7vS/MmuqUWc+Bdx10TIgnOkHmcHEXnBhCdyhijOJUYcuBs3p
Dhg2zTG1Cy6RuOi5HP2KPQoGR16KvT7E54v2Nqzsjf8UVA1bb/6WGVi3Xb995Z1Y
WKbFljasy4x5WuKmn3qaLFZTItLFN01kkBqCJRRP0Uo/GWRMMXPp9ZQSGZWq37BH
+A2ctBx3hsO3jVYGfvx4aPut+v6r0y2/h3OnaVyPQarmAcC9rE/RahLpiCh4fbpy
KnleEUQNEFBm4BqdLCBx3IrzmxOG3BbJYO2/bF+doXRQ93Vs+1HvIztI6tUFgQoS
lY+S+1UB3GPoLjkL8h0dsiRjC4A/TPD3v++caE68emMsg9hNUv0uzYW0F2Wcll7T
K1H12JxLY8cPkuV4QMm3O9oqvuDGTRVjFsDuoZA4P/U7MPGpscjmgtSHeTJecU/Z
5d3CpGT56ZrDk01k9YenI90HL61KMNA+zyCui5hijdhudGEpao3mIr1BPVPTkCOE
vjrrg1ksVgxXpV2RckA1bOhID5ZclHVl+F81WMxongidnGwZQo1BWUxA0c/myZU2
WF/OGi657o5XKkomeU3qmm/uQKx3CjemA0FIylywN4hbPRUTRAJxRcrfJukyeQPm
IcbCUXfNNqlLRdBrNOt7ri0xrTklS1reiPQSn2RgsSrp5sztftgBEYm7AMpcQ7Nx
UhGJ9dEXxNwCH2GyPmnsh8lAYAZYHtHSye6zznnH0pxDT+sIqgje4KrC/Duom+WE
AaaU7zyG1lcOJrdA54g2P5QTo4mDFgucF3tzT8aieAXNgWhI7WmoerVzL7MZWXWv
E/L5rs/tT/lEOL1Ljw9rbi91iyPeHDJVoz3tvTfGjj2pktgZPVyrZf0gNsB6GVPU
iItI5/7Jwlou1HySFxx2AsvcD3wDxkxuh2kL+dNe5G2VdYizyCjEbVWKC/UmcaM/
gJJmx4ggRfGqP4ibUfJQJv7J+GGbH5Zdk/rgOtrk9MC/i4/oVRuScZdLBQRAkdZ1
XXvwsMtqDqRIIxJXlN8WADtt41lfREsOaZLcZfcT1ZSjoPZxtEdTu24aSqv6V191
BLCR58zy3eCFLWFye/eW4UUIbs+hkAMbiQ1315owkSaUaS03EBgQA7EAhlsDMhrR
/wL3huhsZ4TbaBWYetHfRkV2Bxkg4Els6ciet2YW8vK4nEdoHreiCFw9jtZXvb+A
LmT3+zacJU5f6qJjvhQkVJVJaWviY9sVArUzC8bjqz00DJw2fshu4rvICezSGYGz
bbn5TcUsbS4n50ETcCZMKLy5qQOwwqXK+ZzXRPUpmMK/yVNMy0IdMlBTIe2MYrbG
xSG9HP2wGBrUurT3LDR3yFh1M+a6XwkNPLjhaag33auxnWr3QsISBoPqvFaZjShl
oc5V2w20zwDAvnnNj5TY3BbXGqtV4yljIDaJhbDVMFnjxJtOSkT2liBfrEIgFRA5
O2qYxHreGGiAim0ZJGuhho/0arquOs34A+q7eMyuLylUdGpksESOJ4zn5meBU8x8
ww92i+GVHskYFn0qUlz5fXQlHWlxhwR3o24/M1ETkP3/JNzkIF7BrtR/IJ23gGlq
cMscXgF4nBDraQ1CHdundKrLkmCr2GuvQ1y98Bgkx/AaWzY7vEPxdXku53pAk9Zm
i44u8XCUiRH2ayASmilqIWjKXKn+7ePOkKpxIONWRshLBvCivhc6XuwuPwoCa7ta
HNJo+A/w5U0FLBVoxDSeLDx1+8CN4oIL2B7SOuO9U6UtFy7M0zTZCk3no5rZCyEI
zzBTmcI4Eh/I+p8ldNWdqGx4PbtJEHkz1zKaDY4mifbANNWlmOgQ7LxcqU6eefpp
bJzz6sVahyQjANmPA+CRT98jguV67JsTVqPlaDu01cLT+tHQ0Kv9T3wyHDn9LTxy
YH/jEX9qK6dQ/kKnmbSiv5pKfqQsz6qtlh5zxMRXzRI0iTLq0Mf1wkB996HxoejQ
AYVkM1pLM7pFs6F2xalu1QRteZ9hQoXzXdFVBEouDQ/JY+w/VFrGdxvwpBkwUiW/
rT2mr3I7IPddNSnPqoUzdcS3MP5jHs05+j2JBO9Z8DIoIV0C6cQG9GXFXYPMx6/a
muh8Y5OYAnLN4tXdti2pRWUruEpgKC4ty2SWb29tQ22nd36ygvafOr/sXjRlD9B8
GSKh6SAl6vkCVjRpd+Hnlr1k5axujjGLlssOh6dk8dhpzLr8MLhcSocI5mjfykos
Ibb8ahWBelbTUUu8y6IZLY/HtDSWOOUtKAp1PW1E0Om9WrXuSjtKlhE+pmazGBcG
G9e/xooPATasnEQSHHYn7m3+zUJyFWlgoM3tm5jicnyu1yJycuVEkROrev7qidzp
pxkKZz+D6SslIqYm8wHF9Ygd5mQFzH8ubmkxA3py4byQTtvdoOy+qL4qNvmg5+eg
y06xq9rgvD+qtPqcbn4QrSv0HalfLz8SD68uMwIQqy0I85i55WEs8FGGVXlaKqwA
6qAlBww61y758cO0DUl2nJt1E0cRC2gsJyOv4TnFlQlqcLOpzVgm2ke5JrtRGiyU
mPPN004w9+EY9gLiWhgHqbTjd++b+UbNv1tKxUr/q/m1apfSdkZxPhziYt1MuyVr
uqVoS98SCgrxkYFSmCmGBFd9WKinVYiJEgZ69rZ/8jl7lodj9POjXplmkw4uIGay
yB+yeTXWhhR0VjQVmudgfK8i0l8671adVmplFVfZIfz3hmeYQlvGe0+dosal2z+t
VQSykkkV7JRh7fXKqPGX/2TmXkENw5GJJfmkdKSOvxyhwRZZTg1mhAANzTDpjXd6
JfaBOpT+lKzpcpqH07CIDV8JspF/SojunOFjg+5YI/wZ4pS+ZGOxA8Eg5fkwOeBU
Enn2fVeS9ZUfBaO5rB6jrt5qBtfuLPYjJDRSSSQH1I+jzFgaoA0Z4TcfxHvpuuEV
W7DCWctuLp4POxL2Qse9sByaUvI9fanaTMibJjJIWvuZcdHAen15YcCuZTVO39W8
LVqt4EqTKmGXgCP5r12o1nOxgnxstrVJHvTPuc0LEJZjX+lxsnOpuFoD/iMLdSnh
Zu6Dzbr6jWj421forpUARX5zB1InGPZFWjPmtHkPyuxuRDTU9fl0RDK2KLYhrgzv
lakhfKW6b8SAG0PQH9li/poXwBJNAQxiyeSP2kv+4lbv9onfoXz5cceP0Z+QnE93
EZu84qikzTxQl6SxqauGFwS0aUbAR0PfvU1XSwhBByy1PpwD280MPVHSiG0g1UQP
otUTguDAsPVz6QNLEXNTk9xkUla8NLhQRFQVPMfS3W3pgorikiDMuhrRcDP+fLfN
czvcz9UxpI2NkNjm7skm37rqW+stbsoVropF61HC8dLc4xWRulR3cE/2m8wHHKHr
O4lbgo7IVTHIWzFIaVKvlXcWT22vIvC/gsm3aeLbQU4B+vqU2y4y8V1F8NH4IPi3
MTVvB1rRhZrfSVuH6h3/d+u8e8uQumjrsUs5DHvZlAyj8XjJP5PV7KvJ2aQgGHlH
S/uxx00xHHA6GhX62tfyto+5dBRxNP6FGnufz0uVR0z5MdRWCPg3jjLkmNBkx1xg
M7ztC3Gdk1kpDCOL5/SVYLCIxl4pQovAOwrhWCfMyYxHVqMkxNFNzrl+ugCqoWlq
m1rWZJfmaZxKcaTsRo4YbZK1uQcMqF5WDuq7+05AdOI/ArlQaPZTlAMLfT0/g0iS
gEpa2Diw7QCHXv9aNaufbPvxomkn0g1NYkl81Z4iXr4YPtuh8V40cxwe2cFd7iRt
QYB5IerA8Xw4tUEIcKnnwL65n8dMredGw+j+EELHZz5f7a8FeGsgljEyDDlIhXD7
dnBCWAywfQ+nkz33+e8MyBxglIsYLAOAnRMhkvPjIJxaC1EWD1UyhEm9eWhI2Eai
MZihk1B61i35ncjn/cAFcJwhZZDd1PRFUmNpbjK0qZO0XXG54u7r/695//SzhwHV
KwtswIzVmpSlabp6JtoXEtvNVGiNkIRd2ERTLOvc7gTCw4mHEA8Qe4Mr8LsJp9A8
ieKBLOB/Zyz3U25e9uO3EgtrJ8JveYSoKEIgZsB8Jxzsve4Dg7buWq9dcbWwb/pK
NT+h6XPtWZ+A2TE9tYSteHQ+qUs35PZAVipkCZHSDgre7fHfynpv6RatdCO2aYHd
dF2ApxaStSFNlD0/frHsk/kfsXdF6PYJb5iCcfIJB+lCqWGRcaB36LE53rV39glo
Rls96l0Ad41poc2QF8tXD9Atxq7htT+kXgz4g1PHdvQAf8BcoJl0NoVAsws3DZHI
/oY1nF1DaxFCdUXJ+pjtDP1dmUoM4U9BgcupiVSU9rhHVo/pNi9I1LjZ7QRGmWXv
l2dWjCkUilTzpVez+ACiDqUb5tbp8NwLJ3Yr1JImtExjG/vqFCYoq2lkuokT3bmf
8YWPaE7v5/7Ox46dmILX83FvXMtRn2x9ckCtwa5qFk2otZwW05o2HPp26x0RmB+W
H8q+kSNuk70Koz2lY8YjtTmJV5KitbWHk2EoTV5Uxdt+Q9M5K5gNOomTfbH4AQGG
bZD/SDtaNUxBbRm4XP/5qdX4YhuKCgOD5PZ69U5YB5TvCtImWvnNaz56Wa5IG0GJ
Q/pHn7iIDuzvOomhbWaviG+EOARgbX1T6lYS3ID5dmWdAjJNXfwYBupA1rpSJOU/
/lDzQbe8IG9lBbXG6QRqF/p14/iQLnUm8cujY+SfIkeg5auTqMjihZYY7kb5eFSS
mQ+ekC89fPKmJwhPi2904VOoLNZlbt+Xx6AKX5Vgqh7XK0T/BR6XRXBSQWbZQ2s6
I3GflktnGh65CEufpRUJhxJsVvmnWLNyshiVV1s9FAdD3H79Q3+kp2oWIcFfeUlZ
nv2Rbx+1SQMHXxGUjtjMiGJ2V9AndjDzKnQrqtM1lbjhVwVOnyKCwIfUJFpihcow
XB2ZVo0Zp2giWzBu0dNGs1VcCb5M2SFY027odRuN9qXDJfiUKCrq6f3gmqYj++1W
GbqmcZdq3iTMg+ZyKszfVygjzJtR2twb5JB9Ywyj/bvNNt1b/FJ30PtPWFAAKZMS
88fvTFA9hYuES9sYJ1Z8D5TWpf9YL9zKp4RssnR5JvrmRh1/Q20OmC2spaBpBhr+
ZzzPRFo4EOm0uIz638zOJUUcYeTI2r0ausAGUYCWcTaiPfzE0y9kRIfInYJeMt7T
E2p5IyiLCZf58521Ejfh/S+AkL5zSy3kUFvkOQ6s7YWDbWXwOEhKA38ce7VOL4MQ
aXv+JANMUKslqSIUEKZl33qmhLBW/5nVIM3lzXppB8yqgbVwBGctaikQPbmmyfKj
2XykJ/37wKJrXdclHiVgItZ15StXmROxgZFeMPGfDhLoXiWpSNBsAJuJjYicJIja
xUTSUVSwUekWsZedKZq3RRlQA5+kcI4nHyp2IS2OcjpfUODO82P5eLEjBoRbdJ9v
BDHpaPPDlhq1biPadil7dN2Bn5GZSgKYK4sW4SSMNWafjqxGc1jDiAtIOcyp+IoJ
m1Xz3LI/7LzwmopVS8qAcHPOKt55ozH//ZvUxVfNSOlqCjtEmjq5VNDK4P8QtuW7
DUAj8CY4iYrzyxLtvcm7SbafFzHc/lVY0gHMN3noe/8+ydTk+pP3vfd2QFBNRfC8
QrNj+7kSx7yABz1PORwzkopHvzHSQUeQbsRb/XoICcwy4CwORlcJfD7736BEF4O5
GDo5o1EmpImQjUvqoYCNby86Kk6qBlKkoKgZ2QZwlLcpV5vShZeFvnq7/jyL/TfE
5acrod2tfSY4NFo/7nahoH63N/12uah/I+vT7FdnunEnhMD2OUU+ALljaRMGBcq6
g0I9XI0R8khyFWPmTo3+EHekT0Xzw5/2Nd8mg+s1J7p1QTbtDYUrfS1oqQPgBa6i
W1ylE5cASjBjitlghm0r+77UwI8UDOAaKk/WsYGbf545UK8sHNd/7UJwGC369E7U
YSVxHXkHGbKCDZ/m1Wn0brEqIxuJSKdzpx2yoYUk3fh7v2ThVh+5FUAegXsKjNRq
wY3a6Lxe7wmwKBJk7bG/8JVX9Yb9ymjkiy1C0Zlc5+cFQ+Q2SuFHxRaJoqMHYUz7
bd1rcFbhg8ikRsNaADVOtXXgJfRQqhDYAOGuegJ6oyglloyCkPRU/jnRa3RVt7k8
1pJ5PITOIX8gLh2ebVtBEKTEj3YljaKE0U92v5wJgE/11Zg3m1XkJHAtBJGzLmGB
u0h7Noipivj3VxSPAiXJfRadczNilsTLMu8r91Xui5IT1knWSDJjVdZFkifw5olq
VwyyZg3mo8QUr1yiKGTVS3/ieirce3hfdaQsCqVC7YVu51H+LuuG1nzWmkMnCRdB
cayprsQ4MYnual6xu9VTJklWG3BGwyBtHpXNG1cWgRIdB4q9gvw6EKSoqFjLG9ca
+NIRlLZ1kXfowfwDRGMmAfmwnCKXboJL97ZTTb99BEiYtJKY+KxIzauz2umJcoU3
ZYw6tPmL4nGXeYKdTmd+f3haM4/s7u43kl67hM7NcB290MJwBITg8fcDpMQ350Rz
kSepjnEAh/ENf9wKxkrZwWXrhPmIUpvwAjHq3erOXjDZDJeZbsTmj1ozD19GlKNQ
mo3JMJUCqUOKbHqI9ptoVnugPVWo8UAewqoRp4/zyfoG6D3tc7CHDw7PhY7IKdLQ
S8nI2aO+ZqtdSk0qFCRdLE7PLwHgDibuVP1Kj+UfmXoSCFRcYJAYddpW89AtxkK0
NMLRv3nATtYykdNc2ORHXOG0jeSrxCfsLHK7ciHXyLVt2syQNAUnLJXCJYyQNR/x
LnrQn7Gao+eQ9c6fbE5aBfovyKoImwBy6lWGLsjXDPAd5C6Q74r1lo5iObesJ+k5
VM7aM3XJjK7eQms7dV0cs9JeS+fgAMHIL/CQvomMs/4vXXRlHnmmK0uZ8uJCDzE5
lM+AcLvfg7grItSgXGfQ9A7hVkojzt0zxbsXB0Kzz8tJ9hEE6oLGHbGQ/Vv7s2Ad
xPAsAaPifeDeJTRGTOSwGH2xMohQIORsE0C+0+T6hclGjuqxVOepXoJ4Rennd5V4
ubD21UJu54cEyscy8p98yJHH9MRy+NgqM4J4J3+Q/e9734p6GbH0Fj/HnUY6xvDj
Tz0bJzHtn+XN/B9bbMWiJapth3u329L4h/feL8v/Rzz0j1Q9XZ2gSIvOt57cdwWs
B7VvP/dnYzOgpui3Ittf63TFrXExQETeRSi5FpDsaNHog0eR70Q7+k7WChNq/giW
DldVEyRhudzB8sUWvhdX/g34+e/NOvCtEpt4m94c/3vW/GGDn3Fh3ZJ0Hkxw1ZNO
G9QLqdXsIWNtREX0gpRjo0J68R0ZpoC3r8vOglJPIcUtji4pgxPqQUetA3Ae4GpZ
HFar+aN3yXEcqhHoHnCYYPsCQxz5FAXXkDdbjNlyeGkzGvCHRi8Z6LzNNF7jYJTr
pYncwZDt5fNB83xDcTD9NcRGBnCBWXNixbUO2VTAwFc2K3gPwwuEPUoVPmF1CfxX
lfQnmIY9EkYb2aUv6tClpgGRomKZ1LRXwN6+ZwxG+79a2Cx7Qg3DR/rPKUc3vlLf
Qe0uoAjzATZDIOhueGiR3hi06Df6Cuiyzq6tbq53Zdr5a474eWpE4J2rIasAJ4mI
yRXr6Ti6ErL+klO4hgg6YKqyBunuNenFLdLcFyLP5s8aHcIHtG9A0OCKyWrFnG17
JfbItbLC58ldL1cE56sx0u6Mqw2jlq5dZIy9YFjDT0QpI2oNjaLJFZIV/Ufk+HAj
uE0QKrVu5cNHPw/CuYM7NJbwZnA1NT/Ei+ASRDkZeCr1j/RqMGgLMWtxMG7MJGfk
k2WOPYatvn/5G2Be5SQFUw9GhnzLQfWXMrLftukWLlivXD8dzVMUyV/NVwklUtYy
WaWTzzWHUvb9YOnGKh62swky/I4qYYaWgM7kwrtNYYwkha2wtfqPRovZ9BV6IJx+
F9PiU36etkIwBvVZHIXXq/yjl9OLXECXPW7VPWxo2XWLTVsUjqx1gS2hcDWuZQ0F
2OxTcdjZZjyWPKkvj4JpXKOB7t2BH3jbWQ2J1/EO+WAxFz1MTFddp3eSACn4nVr/
fLD3QEd6okxYUbyRFrmHyveVpVOxKCSUpkz/nXzWB0D5aJyE2e281vbgEeDFqYxe
gmkDyIw47/zDcYsJ1ycP7mP9zOOLSNDpw4M0rxtioKFNjKFAKoQvSOir5gBqIcAM
ir6yWBDTNOLyOpXSh0eZ86dK+/U67U9+Y2PRiEjBa/uu3V1oQcmbj0E3Y/wW4Eoi
jQtZqtHkrQU4O06kgOfbCAhK9v6Rk1zUyLPwXhmMgTEJ6GHhKyf5EI36RVJMKMbG
bdTNz2DcTTpQgHoZgn39jXv003w8j66ZBkZ2ikjkpPj+JgT9Nt1MbzXS2ORP/u5Y
huqXmFdst3Ia7L2db53Ly9G8DCSvuqdYkIZiH776LDwGVVwj9VKxmbzvP/CIyivn
BuGr197gxHnxOfy213H/FN1RhDnp/8GanNiSvDY5E6PnCFuaWap56a5y15871sAU
rv9GaZ7RxLmw/Ct1kMqLCKNDPD0r/GLLIR7WgaBDn9PWXoimI281mmuMOf/ukicI
La/dyA3R6tvf4uwDJdQidTlnuo27uoj/krsnJHJhcHF7cbc4GtbbRqGHGst4DUZl
4Az90rJJsRRbnWUDfoR0l7ShgJjcPVrIsHoDVEGHn1UfO7mLFkCx4MahlI3gf4mh
xKp1xhf4HkIdHXtLJtVsh8JzVToQOj4J0umy1rPIoH/E5Wt6xaUmCEdfRHXi9Wd0
vDORDGO4p7UL8O1SgU3bUXlGIt326am61G9c32OZF70s9JsKFIIDJQM5rOymbg/C
yr0MctbCiUyWGIeHLHnDD+BKDYSVCdEA/gNcEOvshHjgXDG4GxHtDUzxVa94mfJ0
oSWVfpieFM0GN14lgy8jdsyW/tldtGOs3tWra0FBt7A72zk9m68bL7fJsaGQ7mOg
oZf+3iKe+zMhGraoFpH4fWceatOHTxvFlu5UrXQEn/zdrBrpUZ79tR0Jp0AFp0ik
LxLYeeNnNKGAY+tOVHz1nI+/IZMTjmoC2UuJbODjcKnv/1FXsvOy+IwOfeQ896Kp
Fiwza7+63LgzEj+4Os8Ns56X9T0lbruBIrYZdNAGu6xnJjyuppWL9gqs9v0hbF7y
Rt1K62Dsfi2L5ehHv+CArVpwl3l8a5Uw38M3qmMMu6pmY/pCiUoHlEaRoPt3VBEy
1sP6sugggZHkrHIzRIjukz6MoZhJC5u72MglRAbEIRPBRm3EEt56uW4uFXbouCyF
0wkXA1LMOSspAVRytzqcS3L7ioRjWU0tj7tuZK7Ym2i1WcymPvNGgzQfnM4qxEjb
lwTRtbKZQHmxWvFb5tuwiYFrgeRJdih9DElpJYE83POsq4Ou2KyFKcXXvw4O8rXr
m8qqCJnknzZ2rC/2whAYiR3jP18SpxxjcziHkYUJzRc00U3WMe5gJnQfZV290EHO
hLew1bgJdNfomAZoV1RXQTTSmuy/aIhrbNvU9HeCWxOErwcs6geF9uh58GWFQwdh
nM231yxeZ2rp29gtBeqvweRHGcxBhwd2yvYQukWeNgQVSetGsQUz6APV2D3XUh7W
sEL+vKeL014NRfO984XcroP3fYGck4fD4Iyt4vK3jW68Rpf0wJFaSBUQ7+41XiEJ
fobXjqUSH/EpERRyDvdOWQhW9uo5Jdic3By6nZA97R6X9l270o/xiC4sua1wmp6R
Txx9/Wa+ndZGA/W8gfbGLEvx/7LUsTeelwVuLaQUkNI2ASy1mJ4Ab+emaQVZGUwR
Y0kxJbV03TBpnrjRW4CmW27TzvtitWVfZKVD0ezC00/xL6YfyzhmyG8ujrRYWl6g
qMQji9f3A7r8ZJjbM6GpAEvqGkPEve2irhpfyU1E0pnHbYab0bBgwgs409N7mjD7
Y88fKB+2Idpl6rJe+Vgr4y9YlTtTahKAz9mCoAkOl5XCZ0O3deceZ5yHtjaxsi5Z
KqfP2GNxDhFaedDtsyurFOg7MIr+7QSk7c/l1EvLoz+gQXwph9LG3P0gkj11Rij1
PlTU4UgSS1oB7+uYz6sJfSB2NNCNuKdohRVLZ3OGFX71tjMDSYLIaCZmiR8GSO2U
q+YjDUSnD3/JzscAP1Mll4lRRK49r9jqrAJftJDnZ+mgGMF2DrMqar8C6bfZfiqR
mNDLlJ92aDwGQYn7hqNqK25B/qCuQDI86JMRKJU9QYLCc460/JlfqvxG/C+mlYqV
zwXx1vBzDTrfwGCYiT+bnE7f0pp/bH0V/tjAJTghqF3orfjgM740UihN26EhJpZA
ynapMzc5r4vtH+30nNXKtipPAvK8luz+DxkkmvA5NEpj56vObEILTYYWzIOOggPP
SN1v+1/xTG832rjflI5JJDDblupSfIDCwTl4ePlqrWmIxaKtB3q8Pk+IyxLndunQ
3DxsY69MBQYkU8XuXVAVoRQEbf1MFMVDb2m7fHnJRt4TFqDjoYq8eZg+Yms8UKSk
Yk/CCmlHAxl790inUCi7VQdn+502JUB+LcbcSi42Hr3QH4EAxxoEiQzTBewc6fad
ZlWeIYkL3tYl+BajFRM0sgXdFCfHCB675cHBXFiEMmS68RfYc+QBEd5x8Qe5vYg9
F+BclejkujgnMOd+CNxZ3CnD+Clvi3rYkd9Zkj6dSgOG0n9UGct2ELr/Y3NNOJlZ
2HCdrMjt/9s6Xdxmnq9MD/ZIENHu/wWsClCLIXz57jlvORVadbJPLCoYPSc4UIXv
/aPPyjwciho+6AWB7ksy7GYIUeToHXiU1BLvZVEkA8G5PHOTXObXdNJREvF4/Fbt
kTeU1niZylyD9mXDqHI6lX6XFlnGOcKbuuVdajxPhlCKd5cJNAcAz2jAUkSy1Kgq
g0iYehBOLXYMQ+5HCqaD91XFlKXOnybaYb+1C3WZ7PavroYh0VLff8hpMFBEn7ZR
dT+O3/Hn5XC+boxJ66TpC2NK7EkVCh71fSJrz9bLeI4bd+UKQCDzxxas9O5SMjv3
IM5iZNy0pXGC3kQoVY4ld2KdUFm9RbOzbqzMpzSr9uFFz8uikBOnQ3s9cs03gn0D
C3Vf1xRouSTND3b5l3/vH1vO/TsHRejlpFNzE1KavaGrMm7QkdpCPw72vPOtbkZC
GxAtSStB28rDQnXIxV0YD9b3Du2HfPz5gatgVe4RameKm8fYeWBxGKclUAlSNcYy
+k+PsY2lSN/QZrIyUugTp5u05sDTWRv3N+lfrLiEQMInPaoiAPE9+HtyB85Q7L9m
yYp6ONInbxgeBv4l4AdbRy0VVW27tY6WjCXx4mYhh21yyjz7Im0km6CQGZZduk9H
UYlwXVLZ9xGSAVo3goFpqh2mbiqA+/YM51eA+FyAYOyVkyQG2zmhectnhnDb5Tx6
bE7HZ7ZZXTirWLG7r03dZzdLE1YiRyqn/QM35OIktKDO2UOeW0fiM2yGgXpv50k7
PipMg1cI8u2ZiKTRa747P08RB0eVBiYXDtOws/mVTkjsfejyAicoW7cY2XckJOpY
vgyaUGluJRrxHsBzgUmVgJSO8Nxarp41Abz1rktlhYnL4KKhZqR0w2fZDw1dnHYE
F9/k+zfvzONAq4PVtbMgHYy52IlqD//uzem/4wgQ5Ce8MPOC61ASkYBAXfi846QE
Qf7hEpBNJj5KkitdmbTeuk77NaaJ00+sgp8IC+cw5waqOY0nXsbBjdXYrjZxmfIS
o8teyV7BEvdCTM1KMZilMVme/h8QTPxdtmv+MP1YZGe4lC0/wAWko5R1bnq1ZzMH
0KoMsmpz3znitgHJ/eHWWXairqNNFmW4Q2bSMxwdWf9NP/V+vMBZa+eHoxd3KFbw
sAC9beIRxvjIc1JKf0wtMEbfvqpBv9P7Zwt4p98oVJAlRLSl53JlCdfAocaOZP90
S3eI2usQ+AJEXYcyGeRjFijdPzaF8kCjN/xrxL3Mw/8WJuQ5eIizkd754F/riEK/
HS80/CyfoPZ4J7RmPZciSDCMPrO6fYPT3DbLInz2soLwxS+ZRMPTl0r/Juf5Y25b
o5cIx46ME4jvLmWKmwYgQGa4pH1Xm/p3WavFVavNVVS6g8Tm/s+UfQAX1737VgR5
Fae3tHrDgXmg67gDG8X+bBfNYcHRfPiGFskZA62M7WaTkgXHR1VP3Uq3GvsaF6T7
amfYufyXrxkwKcW5CceWhejGHlXGAfWYZe+1qoUi7EQi47V3AT5bBWhVCfr0wS8Q
fWDm4r6sj6rnFcapHWTMzp6UXB/74S1PZd+pCKQTlpFJ3Rqt+efcV1Ul94PkyjrB
0NwOdBDkGD/EMXULbvWhg9Z3yl3x+3a0JW2Q7RH4aVFxafZYre+4lVZlhNZCOwkS
JbuUEqKvWXdZv1GY36K0ijdjYuUqmM8cNaaUnFOhdYkiZo9wwQV8rMhBpbkC3yYJ
xJjloO6xWM3d+wn9cmZBrk9isiccSx7FjEXr3cuizZFje6NN7FhToN9QM+bFdsS4
YaiC69/aJ0yY7nYjplRvR93OagoNeW6p354nkuyA0tHQTh66f1lBZTUxVJuPj/sg
3EjS24/0t858sDc2wO4GQfQbZmnopNCxddNhffjgHCqLM4gor1jEY4iBeUzitSwp
zLWMcv1B8CnrDEdDG12EKbq20/vYvXXpUkku4N8pw2NpxLOTekLwUT+9cd1B3wQC
ZCrOGi9yPhOyA4xAvHaTs9O7jEZ5CZ9OuQkPibbserdKRh8n7zB8C2iBnbaf+YHP
oXPAyYPc7ExWmOILgiveBEl9moUccCeUNwpJwCUFzWaDvHsecP8qn46JZ/Oarcp/
TMLVeJG7mqB4q343jDo0cb7AMUGZT6lylM5eQRUcmepnIZ/hSujglRnL0lWnMhXp
9CKAaMVBL4wa3kxcxRlKlnL0A+BlU8VTAeatzlGnpJpydcQa2EHTCjQbMuw66/P6
GLAgxPTW41LAR9gz9XeyBbZ/+TZlhfEU22Y5kQREV9mCthuI/m4Tfjz0bZcJrBwx
e+Wsx1Iej+NXajp1kr7sQActveFwimjjiSyZtRWsc1JVsr7kB6l7T3vjb1LO65om
Q8gEfLnCFRB+Wqx93nGcHRcly5WDGALKAd1WNmpJByHQuEYGswAtHiaJ4IjIQewt
4dIBhhFcOAXb7fjWns2PrdOrQYxdT1d6zM+amVgBz7ww8v0bRPkpbVPidsCGo/Dy
102JOTwe/8UM8hMdImRj7Y4t90IZ5uHRtGnHr4oxw8wWEoeIgp6mwjzCdQL2/UUl
LoA8cao+xULce5I4rEjb+c1AMYFtEPdW8PVVX6flN7OE2kmq+w66JKyClUoLB7mx
qDFykRFXrI+i/e4CRgpxntyMSdqFpE4b4YlxIdxgFV3v6nyU/9cUM869AXYfCrsw
2KoPO3kAtnjJrjO8p5yZd0NxBIQvmkkhPU8SE9omC8BFOkjCpquJQans5htoUATr
FT1VN8B8ZbeCcjzq5zWaUue3WdSutH+9IwtHWNhqWZzbuHUCVHO7ewVISFIfZmnh
kDGyVA+jcbs5mLpB1wL+wK9w8j2xtbX7PtRcTqWNX8VbsslsFAXSMuuq0QL+E9mu
yoY4GjZ8ozba2Xbe/4+S2CrxJX06sqFfPJZNGAPQXpVS2EMuIoEYzqmhGZcexTSr
ridpa10TJmsCyQBRDneH67CKeLOJwWgYF0KnrConO5Aeetiv2em6UbZbe8X80HEP
oesmfyVwAJ1KPZhQyVMy/SH2uRnv6EwnU5TctWBmE41cx3WA5dd2Cyzyis4Pu5Zk
sScP4/r5PkEvBRtHVX58RJmaPAb6AN2kC57Ikh3Ue1eBVXsGjwpStbT8Jdo9QcZg
T62EvkkHXNdZ6JNo0K4naAS8tin5BQoJ24gd8pg41Dp49ooc+N0c41fS5J/B8+ei
Appx1xZ0bUav4AfqhMj1mS+C1z5Jnzl0zFLxpGATfORmoHC4bmn7k4yWh1Tn0//l
Qx3EZq38BGLhd4SQz53iyINagTF+/yhjSWOYwkp1EUv3qmc44qbuI/2Nh/4pv23V
A4dDLgoAwfdC1ctS0Sg7nAr5nnwn/VNtakROl/YtBD+eGbgb/0y17m3XZjgh65y6
riys0WoKZKCfMT1qPY+LUAKKUUp6d06sZyf4wEfOMg3SZLXc5eZCn+hEU5E76mGw
RNytVVGgBiTNVjAt7cYROqdSLkuDgUC3O+MiKReRcdTY54oBiLPwfozlJmZDE8p4
E+0nS6LS15U2rsPf5zYoD4WEShB8E9CO7XGlQA5CvU76r/+yKdEMbV/l7VdlmwQ5
QTHUuq/zfPHgotZcbTlWxG8SBpTNTZQKxmhg4UYwG6UTpr+d9TE9ZocLm4+MiWYx
njimyJw0qA6zSj5wBWgHLruzwRATMb/Q4U/VI3U41VhWBkJmzSk1pnI9j3Hne+wp
wByJvfKlwU6vBZyqLMZt2OKvMM2UrST7nbfY695rv7aOM4VcjjxaPtVpCbZng/sT
fF3SVhZI1FH4HMSYn4pk2z/C3T7v2BRKmjXGJAy2/0i9jzC6LNFdEZMKz9jZFwx2
C6RKvPtXbD/TZkD9M4chFJceiaTe8MJgeE1bGGk4FwCBjV5LeSaCys0OV4NsvtKv
HNK2yQLT2Jurs0o6Dm3t/K75A8L9nJzZQQw0wbHIq6Ta1y9rv4dq+TZxPQGWgIFu
hRoXkOIPm1eulquwN0e2URRYN25n4ne4BUD+FHlhmfc9UyM7II5S7sA/2rSMkLT6
NlM3DnEMZyIBuft/ZDHood14MWsqTxVrriVAE67SnM0ADjgXQlmavz++vds6f2+B
6+tdQhuyc01q9CwwqLA+bkAZk+ETzqmaOaBToRsoIKKSKu8B6RIvoUfYFyE+9EHl
2Zp3cVbct6FT4eDooBXUH+pcC3QsSRhBwFi1MAQ6EjfO/ZXdL+7MOiBM6RD97cTB
+X7WeBkptjrLvA/ZTaYResntzw9b31ZaGYZ59A2H4EdtswfF9vETlQLhP0XWfMuG
BSpyfqBOsyp02Ur3kGMj8ftyNeQuP0sjgWvwS+bOcUQVnTroSnTIq2bcOegxk6gD
2XBD/CCqC5ThaW6igoDMjF4ej83EEgn3ZFegEtSFLn2InY+h9GYfXcH/NNq5/jPr
czaVxE1PBYDoaMTFrlm/A7BFJ/DKHciBdq1bYgEW9I7cd9C2YyWuNQorznALPF6g
KE4T0hL+0Q/3UmSyXI40OtPSoerfjXSqLT5IhI8FkWimkyfqfJverZPHAk3dzHQ1
wX3ZV6r0gVkzVVVpR6HfdgF1cxCgF2gbyAcqiPreW+HQ71ec1r7L6G/5x5eELDJZ
NAhr5tDQKHjLUEEjMI3YAdLSn9XMYyGJX6Mcbr1ur4qaKEV0c9S69Ewa3Iw3ROSY
qsnmezo3Z4KmBjCe8tCqMisPq0P+KOIbUSDBDfV2TP9C7c0bPPvJKYZEWbAc2LIa
dZeN2cM7vXuS1i0BoeSNzjf+1W1fplK9nBzSW55HLrvFQYynt68dzhxz87QXvHPM
mVxzdDgXnrhoZUbl/T4XYBciptgTiDr8+39WTdGugKViEcQtWOcw/hI/jZFOEplb
G0xlXgerNm4UIeEvXS+rFKDCJx8ueQ8S4TLx7gV+KYOHnvOt2v13sC4n6W84olNe
hvW7j2C7kEe9+L0L3WYneOGbO2eVp740ni3bP8pREtrrilRhMZTnmyaCiXIeNHVs
5pxFGiISt67QkTnkU6PXwugcUQdYfuG65k01QmTRwLKHjNrVzLSiFzKdbyG1qbzI
2EFWLTbyvSHUoAPk+R6/l4xhzEJuP+oze/LALzUIjR7V6IaT8uQo5hBX452IbUU6
4jQ6bY9MrTubs6AKo4uPibyMz6ZIjIE8sy/fl0Pbe5XHB4YOYQN4ZaBDB8LJzyxj
WQG+WeVSlrDbuVL2+JkyQGQnvlgA3OrWi9dtkUA60m4k1z7x7Vckm6TTGw0YNtku
M/h0fAJIn1z5yCPkBz2F0sn5dBVa0t6qZ8lvQxJF7xdqB64pR8lAbGG98ims7F50
gkFrM7jhMZjpVzdvxPTft18FQ8Sy6tHs53WGzUt3QI4S9Hyv+Al3UGhyoVic+VC5
brm7Yl+OndGu9yRS3pA5E1o+F2/At38SDRmnaPA7AW6E4vUN28wM0H16w51rqIt6
1nUeIojjid6nmOylI3MELnVwbbzoXkGSg/yGooicIxqxT/IVZYDKCOzbGddu2K94
07WvYt1alwvFQdFR3ka5CH4z28KOPvfDJs73PiIv0AWHRHuUHgLizA8cOcqAVwRF
uBsOwf3TSo3ABDHIRRUmEKRatldDjIp+94HGeXtqywhNVT+KVJmR81/ifzt5U68d
3IfzcWcnL2RMjmwpmzOEyu2eMA6WPTedesoSiiSvEsH/LYMZT+NYiNctkqGDB/dq
rcQ7V/gPfWgQxBXF0mWZfEQJGlX3TZy+MnwSOZ2gnfjZP/rR/3vlqULX9xAlQi4S
T3jwm3GRAD9lDonMTI74mIKuvcF4x7RHY1xXEudg4SCo+MSShJioedKY8Lw/4kIp
1JEhm2GyXQcU7fJjVpE0c8uv/axTAJhPebdZpFSsbcBaCG5EwMe5PbnamjdZ6kp8
dc8x0A2HuWhKltRtM8I1BAxzIdn3NLy6kglUMEeII3ddeVmr+uPQzkSLivef4vH9
wUM/5hV+FR4/L0jI22Y40iV2d4XmCdUcJ6RnSZMF/EcuidSQuGi2+IIqZ5Ssch4V
kQTqMknOG1X3HDyImhcBWFgwRCmLVOaeiHM/rhhThJC8W0fhjQazqfuPFH4HB8Od
/IqD6MERD3lWMyUG0Y7FIYpC9ZJRa1tSt3UZPy/oA9NLGWdb8cTAGSw2CytM1byL
4SWhG+dePnTpqPwTVTf+kSLr2CQlJD88/Nm5j7h7q57PtjaxFkcsqG8IA2u0oaVX
s0qGLn84znhUYbjIoAhTh0K70DzLZ70vPPhjxSl+RtJxnIy6DcC1uZJwA1Hmbbwb
t4uTcOOfEi7Hkij9QneR1/V9cwrfyCK1JHczUFs7LKxkgEkkRBsQnj9JGpBOTLg/
BiD/046r5QES/GGE6vzY/k8NO+7yOXfEeja755XeEqEDo7TN9MKZ5864s0XzyeCV
07JfivJPQG8mQpdvaGCJ+s0l2UOtq64KQjigHlggJe3wqSNRtiek/AD/jm1b9jiJ
iFrlTD/63Cbee/rgcACOy4+XNEz9WfV2ICPsPu6cGW0ot3EfVounY7Hzoij3zCiG
2gxoq1pKD5o5APfhfuSvu6V4WqCmJ4Pb/pMIzShvJpPqfnYHw7tT95SSoBjDOehf
F8AF70BAUmDHQSf5ILseSvfXOGtVL6szTMc9ocWn3ciUqAYk+72TiG/n6IrazjM3
Svn2jGLV68WXgt/Lvxon4+uw13oxIpAek5xRA7ur7SJc2VlIgi5wZ56e+W8kmZ6b
HWtDgaQCEdHlqpfsv4Ov7T9WHdgKcUsnQHv4LLCZwmb9H2An3Utn+FOnvonij2DO
VahdZNeVgs+wRaxOsDgr0ZEEtTugjewTgsjNcg7LNxB3pcHADE+k+gFRtGHkLtWk
aUPFoVWwweMszYE+wD01JXsUPf5Fm0Pahz9570KEZ3EUtCBYdVmvoIc+h7y+FIyN
DTDL6+WxoCe+BSPEzLEEhtSmfsoMnQdUtwInP8yf/BJhMOmadgNskPMqa7bCTeQ/
lUWzV/+NkA95sb076JT+ZSXaX7oEw+gfhrJzN98mFoq3ALdk2VCiXfNqTvDtvjOt
PXLwvhAUgdQYhHsqVYkcIQvp2JjQ6R5DlVzCsyKIKsaa1gyyYHa+M5hCZGNnOhD+
0VBVQVp5W+qXY9DzWkXBFsZL9+x5vHqzwibQZWHkckJM8fWN2VDaAfRsk6xnE8Gz
QpIIZ+Skyp0BkrDZqJ95yCITz+SJJsYfY5mupuDUXb9s9xraiqOAjKmo+rJyhbDM
RnHAiuOeRxftQ98i0G5TT/Lwf8pGk2dfstfqEDqJv3/BGoTwjavJ2U0Ug1QNKC2I
rkNaIQKb/PECmflbdK+DUvU+7nHv/IMOINldgv7jq4s2rQeDCFw5LKgYTx77UYeW
UKjF3Nh/zrk6kpKbIxVKItmynk63/Z/xDCNyQvBYtpuxxLQyjiYkcPn29ZFNLZJ7
PO0aC8bqLhBc96qWKfRGAxZvL3hS1vF+jrhr28xi5mdBAjBwytapfBBBHMlBmzQv
dKiPyDku8Q1zsuwjJUE7EEjHD7XY3+MNoYivAnA/I+3is3qXKtGCQoHUdsDDPs2V
QYBwFDPJYqep+VTvsnOYsttqtVTmRMhscV5xgdHMX30JbmnnAy9NNV/djfrhDlc/
9wE4iwbW1LcQVKNj/4ucu8cAbOgNkkDm/PX8mH3ScdwoQgbSt4iJCuPuhKXPg4ci
/IMxrGt9ZJnbGhGECYB3iKpwEYAOIfsm4iwvbn7pAwlKGkam6ZMoF4FEXZcJPI+Z
X1kNH+9Jju/F3OVlCtDdj04kzrqCU6end/Z3yUUxRdGYE0cgJ6RvNfKSpCXuAUgt
BxZNeBIEsLLC8T9caB25G9mPjSvD5uxK2wrmfnhaglvLNZLWyAvQyLYCJewXSW20
JKc01BgH+0cJmGBgB8hX+z2sYS/s8J1MlhLX1EnZ+uYS5RQ/ca1v7IfgghURzlqe
tqq8YJWi1jqVZV2yiaiZsR7vMkAWRZSXJhUz9v7Fn/CdDLI3cBHtt8gUXtEGd6H2
udtWgbmnUiTe6Q0HcEq2PcJdhKa8x9kevNiUcIVo/5UuzZPUPhn+nWcXqzpeLoXt
de4BVm0EAOHPg07vgk33LZsFzRtdYPM9ZUorI5pzB3hTEm9Y11aJJm9TOuH1YQeT
DvaHY7Ii2EuUoQca8GlDXva9UzZUcWxGgnrSCKVh9CsQLyAlMt32QeBhNy+NqXfb
2E7KJzMZG7cs+ytnUXY7PUdQdkGNhQbox/lC0Xbd/0M5ss3oqXGDyxWpJRXrDA2Q
0V8K9hNZ8ivf+V3tjY9A6GoO45I5i8Qg8nep7IBTSdXJaporX7DLVfipvp/L7Fup
oTE60LPXiwUfLTiMpsZbFmLnoTvglfzcAblzZtCzUSbliUPe3wm9TwnXhEV+Yp14
LHLdAw9rBi/7rntcsHKGWXbVHBMpvVk2iwWmpwSCTI3a/ECW1BbRqTOUJLa4SPin
pLsFj6rCFt6kcl2xU5BSDmay4yYpbqk91StQjDReBbdS2GSQk49Vzi4BwI1vDx6C
0Z0I+6Vx38VgcUBH43ILVoVWHOytJm7MqfED65YhWK3JyvvVsctmJe1IPl9eswKO
HaWkmv2jcFDGl/ZVjZKKf83uvgVxPSg9BU0iXXMkbmsQnJDh4vCyPbPVncqZcRFi
lA3hQIv+14P12WMjjXh7dubZz9+XhAmQVT+YkESncJmFwVEiV12aLe0jOR75KKE7
pfxaeLvJ56E2xIAMZB8htDSdyjQqODOP1wP+C1ANLd3Ms+RbZOOhTiE3akVK6mD2
YghhcyNubSKUfjf0DILwdlB9Dbyt6ZR53UIFVIqhN9A6CirSju0TQecPWcxDiUWq
zpQLQIVx0pCLpczJia2RxAqpVN+5+zuuDzAWFxAyPe92QLmRn6hnOeu/bCT/0n+7
HZUeWSCp+FeU8+xT0OM7CyvPn/7/k9ZjDbSMozmC9hCFdChvsZos6g1vfKxZn/ee
fPuSx4FFnuVgAxVbJS+FJEEKVHwdedqLIyYIS0/JkTH8W/RqmTHpH8IQw/aVyiPE
7sOq11ICDtuqT0u18TA3cyJOrYZ2G0/+WZ24NwNQIQMY5w7EfDsz1u6lrmbU4roX
l/DdiM6IAjJhoVjlsxz6XxhdDOtk1SEo9tFVarmhRcskJtRSq8N2MKNl0MkZa+fw
/z1qYM4JvgYPzH4o2GyMGEjEHoeIZFUoaK9IumBf51psnuTwMqssuJLXwgrJPLRS
cZ92FA9JCQ7PdcuP79EK1dF4pEKvb7Q0mxtWTHPYk9eebg7FJnsDHI/vT5AbXhoN
ImgCYnkpbKHEFysfuTOdYoaUVxA38aJHu85t6yCVd+ADiknZZiHXdcTX8ZSD7PJO
DxMpMGQWXjej6SnDcQjhg1TGDetkZwe/U14sED8QcLAgqL69LIFu/Ckp8TQfy5/9
YN22D4kvf0jbYDcYPxBYGrKjqOvbtHkXsGalI50WKjdJSWiG+8NCPP+etH8Jfufu
6PpshkvbbNRpFt9x0DD7SoRyLtaqR5cS09Fm1x7+aPiXIi4VpOKCd/Yk+tKajuN6
HP/vMhePerFngAY8GLAndm9YJvy63ylCvmgFpg7lHaAdz0Yc5rOgRyWhe+UBZXPa
8lr1GKA5O5kkRJmjQs5i5zwsa2lw2sjIxJmDHIT7/kkfuU3rvm8CgwKmbCifsPLd
LECP8R84Xdyjp45gexY46Jv8+HeBd6R+ktzsHNMIdqTbPx3LS5UZQmcWxayM48WT
R7dr5pH6u5oavHUlywcxc9W7TVITJ+NDn8n8uon6HHapLxGAmLjykAPAys4c7pAM
jqTE8aIVQ/rGSS9YsTgGrWpZ6aDM4zYSIWJnI7TwrcSNQuw7iZa21Vi3Emz+RR5R
ps+rsCyfO1BZ0yPmw8zCABwM7ow6g0DL8adc5V5kBur1Ok3KYNDC7dJvT8LXo2RB
SoCl9TNygmeO3+xdI0IoEEcOxw3kNWCGQkB3dG/9Ktv7oOBwF/Tq9vIleaSvGKw1
a0iEIErTMequ5oLWtsj+E1XztrvhfNBZ08UdkrdrmEgeXa4HFXGiIhigOXqYRYBk
VF11cYtl1isSX9SBHM6hz1JyzQClXeqdieK5UhyDbNX5rGex+Z7eElBEUZ9k39V8
1tdRPoww2GZVeC1C7SKK4bxAl1rVsW/ghimHB9Gd7uX4IYrobw8rxtINl54XAsN1
d8bZXKT7rFekJ078dc7K18u52+gNdmVxNzDy7g/LUWqKwkj4Nq5p2HSqwgRubi5B
d5G+fDQR6Maqiu5NtZyP82uZmcv6/t5vWflBNm5NDxjYgqv12GY5JcL7aqio64vh
oOe+tcz4Z+6h7Sx6+yWQMoaUZQS7Xnf1hhqGaQeC5HunYf8lkVIRByvhO1q3sEQz
4Ky7b7R8j6nTmvSrJ2LCPorIKVk29nD12/JbiaLTCcReoOzqtMtLMRNlJiaLSvID
2G8ILgYTgcj6DgDVGH/MToWJ3JAGMlBAFvpZwGB6JRmeEU+JYuY89qeFNpLV5RrD
J8zcI3jKhQp4w8kTie9UycTlQKPScEVmxv4pah5cVQFQcGu9nYHCiKuV6oYOgMOQ
Y1xD7mCZyLFH/+5fJFGGaIpvFtNMZrXEAAk3cJ61jAyHVsuB0L08S4u6kLF1haAH
lLEmTm1jSpiK13rsh/QlvxXuhyPZOYVVcnDaNxdCjmNnGW9soYAgHCUjxPYf5mwQ
grMtqCn941EjR60q1Gy5KlWpq5OQ+yqI484FtTw9mewix/6SJKEPVTFhlntJt5e9
fhTiBqvavKm2+zlnBEVL48WRfmvADWKY3tbMIVcYeLxYMPxc1yv+ke8EXNHZA9Je
TRr0spjgMhIZcMMrGZzDq+/MZTxhFqmGH/1IGx1GCPe5xhJHa50CiB3QvllrMpvD
gB3pVcxRix0jBRKxtbLbPXTzZE6DoLiwJg0Oh4pq+J6Oz5ak8DfPAXzShgMsvkAU
1aIDq2vK/6FqMO5Z/sMjxsjviciPQwTiv/ezlI7+qrWeqTWfWtil69Ffb1BnXgpL
WaLWSf5MM6qclBiOfKEQ3538GD5yzjqiLnwAzoHGyuDfMweC085DMUt+jKFhIpLv
r9wYwEXSifcA/y+AegI7jyDPtKZ27dWJGjuRiNw7IOoqcc9Dnx2OUAPASpk5WA7j
H88/odUOjeF5cY9EiWn6b0z9AHyKv8E26Gbx5m/4hvtLkNI2SN6KtpYZ8b0Wfhaa
dym4vI+A8c//TY6AkGHZYkSZBVLP/xz5FUv1YOjywCGgTWoTcwxLlvCLBLITy7JK
P7wXgrt10cWE1keOTOKc3q0HBWSadnjK/Uvp1XivOtsf937raBzhIewdrxb+cliq
9zjfG3zcSbfdpZ3YL/lBGlGoeKzg1jj6knRw/9UNpd3OalnyOTOF6KWdem/SYrVj
7J6DYK4LAlngt9pX1W6SD7P7K+b/TuJg1r99jrUUK6i1yqi9xYs1zA9xrpRsA6dI
cAnAZQ1vx44NNPFxe5G/77s5rMFWGkyZEi9eeCVGoSfzgrzcZu1QxgGWHqyMAJcT
yWBIhcnQl6GKkwSTKGhYPmIcB7oYGGA8fuiGzLA6Qz0owA9GGndHNbFxYXbjEOOt
ZbQIeWyDnXbxEX6ySlO6Xd+jdEy46pcDUni2M+DFQ/Sk6d8BZDF2MECT1x4RcC8H
l992h48QJhWmJGLHBdDnwyQnQUKY7t5qrcB5tDYQO3Nm1Bn+2GtgIgmVwgcgUJUQ
2P/bRLdCbbRlUDMuJ7UJOfa+TD/a0V+pzicKSbkIIAZH/xkO74I0WiJ5ZEvV7wdo
jH3AOGEQb0A8EloC51yGsWdwpwoUkPuGRn3P7fDXhHeyJ2LFFo7NUsRCkwY1cGvI
2Bq4AX4rUPL03FcZ2PAnoCE7cEPfmv1Trx9rmFyT5W5EKKUqxCgoaWUJzAsZHW50
N555wiotYzj/fUfbm98/mhQChFJkMTrC4kVdGUvYtO+MuYSUl2s14gikQYPCghwn
aHJYmYiPjSJnut2Z83FBQca9afIogPqu89l6IBekVCMaXKks5Kwt2HlFCpL9UxbI
83eUj36VIyao5cBN9OZfX5hqKjP39EyxBQwuQlOqLLvubduxk2vJA1+P59Y5PFe8
4H50HSgOOGFbnU7VHORQgkJvv/LugWjnDcLGi8N0bn2OABJMpD4lFQTo2ez1ER6p
w8tMhb7mBrZukR27ArKvi5OBnu/aWfnQMAvCYBUFPjvkyfgfYr3lQytQcbUccfg+
r7wdFrnhs5u8tw972ti2XZ8xEXn4IQkC0/veCUUT+x+U/s3WRkUSxDiyL1SEetUj
WDur/keqDLmqh5KX3uSkHlFJOa3NAHE2Sc+l8FFXyZUgsPa7XLmBJ9GxI+kZnuF5
fXONZ8mUyKPpSE9JT2APqilZxD3TwEJQrex3W1DYJcBRyJugc3HxxHbXXIZEGz5H
DEE0pTbgggJgJsPxKzaa/YkKL7qqGjNt6JorYGydCnsdx5VDX55Oni69sTH2SGDq
358bRPvAP6NhRzQmR9zm/ppK0ALHY+rCGo8HU7xxaqthvYC3MmgneYmUxCgUsNn1
aQ0X0GGB1O8UXFW5q/wTSmR55OwD7Th1ey3JCZ+ie+92SapH/aKHYEYGtQSi5hFa
w3vcE53k8ZO6RFkLQqMeCwUGLnHl63Es0fx4R9a34KoU15ZtgsaBdcnFayPJkNky
Ex5/9kIO9LSXxFNH0kTNhpSTSyFmvGwp6eZtp9zchT+EuwPRtsKqCSCh0yzI9h9t
OETKxBQL+spDjOv0am4RKsroFzR2Jc4dPY2sT0+zSr7Dgx/N5txO9IMgsV8gDfCt
FKjnGFONWVIwlzZ90O1zaaxqHEFRa0J4i+qd0Kal8+BuAa5y4LbmzfWrsmLJlX5H
7A2UOh8b5vs+E9Xkm13BBuJJfjJPMTkds7WJcIrcKM1VpNuyBpPji+qnG8uRMj9n
i9oftocGSCuYRm7otPu+U7WeLYdxma3NWvVoHq6t2KSxp1YHmXeMJEY+7xEyJhPt
XGQ/7mnKI/LHti9rws3a4sg4ITKHVKC73yRZYuge6SXiDcGSekxEKfdC9GuoZrh0
KZySBcOCzOov+GKqRfntfnc9dfap8n7GcbEDLoDZe86HTExFEci5gaF654ZsS6xJ
2jaTWOnvN+tIoITAuPd9Cke/Zudt0mgU6ieO2jepDGptLTggHOhiuNll1uoQ3XIl
mqW1XzCafhQBLnoFTLsmcmeK8GqEpJhJW9jEfrhbZAvSkCmdyRP0sDX5EpHnT35x
X6zMKYB1Z5lwQuoMk5ueUSpo3c+CS1MiBElNr4le7SplUTK9eBeUivPETwrGqU7J
E7xhBIFuIhbugLIqOXKnRQy9Mt0J9viEzuV1TyJY7mk=
`pragma protect end_protected
