// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:07 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rd7tijiqYdyiFPYMNBQ5DMd7SzRoxCLidTwF+TtXBooQKTWAG3IAcn7e6GLZsC+v
5tG+9fthZ5tKNVfaOJO0wLwuA1o0O3kw25C1vZqN/OauP3h+/9X//6Q4xca7C0Sc
lug7xKRzELADEdAlxUSpyxUa/8fR2mIjOmrF0O71dZo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46928)
mElXGqeZYu0j3zjGQMbO+HxuM7x/1lhLX0p7wXuSUnlPiP13OmyT2d1FBI8x1jwP
Wh61DVa2nua10epKwvMYcIqWR245JOl6IZORs0cPufcmmcNlm/qYGkKblaRqVTA8
M93BeTkGCgswkvQI9XuJpQhO2LjJzAPo1UGPwI7iD1AmmLWIL5l3y1M2fB8VWjc+
a1YYhSW3Hpe3Ywh0JZU+AQBTSHACaBluvbimCJoKLiQ8qypyHdzFzbM48C4+//DO
l51yilahkrjYo8lnkGtGRIEsdQQ1Kdw0MdLLZlsiA5WhbzPPp0LEJZtgcY4Aus5T
MwRCCRvcRsg+7g5sIFd+OYCzHMsbXZ+0GcjXQH+S1WaVEVIizDDPFuy4n/fEGLI3
S6gJsQThSUU1AeOk1lhAzbt71LY3W3BnBcJ33qUCg1Lorr06eTVBcoqrr1w5sE7B
hchbLCV0alNEqR7dAkuIx68YunPUb1paXXJL/deMgVBy97ebEZI65BN3lXwE8rS0
11i2AVdKeE6N6EUyOYXyl9l4I6BHrBMrKGVZoITTqUpbgE63hqmHVghQwGAjJl0+
uoQADhc5hdTzDsic/GDkhcOgQquq1/aqJug17vX0LOCzpymuBrZN2p45PHl8yK3r
bwtn/vtkuHnUYaeYNMTUwBUhHc3cIrQnTx2cbaIiIh/nndKujNPTHe+vBu2KnSVG
fJZ1y/1udHpa/IDCE4+IoL/MVQkKvS8DKAm8IkX9/dlpBnsjT/3xrVS/o8pE5NpJ
TgjmjRRvIdVi1l6OO63l85PLw7KPfJnH21S7SlQhqEB5jO7a9SnZZ98I/vqI5kCF
sg2+PigBLT5qWMnuuOFEKYxt/GwCBYnIgrXwDHDhOfUE9RPeiqxS1X5knl1aIb7v
CGtCEbSesU/JZBFtPDNWgTtbfQo7U2QmiUFzJGB3mMqfnsp53X3R307snVJO0H7D
H8LZ1f/ZU+FTz3uaI0kM1ZXrBLnkgARl6FCP1EvxkRYmgyipT8QsArW+lEvCLYsV
tbe/z+kFfDZliHerUulv9qbEMVp55yrdd+0cz3Us8m5IvjkX9XH8waZsx/gjZPe4
+9ZD5iHH37WXv+duYp/dHAx8A8YLXGH2CoZBuKLN0+r9odE9hIVhFHOO09qkElUs
2PGvu7e0LHKrgG7DQ17hH3zbcyCVdZLBnupEzP03hTl2uQu16dkMjWvqMrePXo7Z
Tdl31tAI6lG444yU2oO0TgrsnLod9sG8JDBDF9yF2Uk0kP2hjz0M+yetaZYPsKAD
U2dHESmOZuEE4HWxRAM13OvV33Tr+HsQgEOLVmUbiJXyk1fG4IuH8D5AbrrPieYe
AElxUQr3OHFljRxrcrv4sqGGkUO1TA+N6flOwJvQp4Te832jmYECaKB5nPeGZA4g
kjJy3/jYeJNWyfox8w26oWP6aUrWdruO4kaYoio9TWafBw2tKmNIkgsI5QAddsDi
UkvKpCEFRuwZqqtQttaLkretAlFjmhyNq67qb0s7qb1RVS/BQG7XqTR9aCtTYb61
Lf6cCUnANiG26gylCscqXgLcm7ssFtfK3tkeHUIEWoLWvsHGWw2SrsYj7saCi/qg
vpHzXuxahm/aMnPC/k4QnLhBTMcjk2QqWPvAT2qoMA2d8aB5Y7yl4WBtESUU2F/I
A4yM/VrQ4iRVPwc0uZZUz9ji69BpLZk8ivivcv57Ti49gXl02Ra/UtI5iUhQ1w9j
okkMKsJRvdd7jepjnNqFu9bb8A6i8dX9FXmUTh5KnmRYPr3/kg5ha3efdR4cGgKx
2SPTHm40PlylEYij5CkD6ZuSTzJJd1+viohWUZjHNNtFggw+GuQM+9i3zxVg9MOX
hmRbSApgh06aHvLjWQY5LpQdep/CUzY3NVDm534DE6NGo/4UCY//0YkPMmDoplfr
ZZc6WW3gky3SGvE+NE5T40VEuBRCMe4IAiCEvyCgX9HD49vfYQM2l0lhl2N9oSPM
fjJSYJ9rWMu/pezdJh7hGGXxGQqpFUXsYDr8dMpVGOihOK2UDuuUxH2sL2oxMY8E
8pzPZmnDTQdolE350inMTM6t/x9k5iab49ixFTeQwqjhjF7oU8ANjLuu3Ht0PYSG
1Ya8BNFPhoejGZToENQMNfgi4d1HkGAibygeWGwWZrGvkYImTeOTfIR0S0OxOw44
kxBbYnTHkKqPGZI0/Yj521myJhvwbzJnXohvoTmhLU7YiW+1b0x1lHRsAoB5QVUB
XNPXLMo3X5E5Lcpp/NGEiDwplUMq04+UyLjYuaz0JbrAyqlWpAe6UbR9AN8wDnTj
s2Z9ODEAzQlUSgUJ+w3GNyJH5FFwiI7181xZ84wxfvGmfg7DL3nmg6x+ciyr4XKU
DDAgYq/myaHg2kll1T50/dUWZfWYzSKOAFAOnTdL3DgQEV7uNC1bZFSBwCpzmcCW
KE9X/8x2cO59XVLsfciy/MCP23dEI+rWLHTfzVXaHCvW0EjHGadOE+qP1MqidgZB
EkSrtXqYfueTp1b//j6MPIFDURTrnJlQyM5HGFZWPuiul36Vk1ZCJjPTOwizEBk8
peOu8HX81/amDyTkUN/zMlolgQyGiFf/5HoNWYD/mI/QfP9w61KAr+5Llg9kp8Xv
ZmTnxddLD8M59Hg0ytKHL2tYsMto4E/EnwPvNZazygcefX704C0DBk6vHe63h+MU
qToQHszshjU5vmcElau/BnbfpiEu955M3BHPEPUFBoPcO3uuWZduQZI+4yX5Wnv9
B4XhhUxuRuXi5yaqbcuFGBKIcO648O6Ex9DKCzjtIBwqfP4vzOuoJEcT9HuGXdsq
saU2jajqJ7gmNlvy6UBCKXBM4+Ij825rZcUWSNb3vydMTTw6fwe4u2TTDK3VCrbQ
Rrw5HGiR66JNH7aI6QL52YEf5f6GcSpgdMwGqs4tKipvU21p6+m3NLUlEjObmOMm
5WqMNsPbgP8CAETHsWsxRQE8mN5nHm6v/LPqGoa09NGalNP5srxIbqDkh5z8fMEM
bQEaPYL3godIflt+6NRLASTBgijxVUgw92VzY81NVwuUgDhqU5OViNP9OskkliGQ
8hcGClJcxe7UwZQPcC0w0oL9SDKEsm1r8QmaP3yuChAHyY/+cQxKibes8Oma9uYc
DJrOiFeMBjqC5WFIo2lL5dhV6w8viO2kEH8yGAtWe4/tLN3o46MTuReHRj5aMfJX
97yqDzxsKdC9crbgEJGROuI6ZAiqa4tvkvfUT+4u/HnGL478WBIpv7diIhzoQqSE
BkyUMrWKAMWUwktoJzE1Hnw0Tkabugc+eaV0SlraJL7fTr6y0nrY8C5PlQO2qwlY
OG5czVsdy2jtpxll6w4PC84NHwO6duP7deMNSzal+YctmLu9rxHNuesz8eC9ZHfb
7NDgjgcxD5iNTNe0B3ZuP1lnIu70T2p3Hp4UGFUoq1t8lrf1rGdJ/bbt69yL/Z+s
5edlftqjMAY2V2y7wH5fZS34bqvEE9hlUFv4vm7P7yTaBv21gt3W6D8BURXv7B7W
ux0aKSll0Nv+Xn1PUZu6j1+twnRsuYCEEeU+fZn4kHf57kx1lW1wq+q+/u+MyVG4
qrBTBv7EBAhLsIeBwLb60L+BCscEfZMYjxFT/7auRAo2JxfDOQqX2CuOnuPm9w1+
rHxZVxqpvT8WuuvSbP6zZ8L7BvhXq8mrdyQMHQl1txclJS1lYKYv2tgVYoS+T6oN
Q/SFOMvGl7FKoMfbNyZiZrTc41M8q2wwaG+Zr8Ddz9vaQkvHtu1bCIwC4IcYkYsa
YSh8XCGZfqqDTD7vU4DJXXiaeugb0gDEV763V4XGsVhq8jc3zBUQkFVsvyNUzExs
FHx6umcVpzKR3w9ikeYJuvlpryoCF5KO1LVz9BLQXbYkqu+MAgyt+3l8VPBSnVC5
E61u0RVQJEV9XoHb0iPCkdCyBSyvljekDvtId1exEV9F5ig34kGrKWcPBfpTxkQJ
Mu/We7qqDzPR5LBxE+SiJVpXlLft+m4e77SfcYLUZpVlhCQozn9bK7STuWE3Nof0
uqeQ00S6+eSGFVuliufZnk2XUFvdvuupdkVPmzo7deTtdyAU42N14jRNxiFIIgSt
c+7pjPp6t3cGo1CsMWYPyfzXE/XQfI2Rlu/4dtEYYFIQMAFP0g0OSvTEy7kw7jM8
lA5fn/kTX8XdEhBSqMTaMKYca6PKOdgZmRPFPZTRmBLa7enFfO1uraW7+6Ztu1qf
lp6baYt+Xkjr4IQTghx0rBTzYFPHH9XKDxg87DtTb26/zAHlYwtyshVKOMVnQr7K
Wuo35Ho89yYV4gqPy9NrBGmzVsHuF1r/m8FOOZrv3gVNadQqQh7YJEhVAozQSPYt
DQrCR6vBxspPqIK7aX952Lf42ajOId9TPzOkJxqtzLXzuJvN8CkV6gRXD3omkvO+
sbHTdPw/wgn7idpc6tWH7+q1lpcNE5xHUpUF2Fn7p5bGPvfqnK8kdJiKViggW8Pa
bRaZjGWEA36MfduA9mWl0AKdyHy5JjNKEoTpyGeWyir7kU11gMxOD84hhXj6tMWO
fSNwupfebVRqX1aRuanzLoyEEji3BVoqh722WXTLrZ8CAtbmOn6j2FeyN5MmPxyW
esaReHSAzxDKs+kVo7QBCRzPy9Sc1TEWKEmnHlKWBAXX+enBKyly+HOt88vlN2DZ
1+DhLQMh8gVOSVdRCH8iDSIH/p/ysPDCEi7N3mGEPqbpg2Bqou26nc8CcmTXzKlI
FyZcaKC+NjTR3Kx+Sbyj55p7+OnH2yikpU8Fchkt5W2bpkrEPi9tozQW/u0y0NFX
ELIHkqOlsppYs3JddY3vMFUTpCQyDqejtfb9THsqJYdVixjONDkvILJ0RSWaYZHl
wjXbMN9R7iPMkbExWcLQ4fL51zDSLU/9llqOMKUPCGlGuuraoYOydCCqQKqw3eWv
23uEGGKj3AOKMNWPN8mwjXpkNBoYVLJKFuDa858J+UTsUa8m6JWxXGwYxsDQJS9P
1C0NzWkC2HLLj9MUat1H8ZwGPkJIenMxcPqGAbGDdQZahYA4DrSx7IFKcUNnq30G
U9yTfoC0DYxKI4oIqikiowCfcJd42beOoYIWdZelht8VfzCUTVsA740D22BGnk4P
GYTULKMeBBmg1FpKjJO2SL0i4QA59AwPZfJVFHcns2lQxdJnza5KmwKgFi/Pf7+V
S3QVhS9WXEbjVqTvNfudtZootK2zWLoqmfxSiZ4YtXxEq+sSuoe0gwmg2t0AEydb
KCPkBfRCDFVyWZXR5cKdWCElzhbH60XXvlUheIDZwGDNy78UVUQmTPVjS4QbR3Pb
/tQZSAFDUAZHY30rCA7+ZDulGE3uqzT9C7StkfnkEuZbEzZeRKIf+M1baSNavj9/
ZLoKt13w35himjx1yvLeFHGricxqVaf/H99Z412sxsr93RKvXwmz6l57IFkRsjcI
OWmC6xISReHpyUYGVrSgH3hDyj5HaMbfJWrpBMvPEligjmmhioD60fj2CS4u/Kj/
xUOAOrq1z3rPXzo2aR8hwH4cGHwPQEyqtpKtSbmAMWIQ4UvKPh99W2OzvujQnEEq
HPW/YyBWeytSEbzOWRQruLg5voeEuBvW09xUo38/1LWbYFQbX3vfjSBqqj4yJMjC
HVAJJs424HRkqvI6bzMUgI6V5Qqgw5SD1BBzI2JBH3IFdeJNqLbmJ9VxvomqHn6N
ocQzCUjsx7goYtm4ezKeczdwwLS8Ke/HWklBs9v1wO1CWJAW5sKOs5z5YZhYtZjb
0qJcMlEQ1iJCc5FFo3nglWxc62tqd7zqUgVlqZTbWQwhgSdiZ0U1Bv/14eSAG0HQ
wFrYMrhD4rgI98rPH2oIleot7mXxgZBNcorubap7NPuzOAwHH53NGzTZeI5DnS6L
Le1vkGIebHjMG/83RnATG7Z3F1SkxMuC+pYYXJLG/UbDtusXBZYC6leFJKWitiaf
duOkOHIk42gW4W/UVWSYP/TH3jOLTZ7TU3aEnek3p4CcAQP4nN8TlKwCjSv8Kbq7
iQVoHjwVCrMKc22TipXDbWAQmtHvWpsON5auRDXSgRAsPkBSfJPhJxdkSzBk1AJ3
25ezEJiFup4Vm0MUGw4XDeg8IjbR4Zm9kGnQgUeuizvdJZi52L2cd1RcvCby//1r
vwca50Z+HrxmqpTCdSt3nXMs/B0mdjVmSkZfsh8guKBKsLgxPaPYWhFqLA3laD13
7A4XkEkq3lJeKmzWXNU/PNwJLwty+uSWIBg7oTf0FuyRg0pTyD3fiE6xdmO8G/Wa
Okkb+7+mjpoW/892VuCQcFTmeyeDQfmXtS3riAKcnsULsRXvidMlmdy34FH9YbPZ
cwbGh9OywU9NhUVR5zxrYklt2Sjazv7nFQEIYDP3ItjQXCOHslT0zenTOJQ2bXIF
WhGcDAkZVsUsMtoNnlubIsW+JhTC1q7WUO5KuuzLCnFdzJzugvkxtOcw5HiP++fk
HRptbxuiqR/txhpqdXyM2IXiE5QWhCwayL5m9y4iENRt/Rq8o2a2/cSxv3AozJ1k
sLEAIBr8vNALYCeo3QiHvIwLPN0ScaVHJ/63aaDfBAgmjzZFr4g45pdS1hILH04F
WKE66zmFrt1J5xRIvqjCRzzzOXCWjpcqsq/yVpw9P9EMgurPnrXDKNskyh4YMyxf
arFuL+VjkzJI4/CJCK6S2JZ7q2sutYi3ILuRiSqtEqp+kjLD8f2c9fzG/0zsG+aY
WZj/7jR4k2027TbTUkQogbLheBm/HQKN5fZNwpghlI/6CeabKC00UiDz1slu7EoL
h8Szr2I64YSrLcrEZnEosMbyc+bgWsFBVe01/7D0LP/VTw760zOdd54ZpPVoi38X
Gugr8lyteuEtsAmQyBAsfom9/fQNLuwOxuuen14zY9TY23Ak4JDgxPDLRQKz8Fre
Bq5dvyFuANGQA5msOtowgzJgiEBaEgWG7XkZ65xMHw3MQO7u13VoaqIOAXhzGp6d
I96XIAWflxgw8/kcYFqg0xV/+ZkUtbkCWSCF71RkC21D69tKpKltimj8M0Enk7fc
cXaWGL5t/75ILN71T8C9h05RyLAI+mWC6tfjq54MTkfgr/YZNgBXlgfPIdeZhpVt
iJ5spgXcmOY2j0g0EA4o+p/41/4vjQuCHLMKQpBM9dQWEcXmvMxTL/FfCL462P7B
Zo5jfr81hx36BkAmVfLrUmXbkqlDqfxMolIT81GzRjW4qiUbXBGZrtUXLdT2lPCr
IlUwUj45ISRLJO1ndJapnYzLImnbs3hozYte1L6vsPWOV6fLzCUcZTDQU9Szs3UU
SNuhFVzOlU7+/k6VNOTBXTCi5N0noVBEFHhOFN5O7F4u8qBeCxEzgw0N2Vls651Z
x3KYhicHATJq5sE54MmZcdTbRqXyZkRaABu29d9oEgKnHjpayFzc7NJX8Uwj305z
estgNBUJxLCmE1jGeGDia1IvAXUuZbQIWiropnM2H9V/gXfKUuS2vv6EOYbsLjwH
4FCvfRoqg2YmKY1lFxKPuq7oBmCb4VR3Lo0iQSEjNOg77UpTSJJTPGgaPw5hGAh5
5JH5u70ALeH580qeFz9avHrLNec7RLoOjrA7jHPNJ9F/3jSW3MFOelb6IX9jqSIt
uNd6mG486F4YaCriwI5SndAxcnrdiQx5Zyf7vp98KsAMDTez0JYwPTRq4US9T/fW
81zb2r96Djr4ft8rwmkqqhthIiMC5rlB2rI7lQwl3exfcbGAK10ocJs/ajfA+GqE
tQlY7JIZLR0J+zo9ddEov8tbN5BKYTKejro0EhLM1sU5STTRVOeNG9zRMylTgfMk
w/okCxYM6i47MVUTvD1Qo4sMhgmsUfubgn7QtgNaA4Ye5wdyKNUhAQTH+2HnEyNv
BibJ9h26TfafTUrUr6xsMl5T1qypnhMdN3E9HdQ0nQR8WoWIJ9zGsve+j0VRO2eF
/zpr92POq8z5Zo3MIeA7DaCxdI41hYEYMoqJHm+fuiCYRPrJ1o9bFo2jonvbZ0YV
K1igHZ1RUNns9fadxFHn6SkwwuXWt50ng9pYt630VV+pqkRXpV3hB285bGfyqHZt
Qh5YW0bMfHeGexT9WZZ7riGugrvSZ/ZrHg4j/ESWKlTwLt6A+JgyhanNARs92Ye1
UGRRIWKgELH6tU2mh1BqC/sa+2m7Ucrnh0MIPO5V5HOJqWdH7TgtGZS88KMU79X0
7qDcUGFFG8zFyjwE1AO+SEE3jiPIkMPoFHkKO7/gtUuCB/TmWNLYRzOO9MY3CL6c
BscfINazzAs+OEy5T4J0nCrtx1ppJVC2QwMGBYaMtLEl4AGq2CoMATIkfZ1YxLd1
RvTttr2WFKLPsVTlMnmDnYMj6eD8OFURjoAuJiGiM89CYdUwsT66iEkVbQlSnBaq
BvrLwy5J7LFIVMLPvC1hlEnhoO/N79P7Hzkh/2B9X5W5xL974zxT8heG4bPbFt4c
ghD9Wn/YVi6zC3ivfTiouszgjr4Z+NxlhYvhBCfzJqqzsWVlD1CcyJaZfoMmuKuq
tAATLL6gqyzMWGz4qZB1IQAwppiuvhHDbgpvtI1pkUfYy/bsSbXVd83YhPdWlw8v
QBiMRuK3j3o+n6IN4Yqr4/xNc02dPHCrti9HWwmlodSw5vDgD1xcstDCvJ/aT+KI
TpBdAqrxLnu2KO1FCdz0ubJamrSa1HfnyUaRXWSDFPFu/9ebwR+ZKH84HdfQN29x
glIF9KTfoLnjNCGfFWjWQxWp8st3DYRtKYEhVCgtY6FlHfdcKzYXtbZTOLT4Zpur
+l4ymQ6h4VYsnJjiM2FpsbF8kvuOEUmSgzrw4TuL0PPr5oTyoEWGJkd615fntgYC
Yc4TAaqqfJldexmRLnALwVCcsJYEHJzQ7wDPmVxDB6MlZhckZ0nMC3gzVvPAPzif
WmNMR27aUNpBsWtEUeJOSHn695pVdH9zDNZQJ3I+uu8KgY9GJWN++sRYDbeLrNyR
2Sp8mTdPR+LeO3L2PXbzxTQjQGZr/eU4nI2USowr+SnS8yDmD8XHJ8NtqfRzsjKQ
PkyF32j3MgDFY0z14nvCq0TCF+sHC5kHFJfDmOfx250mH3J84BUvVHQBbphcNRtf
WFzZOcvQ1OjZAWxMDdmn7TlBEeEMsN3zvCVlV8Td55gznZ6mTCrC+MiEsKLtrItv
bAW6XoVQ99bkWM9Q1WCTZE3tlhUcRN5g9XtbTA6QCYSlyhNOu7FSnHWZGrbk1Isa
ZMzYNm09as7V65F82FvcBkm31z7tie656HmebqLvictHHD1MqudYw6CYAKu0Phe1
ldfo18rgzpd7/l5xpL+D5gJIUQbXej9c2D1QChCokKjt72Aq6DUYR6haLuzsqf0c
N9rzgjHmvgQBVOBNBar3Fz4AaoFcD4oGg9dJSe7t97LsbXcKQSE3Vqn8+3eRcT3i
otXi3fABv54Um4MCS3kCdTYfXqVh7S9KlZ7KNjWqklxu/SQWGLrk9bAKhdfSSvVC
jcNe4XK9sqiC+Wb9Aih+C6NSNOPFOfuN8zJNVwwYlL8fLvFoohGLa88zqZhDuVrh
wuv/6ft1e04eyQcfL0pIZlDlqq/PXlfDjYjLzZeBMQymSJcDbmqMrsDrUQQO+pDt
rhuuTyqXE27ZBM7Spf4Et0x44AO710s8Et/trwj3lVwiUBrOcaO63/hYV5geVjRd
v06AeO1fOmyr1DvnmHcyciDkme/Bqg3TFlKV5LnVkalB40dZL4wuiawvJDReh1qU
5uqNx+srgxUwXWdHgPvpBcJqaBL46D6yx/UHlHUKw9TvExYi3Y8UUWfTXrFO7uUb
dZiFBtBLvnHY7/Wpw6pY5aYr/89OCWY/u4VvcAVeGEHqXTIrCWxm6h/13lHAAmtc
IP0qHnuamjAeJHLjgB0V6vnCDOkurOM4n6oBws7NZEUD/MLkEs7PQDoz+NPdvziF
/Mt7FZm9//WWOi2VCzbEh64uYzrzkEbQBosGHjnKXXlP6BtyLrwHuveGGD4xWQ5u
gILmmjkuGR/GeN8O24rMn2/jMBvzt+lLqrZI0oHbHthotO83VyJ1hCtpBC3ijtSb
OItvAib6dSo0kZAnV/zpf/KEbLoawnssbbYS/ZWz7/c+JctD7k4YYnpGcjwVHfkK
byU6RkgRkMZcpzSgJyMc/ai/CSd9CzUTHpcZflpm14yE6Qbe0/RcNCm7BpWmBvAb
J5hRGLL8NHCKy8ST81TNWevfczzqeb/9RzUpwlse5aNIZou3bNntTDIQFfQ+brCE
xuuinp4kIYp/EFFGxT9EaGYX+ttV2r8Bx5bveyDwnw5L5qWZVjds1nZJbR6TjGgl
w7B7s5i+p+ViAdY49G1E2ENXwsAYLtCRICNSMkS1bEbnYY2mcocBVUJ9VoRcrAad
SBSMaK/VvGs0BuQ+IDhwc+JftWPGqq86dkxpXZnSBdd+0a1qcP7PipNLt7PRoEK4
G5z68tJKa8WghCasU/h3a4jqtP64Od2Oe+y1H2NPHJ+pOGeDNQ78tQZEqBD5/a7I
md0ZqTDMXxnn/1kxcFl/eY3RCTveUZnDHx5xhBBKIwLkIBqiASXWen6qfPOnPOYr
7KFTltHko1Vy+W0Lmf8fT5l9h5TpFvlnlsV1U7auKATlaFzUToORDU7Saw+1k/MS
yCnsrUKbAuz4DNb86h3jTbhwXzS6w8y9Gx3QCp5S4HApimsEORSzbGWg6jUaN8Y3
rUKjdfaG4rcCnVIvconCedoMrpB/J4zntRk/2dyNw3RPDqxuLrfoDqRHOTtSVLP2
qqhtsmrQnJpwtAFA4gVgxj5ItLhEH7prFBxJ3m2InnnaAHn3Xx4hNm8Ob7xPnq+b
NUtU+8QYvZNAHe5Qx2xeXwjx1lPi5KXb6IcxpPifSNB2LtTZFhRoT5wyfLJjK+fN
FIONZgusSyFW/dpLq5S9yrZecARQ4zWcfTTJ+IOQOLmttE0Krpr6WFmMWgM6VxSX
XFoQkSxHP77Eu/9QJKu+EA2EVQNXs2P6Yw+2USNMoRHs504vymyzvMCzh7HkkB3S
sbB9Z3UBUMGyyvrQmTET3WhDGdHUXwh6zF4DrOicChhXiUXp24P09mwsNA7BxEQ0
UZ8Q0tBQcXem3LoDAaYD8JO5aHw/zGaZeWbOszXHs4u9hVC5yGdvUCD4YWR6Gxzm
X/HDjWlnZmRmt8Q7L6dh/CvAhY/PuptyKmF9+BoKHVwof9euK65dNxeIHBCF+p9l
uaUGzQcs8khE98L12a/Z6jp4V3KxWl8Bv9Ii3RuW/I9+WJEE/Ic1xxlj5+L8djx0
a4x+Hl5r7sUme0DyOEGcivvzMhHz2Fy9SpI4ayBfo/nQHVOp1i4B1OF0GWLFzUZ/
sFE2mc6RGg+IKbp+H9y241vKahHnOcGaddaAyJ1AZPfnJwiLNLtfbBp+DihwdEaR
aYhMtzD/l7RiFzlP4IAvQ8Zk5zQpYdl/3pjKhX0xcbIUX3D+yBMpO2zCQSF5Ho0n
xjPq82vXJ9FMwrXRh+EsCfYNEbeKp79V1f3prAA3lRAP34xYz41aVofbXMH1c0Un
C99C0cEOcw993eoUi8eATr7gs0QJwfx4WzDuwOj6LSyIud0NVBxiHGvmj/kvVUAr
JZq66s2n/t0wTAcFNqHV2Up0ZrK1pFgY2eWkzdYR/rOywxySyGpqYoN3rBSD5mxW
Mm18l7oa2mPEheunpw8g8LJea8LOJxX9vWjEVLu8xLTnGmOVxLuKJGCCEHpj4WGK
bsufdvC4gyMLqK6+dPUvRIvETSATGOCHqU22pRB5LjYWJta4kxA1LBmrSwSFzgc4
18ueAv3JkG6aVyZmWXqZNcBV1ZLWgQ7Jrwxv+iIFkaaWUxUG224l0HFsd4SeK1im
KgeUEA+BgkTV61LOzIlfY6Np+fVzBSYSjk1hffj2+wxw0SSjQFFCVAxlKzQs0D5q
TAaRyK0PVKm+X41Zg3P9n2pxc/P7zQT6sJN6Wn71+LZW420Lbyn0OW+gG1zR/N99
p7VR2yuF2FKfFoQ/qrMm1Mmq8Sf2Ce/Gij1RBs3IYzz6Z30Rv2lbXgw2Bx0Ozzcg
g/smP/ZlNZGSAous7bwUWbRYwGF44GDAGpPNJ/CI1+59N/hX1wXhvtQus6GTjJzs
EtdlcIBdBza0ixO4KTV03J1vbe1iRVtXmM4zatRVzZn9Urh25rDgpKKbGUthfQmD
qzuob6uvmf5zxCT0/PzUBPkwqejPgWYcK6vb69POXDnSOm+I84dCr5wk0YWGitfv
eb7ln+EjGO1He1tnFGWxpqpt7zipOU6vJz1wW7Ec9d3ZMqywa9yux+CGmsvMVAn7
uKXv/DgvUVdajXGUdRPUHXEiBYjzXDEuYJmwjo3SOnoMdkE6qLRwFJvt2/mUDhix
/J+8Wbpc9Vft/N+6U17i+WXJEC0/+VpyRssKqvwi2+s2Gpq83StwGh3RmjQBiau5
58cBixcxUzxghtqGk/91pwYIUF7b8Mq12NyQY8VEJAvbiv1Ddk5KMHPcRLcicOId
OaKcJFBpB4B60Imr3aMvWxasVgHGFl8zWrZM9IPHckEEFKxSf2Y80W7BfOxIdRuO
U1CTOT8teRdGgBTFMZzn4KHuyb/h+R5xtVe4OSTYKdFI7Zy31AcnA0AvlJyUQqsV
F1rA1dZgIuwJ5N+J4pOieZ1qvdHm9/1JfWTIXYMLha6lGmHlvywKWtOw4nAMtYLw
mHkBRvRLqVrjeis6bcrzXEUo4xdHfatdgCwQVB1gUg1mogD0ovh4Ii3hW+ZtkSJE
q4NqdGkJgqeFRcnSU0xGIPCmgbL6i/dbpkga9FxZeSRwuDLUO3e0Kx/4VPIKXMcH
Ej5UR8MFnbaPpA2geP6aZXIEYy/Bggy4qRIwTmv5tZqJrtcKqjmR4m0OePzLI1OL
Ak3emfPrS32aUVvq2wlFnkBpSnOdgWrUtyaTFfaBDqe7ouAP9wJ2hjvOPn5q2oUS
JD2Nc3eJDKUY7yeiBWKsrmjncbmhhbTDRIYJff7A1k5H/2E56MvZaXaBUxnjxAXC
ZtW8I9B6Fw8GpPg3mZxUBwMiJQFB/cAWaGSCU1QYOc4tVoAeFUynZVAaXhhBY/L0
GY0iLtfkXnxN+g2ptMCZbWFvSuNdj7Is6MBsmxRNd1drY7dMP9w/XBmzNa/7aB7M
a/btS5gWB316mR3djlU7v0IiJvyWPQaNhxD/jJwxmBDWxbW4BeA4w+/iusvcqv1X
tApMrtDztj+m4+ZvJlqiSHvDuAAPQDgmdbIOidJWmRG5uMFrLB9dMnUn3Hvsxax+
I/oqLdvNIA6Gfwn2MUxH+y1CA+r6HQ3mhETDFNjbXjKIerIFqIhZDmIS4BcjZbaF
GaT8S+E1/KBZ3mEpRNa6E1w1+qNhuIsK0z0w7sLB9o0MplaIva8BuU8uvdi0Zh+e
tGLdidXLKGMlHj+4CkrCbT1h9C26v4JWYyjwpEWllDst7DFd8eii5pNYTFVMMjwG
1tNNzUzkK/0vBrAuwTrwW6Hpt08/GTBVgFoDat3raZPUKnsJLOe8E+2XOkT/wGCA
lp/6n5vC+awtMRJfZaP6zg9yac/2Lf/0++y55ujVQWho18HVuMCpJmNjpky2BS6i
5QV0PXAkHZMf4PgRHv3ne16JuEs9MNp3Ax73r38SLfDAqaBrEjPhI9VEhsk0zG8y
Hl+NffLzZkT4qytCen4H5poFEnz9ZTQCm+oQDrWZCHpdmz8ymdQ3l7oqGhoT3m4h
7werdyAqi9lXWrxBTfguPbpLeoGvfYJDXWmSFqSSjy8ybJBHInJYZET+mEDk5aS7
jdN3bl9C/NoxPZfZebwHHgK7MHnz/XN7//bHgrkyeCfTLSl62d8Kq4L64Twv+OCz
7lEZU/yFaEZTg2/0jqyrnWVsfz8oM2pMuQ+yWsj8FeDW5OJtgg2zWEyf6rXYkWOe
0zrt8X91Mmoi/MYVO7UH1R0SJEA5+HPNGcLg/JRC7nh8YAWiWc2vqpW9f6B/Mr8N
6VhTZXjR0T0bdD95YxVXqwZK582ctKoDHcHO4MzocHWt5UqjTWg7Wy4ez5+kgGp3
vHVxXSIVJ5snUQYwRF1Q+S4G+JyaFIAouNep8BlEEaP13nHrGqwH+oOnhvQ2Sc18
dBftMz/Lbi5mWcHPP+WiYEukywqxQg2M7mIM+b3WgrNDtL87iBVtTFt+xjEGoD05
at+xGibftrwaalyoD2C1fXEPGGIFYBt6+AA/+OBrUURvcVHGpAnD2UubTj21gKPm
X9HVlpRgiaFCSMR82QzpwK5T3NAHSGicn3BaIwI5fEiIivLoEcrMBQKTMT4aOlAe
dOgF34jO2ZpeNoTuoMRphj+sSWAvzutdPYY2eDWTThEQVFtlp1sGP80uywm7hKyr
0bHQ9fBI8sXCJ8KbV918b5HwKNI5TONsMXUu5jWFmXAGQdywtUvqAGsiXuIE7X3k
PHuxRQAnSFo7yD6U30dp6rKYEBLI22+yEV52GwTIOYHL5OZVv+V1fMjpRtsusqmt
kNhI2YpvuP7AT0GAtOlvM0sUSibXoZRBIjVawOfzfVN6DP3VVCfL05Q3TbiqGX4d
qoljmu5A6qZIJHpmOW/XphKq+alRLKxSOcYraEcPqhhIdLJfMo70HB3DKn8eke74
dxOg4p3JcFgS9qU38rpPOOuLEb3aLtLYyieU70nRjNkOtGmSL8aWSAEGusB9DOt+
aUcxQ7//LGGZa1HqZ531XbPy18pa7VJCKHTEo2ViZhr7qssZcwgzdjgbYZosyJX0
yR/0g3AHdfxNqgO/O9xotZd3A3j/wpQynYeZJnROy50yAKuVfHbtHq1VOZplbfsu
dKhTuvSDnPq3tRaqA4H3PfMxeT+DS90YT64Vc9B+xWuSjRNjTGhk+RRE1BYZiIwk
7l92L7dL4ut6CjpzYa3ikIE0SZYY7whHhi7sCzNqh2LHio9LJwcoXVkDuZNcHGgw
8tOOc82otUS3qtKyKdQiL5m2QzVqOnV2vNPEZEhsYtM7TDMKqtr0zayiOnxBf42a
/TdVsHtVmwNWgnhPwhoHXPp6LM2VRCcCGSI3UCY6jRzIs1jM/FNsToFsOZkN1LiD
b0byzU6nYuvCi54roMPZwCbNPmjHm2QYwLLAeBjVBoo+NX7jpqCA0Y2QMG0Q9APO
xR68lYBOA2vheeNrsn1rHol8l3vEJ6WWqOddQ3cMK4aTWG4pMFXl9hAyIA2Pp2XW
EdcclYQILttzxybeXyPXPCp6MlURlVhwJMj1GH1O3ZBGZQM1N8c2njJIyuPYZyKE
htUleP5fGNsgv250CrZOdaz1bvpGkBY3iwABbLW2SF55zQhksZJL1TvVPRZzRkDd
UuIvalrmHTF2HuX5DFdd2xyl/pcz2V5m75k4dNUYve5hg6nbKxd0kFOpcriVvPfa
re7V/uuKVbzdwEDhKzIQ0lO/ttRAAjQmnhXOO4+jVhRPnU6/iKTNkTMn8Bs3RBhg
ByKGud7xWWKuAvorwPIP3sqOvUdDan70m5lZqcS7+abuWxQdpNWOwf5pfhY6jW8q
Hhk3bLI18GmXYgj/BkEgw2r8qnQ7KOCJEYTouqzUdWTR/ogp6j6tbLNpiOzXOp+v
IJWVz205wvnpRBVPz5BeWEJkH6c0LtD6FvmT1d9CMT4K/QKXx98nhJYOiOZRsEh8
6XbjqSyZV/rRGLIjuRu/MqzZIpWh8G+kFyqfStFEhnDU7HEGrUPvtUI5qqi2qyhz
XDDlYc5TE6SYlqEG0wfzGOVRDuzVgO1u1gGL90gTbISxwmhj+HS5C1VYyy1UuVJs
ZmgpWPwhvFRCs5UhPT3/KQjvQEWJfk1XWJ6W5AbhlSVNB6oXTpAjB+2GRQwrQqrn
GT1yYWrsxVhAxvELxTDb5q4XoSwt8t9C7z3/1iQ+IIYQUfZBkd0ZSSvfcTz3YxKo
6TGNNhKLwqwgntEYY9fthBgsyY6QOrbEQmURyj9MQov1AaSQicbtzg2Ww3EXgAtg
9s1vVJTVcOJGYx/OH4gGYw/UHgnq3wAVxmRp369O0w5DZ1t1WBXsZbdwbl2OeqaL
kPKUvtkg2/Ah395B4jq+KSxTeY9B7JQRR/MswQ/0b6PqXdiuxulR97gvYRMOvFcC
mD6yIREvsnCmWxjwABlGENJ0nn9zA4uLnSnz/q+tSP/nQ/fnYT7GRryqU3PMLq2a
fkW8RmS72yAGgya3CbyxeiQ+I02tlaaVXERZ26GYKWznMQpyhFoXg134P2JbhCzS
Gp7TlWpW6Y1FQ1E/oKXaFdlyTa5qRvzAMcnIauFdsLZdsqQILsZIDXNYnwrn4Rl0
wf8/mpdc+6wn860MEI7AA+r3r1eb/pOQt2t5U3sa+sWOqS4BE6m/OLBo1G2ZP1j8
o8qvfQR9QdUNUqZvj7Z+z8PBHuqgWHspv0LRwc4b51RYDTlcGpjSvLBV1qh5U1eB
40f9Tia9XadLeVMJEiE8dIbjXvAADCCf131sboclEg65nvELb5vf9X/wSw8KE2nD
daYHQEw2jzrVNsPk8o/j26qUtr5MBo48sbrJUFLH5IONKmL6oe/6hxke9tDYW85m
zXQULT0JugF0OibVlwyEwssip4HdPTARLHXhudq/HbbGoIMZjfy14HWIx9aZymGJ
i1NV2FVktqyUm//KDBqKLlZftYmSRhW6A5xxqJKLL3VEGU/iJavpJfl+wA8FY8M7
llruz2ezVhfZMXR9R3eimkADwEGmSHqsfG2p5pCpMSqNhZN3BsKgaH6CUFZey1ci
KEhR4O0s5hSXSixL9K688KlZtcJ8/3nszz0u5Rk8momxc8k4hQc1T52+BzTnT07d
mRjK+JuuW7RJUigScaNxzJAlscSIzahBgIcDTtmyWtg6konGtjCxmPsNsPsHYqqW
NuvTNJSQx7xskxd4rbxbl+PgA57kcnBme7sid4Q5rvvnVzJYZohLvueHBL0H1Ara
km6kaa1YFeGZwfdzN+VOT21ClaX6Lr+igXdDusSB7TZv87hllxRG7V7w5yLAwDiM
Niv+SySmGNLq1hpu4yCGTLBGPKhc7i6+neth469JtokwAaG2nVJ1CrkS4aoiUIle
xhP1u9TLgVwZIuOaPM2Zu/cp1Z0oF02TZaexgqFeaX69Fyy/PvxkKOJJUKW4TV16
mJfpG3DtBLF3yskSDk4cpqAIY1HMSbU7kfroX1IlOH9FHoBoGhBawz8ojsSKmI7j
WfM7sqMusI3dga7LEnqbwPvNr6xAOHVjBx632o2RQ+xiIkdicmCPlrwLqtBuQA+i
Px01rmJ/uOs3/vixiIb9RTh4z9TnfRiGMNN9uK9G0vJlaMJvbYT26eRGulQhK3OL
quIrxzpdwpFqEUpvRKO+Go7/QDIDX+hzs5JaxoArtsfMhgbboCwDHfIQ4lMpr/+J
Bh37WExiXnJ4S2oHOGi/f+voEnJv6SRmqv1ZwOIoK0Jk6LiftYfHci9KJtl1m27f
N1Gsoa1oPuIJWKnMLPY6mz/ofRMulCHFdtwNYLgx/i07HA7bImVlHF9DKhxx1Cxa
vj6lKJtpY+RAGyRIEk2uJ0Dj40iNfsfLI6X0YeBwnNnPSN0pr515G0u7DLTMgo4k
9AGHeYMfGqhYbImCz/pZwFfmtqcTuZ+lAVZiH7i232wLChBYmSdbNrv5/EfZDroz
/jm+EwYsn9CBX7BSo7PupOpTHQlLfmn8KTMXsuYzIG/K1VudGn+dV2fYIw6udm80
0PWXqplVet9adD4KCDGlVvZbmNN/1qfHdAzAY8Hb9Ca+aHOQOe0msDVBhRc2+Qfq
PhFtnG0s6Zf+j2CghGhCmAxo+9TW/dYTtfl4kVeICYmHTKZNH0rn1Wj8GIWjIUUP
/bjQP6kJeYzZhLFWgF7kwFfkwKnLebZF6OGt22X4urhuMETDtQ7JhZhFVUY3Dxg7
5fN34ZsDbq7M+TcWALOGoECjN7wKqo15eBNar2RV7fVfDA9Cs8JwZOqPjac1Ch8v
7Nx5Lw1vYO2L+N+gp+0SWawDGu2N4rB185V6JknWZ91s5k8cUVd4pVWIbnzRMN/C
QGMnI8Hiqy+RuSXv91UGN6SUUj457PdlPWn2Wq+LIxXgy7ve7JCKyyDsoBSiiqPV
HV1dJBeX1Uuv1iOCiJdGag75ZJPFtbsnI2UV4RzqUqnwixUYJWJz2UPYlvK3pK34
+l0c3ZCX9CcgTCRCVn1MYDMRfQ2nROTZynOrsTnDjMxMlC5WSq10Hb1CV45Qjf0V
ZTDqYXpmlHmzn9QnHDHvSxwcNX6WyfiW6qt1Dc0hSNMa95nBUR5m6vgJY+KExPK4
BeDQr9Ojemh0+2TKLo3xH7g32cBdNBQNFM0My6re09tHvWd0+pSGy2oIomqWc7pd
JGRfmouiPBClyX/YYHfR4xZNXPAluNicmdrrnCNYb4odI3QbuiaFbSnVwGQFJS8w
NzgpbdkoAA+NVCxZIcRfrJEZ2wRpxdH672TbVtrAais22fBuBMT8O6XjGPZwbv/s
cYbJRgqKj4mpF8VB8PNbL4Q7DUcUgQDSy5eSAqFtIZ8mnQ4BzfnFRQ7BHDaYRoC3
YPqqhrZ5m2bgk6Y2m4FeeKf5S/4GFL4aIzvmPOgQOuFXh60SUux+pPqMpocc72uq
2Vm3Q+EDTRaS+Kl4CsrGfVDOiTbN1vTAX+ZkX84bJV/OWxjJKl7ipHq2Xn5pwJ9P
2f4xN32irTlO2uOB6cMgeXEYcm90aYReocCuHXJ2+iF5bi6dp7giYzCk7d9rkH6l
seLOjQ3ueSwXfhxSpU5cjKSsNp2Uk10dr5fvH+L5KDLLgcCPruxYUOGnekizIwsl
Qb5BKniOTIX7G6QPQl9PHIbrPeIiyHfPld1adlSQidnY5grNx2TwcggXsoFpPAhY
O2U7cHF4wstk91v9zYZv0tHHK9pFuwvfmDf4xrooaGxTPXmzopqW1/t7SmGr2H/8
icJ8QfUxnlJIMFSLJbdxinOWj0zvDmGU017BRaQk4YygRO5qkw8+I55RxeJyJ3gx
PrZSFMDh/d1z3gPyYLdWU3HkyNVOYnp3q8pIw2VHMAg/h+92RO8K3oM1vi2Lj1Wy
aqxHVaUSmdxl32XMqTS1Dm9oWP5MmDqmbBbPdVmA2P92e0kQE+KA+5iu3bzYqJ5g
GAsMez2a19iqFtEV71t20AkR2DDDrdJP6jWfdZATW7h0RDA93B2LnjYOiy1HaaGL
K6tSE7wlFWz7cDwKnMpgAryqtWp/+yDgz2GXZ1KI0uaWDnWCpQDhVZMOXU3hjexV
e1jNA3c0u/YwtU3P0X/bhF1+diDPIaH/jk10seP/poxawglbuWRm88ghPJjAzXpq
rimLjTQztBLLD0pltHZXSEwiY0T2RUiGSRyetKZx/sPTsNDLW6UlP/Mr5qIRwkB5
H74gjIZiWgs+0MogqaUeOPUzbcwI1UW/MSuE4E+WN2EmJ1SAxdTkJUCt29Wozt9t
/bSVWZTXifSGgqIyIhvksAfS/tNJzqhzxzhvCK/nArOMxLNb2DH85NBTz7K2Kn1s
WtsKtE8H6T2RtoBvPsPSJq5jaQMLZPeJUYjLHoMwcVBc1aY3u6XFQqNvyMithPhb
GlYauEs2UAHFwsWn+IMc7BO+u22FpQOYRtFxdhy6r+C4GBdyUgs8UYbwDQKZBz8D
+tg9NTFyS4r+auCzLp0LBWmB4uMGU6VcCBAXlWquUV8d6/v1w2/aN3h9cnCN+N6S
ScSMQJsou4ushDSx+HYGtLHZ4jDIFuDvTczjgalqltycsA1ePAtuDhJhVqe9IV+h
eYjnUgAJvClDnlj/b58OFedaiXOahEyha5MKryra8vb86woRsOQpRgK5bqiImT/w
QZRs37oVr/WmEsFuyTNLI62yteelimrom9Pkjrq9gm+nHSvtEcTzgfp20r9lg6IJ
GPGjZB8nqyT51EJpktPGNJNKSNbQp+Jc/xLrspLgdYzDkhzyOKBoACnAs7C3L3gv
PdrhaUL5+8FpvFQv1bkbKnIgwGd9Zmgi8/hbpvKvMLRdfWiBHrHW5JscuyLzkmzv
ANQKvzrCrw4NsO+Q3nMb3eMcV02ecGdABd8DP9i1I4sAE/X5g9VaHBzqSBzKB5+7
YtWoSWTezsv9u3KTeIDyF6lUASwfQOEVKb/6WhROFJOBlyupP5evvY0Yx4RWTrOD
cZSElfGVB8pJwloXPaEXVnMEWraZeZ/ywuTy1TZa672UYpCbXx6XP+T2rFL1d+8r
z8LVbnCiT9HX3oZu+H9dzyEjT2RdSRiOFp2NFLZk07kCgAibXM0q7qmIAXzAIgLf
w3XUwZytAi/lquP2qUBGaslUNhdTEjTrEHKcjTBgdLml00djaCUCJyk0pJ0eX75K
RyJnDPVstJf4evozUZ3an+Ja1lKfP4pIaY11u5VwD7gp//uPrr+8kDQrfP7KJjOa
odua38NpB+Vch3PMVjiLB2+RlIsND8wWV6fcxkReFEQuqFgPboGwZBZVTEhHu6is
WMhly2eCBMjVuAl1xfGImje6F9O7rQqZ78fpV2wVK2AM9aK/l0dFCNWmMH7DD/o1
grFXhNA+q73d1QgZXD5F1RHlgJGnt1Pi6TjRz8Pdsi2fLyTUBVXrQ5sU+ZF6IiFG
rGhuUlQGFYUO8KA2xvhhpUbqP8E0wFV3Sbb8a6QbwZDBoh1mOgRsy9WIu9hW2qCu
ThDV1Qr+hnv4nJMSbS2g+pn3NhyhxcyRjqGg8sqqOu2/rjhK1p3LBh+cRW7Jc8O9
aZw9ypQ5OoS394b38VJv/L3AMhinngEUOzAJ6x4VTDUpXRsBUCuwAppa6j29j7cI
aHOqqyfeu1dCRVH51SviHv3mSh8Ida0Kh1XSYVmWl0Fsen+7uf0fSKte1AO1bICR
aH33mBdjeHqJgeCdXVlhSnkgCrjpbZOxpZDPlbtB9h/ekCVUAngzecWkeuJSedsW
tPO4c8dGUw7Vm9svyiZvEvHHXnPastW8rz64+ySB3n6dbJe5ZXwWxM6dMPcJNdBi
DWw3JQ/g88KYJNd5CuZhKtv7ZivhBSMOuYvlaycalQJd8z5L0B37wW0/jHEbJYap
JgIGp3Ojf52x3AK6SLqGcdv2lIqkAkEyV4/71tUUvkbUpaXi6rAbeKFCvJ0h6LMk
Od2mNnL8d5zCzMKVKgsFZhTlKMtRfL17a0dF/IOl/ZqmLEczzn1dbM+bhk4gU2A/
OgKBoWnpx4ZUq0DXrS28YAM8cL/iubrBlxd+tdOjTQF0OBBFoKG17vICR4JU7U26
uIdSdA0eUcFfqeDKeu/djJtC/PMY4Py0UJfa6RjK9F0kdbRb3NXaTyTY/+UN6qyy
KouHciZ9uzhSiMnob4Xw/nLDXyvegqWK4n9yKAz+YhZyYeNDfcyC1PXGW68E3Y6T
xxGYl7ILO0AOuIgOtAr/yOtv2qXZC94MExugyHmpv+iiZo0pSCEFevV34XVOHtwr
MSsTzyIOHhLW+giiwyZaGGd+rnRNoKK4Q3e4rsHMrknYrNIcZqBkKRUSz/UBIEZu
BXh4YWkD0HJIuEET51ebh9+SvGiKkDrgueePJY4Ns3NMLjtNF4LlgarNQfTS1+9A
55r9BX2Eu23HUT8I3hTC9WI5p/r8tvrsZgngj0fFu1pxT8uqCfhBIJFU3lWqq8Da
dRD1PR/R1FTQx5I1XdZ9/GXJCRo84/iW8sF1beOxvs1aDKJOAhLa35tjsOXCeu5F
8emz2l/YLRGC2YpNOaPkwDJiEh8L6ZBDnsIWL+jWKwUp/9txTEp6wasSaQTYAohD
KdFm8ejWljMkxH7JiDT8QUnFIoNqt9ZX3UNjJ+/SYAj5gjnTODoUodThFAiYKC3q
D0kLjMG4NAIOifOJoDf8HsHG0DNLtzD28/QHRDArJ+EHEpQntKX1srdGKOUlRMkv
4jqkMXaZ02t1X8bLtSe+UcOB3IbXcfGiVJ8kMph/+K90UDcqTKPn8KubafO6kCTI
euOgPk79jCPtq/PDrQm0lEXBVE13M2kqSlZKqVcSbrsgHA13DtE7Owp1xtCFItRB
eYfAR98OtXTChKdBrA0h9KIbf8LUSNpUueQ+7RgJVVVL8eetVlj405T0s0X/Np6d
hvkQP5D9viwFrjB/Panef3LezJj6hH0EPr/CRvZ5UH67S5dyc9thsYGsU23kK6qt
Z7rGgm0o68lcO8jY3jZgRMivRjUHoK3NMfntQLbVkwV8hcAYKrZF33dLA6SI6wgX
VBTpgGhbpN7ly/t6BBQoH3BWjcjZdAK67CxzJn8jMRg0+R8YjaZ4s+sUjmgELGGp
wNyhezVZZ0oCi7fQQTqCzBk6TTw5mWRb+F1c8q6BHd4bGo1qdbBqWWi12bgDeqnf
KjGxt1Ny8y+3maK3FhDR9I2l6fVjtzghyFtA6TncOvH52UoaE3T/2TLh+UttokMx
W6T17gno4IM5Tn16X+HixNLcyRh/jbD0b/t/6WH0bhhtJqVXqOmJdfhk3jW4TXNR
GJFpPZwuXDPLzZxs+KFrjAInbZFiX+y1xF6BFMZB4d6SOk1ug6yCMKMkN8ZEO9DZ
Cayo/L4pY8JANFCQwqLDMK2wK/KOMQQdltMkhpumZo5ZDdP3TB8fZaoGNBSzuPip
7YsRR4B9HlPhmyksJLj6U5gt1DfZGNdM9RssxIOlEMGBcDaU3IeTt80F83LVTP7c
iGlBY1cfeSg2feyiWu/FuYmn4N6Iv7PJb1GvkM0duOR97DaN2dTdzX4hY+65nPOn
Yy2SdyNF2OqSkv9QF5zpR5LsARGWckeBg9zGpFqhlncy3c+MVpj3rIel1lV5Iq6v
G04h2C8Y85QcKCRSsUVE2k1Q8hHp/70YgZGmDzhA9NAUcBqz1iBOIqSNLMZO1lhi
8zx7D388WKdRKoVumHskUDcvTnaqzbH50vEQgcMlQ1OfmZyC7sAQaE5vwbU9qTQM
a75iUWyV3KqxIXpuvNep886Cu+OKC07qjc7HftMPrNNdSGFL7YwDfBsCH0iXB45l
pn83weLp+MNN2N9FR0hPhuzXeuFIHv8EgMvYIpGMVyYXxJpZYZ0Aij4ND/dF9Q21
jFHtuwe9t48925qbPfWTHcgleNkcpKx1vNrKB6XJZtMKZKrlqIBAllgnpjv7GxpK
0RqC/MlS5dJUpsSVobSuEyGzYqJIVXAPwj+Pwg/VIVjTz8wbR/uq3iVALPFtMGox
wjr57CkIY0AJ//aLlEWZVvgvvgozXHCnammzDiLh4Yq0/FlZD8b9lQcOC1rwb9UB
rBAUesrUEE+iH3iz/WUb13Ws9xGHrRzpPya7HHnNrb2ojSN9FvGDVcXi6q7ncruG
H71Kx8x5Ws95xzngk8jfKkbk3LHm1+WYAhKErSQtiRhHsoRtf7fOGxqHKc0aJNda
LZL3e8zyQzqZWrgq8bZQcAKkfgZDvY5rJuwm5yKFDesvjRKeYKIggtMpJqYjvG7f
xHqYJcrw7ODZbh1SSLIZttSEzzH81dumSZ5wLAXg3UrmQUPD8Hrl+bDJ4ncsVz/C
4Wzx+OFL8OFx+bw6YsX3/YoJdjGRq2eSB0F5A0C8qdoyvgpgUmXJASe/4oTq4eBr
qlsD054q77a9t0ExCJdabquiZ8omLyFKJxvva4We272w63a4JAy/X7aIr5RE2hNW
4rsLYJB12SpfcM2mP/pA00VKd0D+hvtduES3dpuhWexPkepmMqh/B7WHyy69+Zsq
T3yZNpUZWmlrHZF0+Z0RSz0ParMQvIe/d3JwB1WmYrxTJCN5SzfIMswdzq50FDrK
jdJBkWJ3k4OFNsg+jnV9yFdv3Jfn7NYAj9g+V9QHBcuzRCN6yIZb5I9kn7e4SP1S
p/RDQpjAFzADnMkyJCHEdhvQ+Ux3pE+S9KXE9iIPisKUDLXP3rVpKW4lnjUtO9pn
kHiYw3IQIhKS8lHRoKaOZHAbJn+bAnTXBYLrcJfBRWOSWgMr7OOs20lddBo6NYsa
aeUBZJIX9Xa/vfFC0fPPANqWYRtLVP9zchJyQE0SNGaifBJ5E7ZciSp0G77EeY/W
gAVW2iS6YFKU4crK5p2IkooP2+Ir4Y2iaiHKT+2Pb8wZZYQ7eyPqCk6M+jOOoFcC
iUH69FfqqJjuQ1RLpC0h9UA0RtmObdAR7kWg3FbHtBYc5k/99m941YzsbCb4QNtQ
ljwTXc4GPemTC7RVmzNmqWTwoyshQjkHsJOK928X5GLAC6YlN8D+ZLVdtJ6rTxqV
rhzL6Eg3R/Dsji2qbplfzDMiXVjiA8o0+CeQlYa+fKhrNm7VoQ5jVANPG+db6lvF
eFynKt3MGJD21MzRuwO6djJUjhGUPjwW4TwuhhPUKMZdcvc8a7AGx22ZvHiFkB8P
vkS64rSiikO8KCUqikPymHQ1aSh7by/yeHVzySH5fL8wWVsfzU1Wk0c2WSLozAQi
/CxKSeFz4miYVUF+YEzNXz6gegK0/VcAsCTcQYI97VzCHtlXC6k6R4MhUzRQ/szc
7KRwzDkxX7cPdiQOgtrlA95fmN/sz2YpDrrfp9dhV8GKNQRxDnr54fNwGA1PMTvK
h9eO5AvQaiYPrJFntXTkx4u5V50CLl8+jBoV2Pb+NFAJuIHvaFuFk8tXtFxuz9dH
rzCr3X5EOpwh1oi5UPut4gKTFYNp30JSz2M/f3ienP4n3Ad2EgB2tGz9D6XIXgzr
qWzQk2qiYq9h8rLdGKD3VrA2Z3X4WfwkIg6oW7gxqPppVKMcncSHBdw23a916d7F
jikGvrMEMjALab8AujSlzB4G7qSGesKGuMpIqbdCByT5TTNWm3SeKorbzw2mOfER
N5xmPVwPLaONYu5r4jzvfdM9SwdJZnghHA6FGpGMQ+ZQwUYFBxYBu5nAxj7v2WEF
396A16ROR0X82hjHGgxZyAl8XHsha0emO5cTACuouiJ6mR13B7mn48LPr52W7kV/
dGRWC5k43uD9xpPuIdoUc9BpqjY1odfgtbklJ2mLDKAenVJytEm+Q1E4WQk3hH4V
CrWLbxMNnqbsoKYyA6WtXJ1taCewL9Y1pJYxkzrq3mNuH/KxQh7LeFaQi43s/ACr
B6JfNSgLlo63wPYG+TuVbeBqnxa9wOykoZQUxF9nUAo9QkDgi34cHKts+opnyvqW
Qmuy1zbTmF4915orzePL1crbNaWquWYtAV0IMKjNFBzZHTXusobO1cCunldGcI0e
bWM6/RMYL6lAXQTIyL/VNtizeXhk24VhnwXx7PQaVHnAhnfmsj5dJXVIO2oiO8iy
y9zKUTAP0/JgTZupHuE2JCtc2FquXZj5YW1Zswm71Dj8lAj2DqhvVGIvlQZqX7qy
ji5UGaeBFj3E2X3talMyV1kh6rw/eMhJ/6io8i2Ka0Z9krUCQ8aWdR8UFVUH0Wqs
pLEtOBdU8j7Gi0IMRTYXdoBJ22HKz4HUcFCkrLV17dypu3O95jYxdAoe3ns5Z6th
ElbV60I4ieLUKXfs1yE6GJf2qErnPlnIV9XGI5FTuB6UOFNbzsnifXpxnB4NndJP
avJJZKOdjOxnEtBX/imgk2IoWntZ9csQIsH0LH5GS5zrt3TNtAEaSNEBdx2k1p7w
q2c9FAKUU6AnGXwgrWTn+j/dOxvLnvuktTERNTiAzJcZfgA3/8iGrE8R8K0m62FT
7/Fm4cJiXKm+1IBewOh7dbdYN+xiUBIKgfhpWbstzz/zWpUJrosxauHrURXeALpl
g5hOgIwKaAnAPNaQt7qzXM5feempPhDhBI3gU16ESJePvqv3aHVvj2tdwTw5IVDa
JTB2ka4Df4cVXlL3rybBzLjKzWOiBcxWiVQMaCX359ZWrmnnEu0xRQuDzlZJcdpR
QWyH8/l/59bGNWUFKpIxE0b7HpuLR4gRk1CEdAbO7+GlPiIVB7BK62NTvSdD0gPU
1j/bxFiemv1Q4MkvaJD/cCfv1oLVfrWtZgvuxpagB59OIIIhOzGQ+LocJUhtPbGm
4TFyKSabzlA4pNELGE9/fbIT9SWrtFjVVsDGYZysCwIfx1GOtfC+DXS+tzm5Q/91
PaCNaSz+uvVodCC9NfbtdmvEyO/go35ee5nh1uZ4a/36X+7BSGEnKE+rdcix+hzp
9nu0YPbhR9MnJPyz7Hr1jhQkpHOCm/3tUaXA8fkk8pO76Hov7zJ6B3u2tn+2km/Z
xRCwZ9WVZy5/WeeQ7j6e+hQrilJ8Qx1R089d4f4sLmrnAAgjrctIBeMAC1/rBdbT
B8S6hrX0ONJ4k0KJBcAuqw66W4kRP63vHjM4tr23nZJ0V67hDdIrGjKNYpErQwuV
9xKXILjiMM34hwM/hxkcNo3eczUak4O0lhEiEN7ox9iMcI81iUNW9cZxkvjPwUsz
NbnbT1kqp4/zuDtE6jeLSVJ1JadnQDtBgoBM+zGTd53G1M7q8S795yiuyK7kinh9
5Kx+HPDadCy5+6sNz55Rn1Bh0bFe4GhujXYmFAktT9VjkVbqcQvlXKqJvoHEAkcr
FnpArm3xa7jqcd4dyh6RHJLL4fRYYfzgmS69Ikrs6tyUgvYTf/DcO1Nr6wCBRlg9
yLGn3S5ASERckCUyij/d/TED1CH/s9Xb3kN100VpNp6YagnPZQqxgwg0IzG7xqRi
tZ48ItSxXP2GkCzIPRlwnWFI+flKNjcZRHoQD7w60xGjgVAD4zYdz17Xpr2pHfbB
v2z7YLIkSX3uVwApiAz6001PhifTfE8BgOnOJUnrkaNOU7f+16O0OTil5o0CVoux
s8HLUfKyG/6+8X/9bCzU6ht4AWkOqolj6+H3taGIhdx9IokInvE16AQp73+U6baI
hAUG4B1YPNZMNoDtG5nih2KhzVpjuyZiEFaYpkXrQiv+C+PahNHJ+UIGHvvpsALJ
473bhjEFf3qZ5CW19yCYNCcbkUsSmRX7H74vnlgwrRwjTdEXE0scPD2pdfxx4/MY
kyu8y2sNezbEackbKgVpSHtdIpfdiyg2TaL7nmqzVPuDnCac9rYSidPpkzqk28Xa
rSqQB9iZgFZg15Mj0KrB2ZfL0OzR0vsDZ+ZDnB35NRtDSU8RVgBWP65bCg+sp8to
pfYFSEI6Tkjz5ORlp7c6Gdess+k0xFrfQHDLGseEstCy6WBMyJ/gq8FqArGJpF79
2W7qXB8FoDrZh/Jy5K++L3pC+SbSSgfbTy5TbpSnJcwQsxxmpQhrnmIr+rLkkQ9p
YKdNQ17KOajrA4SOlj6q6GWGVBr07+cL0bgJLEekn0TeLX5Y6IbXyP5X9hHwOtus
NcOLwZ0sqcYs6Ka4SQJW4glPmc+JjF5tBgZs23XUgySZGKiU4Xlt7w7JYs1eQhLE
5M1rCT4DTdRwYx9bko81CMAipSQ71rbNgdjayHVQ4FFfXFgdoPtWKtJed9yCzkEt
gb7tmxGmaBH+1nqwp9Qpih9gXrjLpWF2en2G9xnhsM8HJjRoNPP9XC/zijET8j9b
nEHH6/Ne2Iiv3JRitruxosgBwkyNSlHLDATnJ8Pbo7jsFfXhU+Fnb6TM157uMjwr
RXj5VVNEDC41UV51kcxMMlQyjH0+dKGogSNUUvbfFYTiiNnhfQmIViOMjGvDXH7t
yDnTBaUyK1SE8h1S0QAzedwc5Z0TtX6bWQvfnLxcmpQPVvmXhPmh4GVKjbzCyW27
SayH1k39NIG6S4vLABrSgqBc6X0XBYPNJSr+0oz5xA7Qugon5YE8kw8a38vsd6oN
Nazkpsoccl1I9UXH3XHgWKZphkYgCzjzfNxUdLaGOaN0Tx5U1v/kwQgjhN9hbCEO
VQEx8tQANoppfWNrpClb0iiePARf94ShB9XFm3D2EqhsXD1/FyrHUYRvk2CySJG9
62Em/JlPfKLP6YnAhWYtxvo8sRfla4QcgSXPjFC8f5FxGzQ86Da38CbIjwsLSYBi
p7nYIbvVSCrnSSs3Z2oPz89RSqWQoL6/zJJYEZ08z2lvrPDMKTMgiQw6waMMdWy3
NxNYuYjy81E+LzhYBXEQSbp6mL0xX7gLFfsftLxHztq1C1gNZR0SOOovs19wPvYW
GmdsqDNdawygwOM9BBe1LylbeaOtisCcnGExuJFGIYBd3ybG6K9NrPTk+PyBX1uo
vOv/g5tRsNrXtGNpLaAvPiJIui1c8fLxMNincnjzueN3Wnor578aEDtVS20dSUAi
WredbkBAHfAjQAo8FEbSgi8YRk9ajUQ/YK1pu3IBQcnxcyM8cT6O/9a7DAsplWUs
nPJ5LPvILvdYch0Wr9Ev0cMm+HH7C80Zb9JLdba+uCJk5FDyFZ2LBiOMEuNMlQ9O
KXs+B9FHt8nHuGgcp4C837MrmN5OJvnxRUaUjQx5MmwaSZNtKCVBeylTy4YhKw2p
94pu90OXe5UEshTi3QBPBhirQb+CHqBjkKX/vYhMyuJ/rakDHx4nIiFB6htpzgSh
qk/Wh4NDi6YcBpOZUhJoN3aVwskjVWFbW81DIo8kg2EyDUgeSs1WvCZjS+M2kuNh
FYiNEG48MyvU9rynOalON21lEYkalHkNjG50uJrzhHJGGWB5ImEGaPb8xDlwKFAy
Sx8X/u1kR+7I6hgWwljs+Cx1vusOU84Mr7/7mkMH9QYXpCXTeyIyCTJicLe/vbE9
D4i5LcuGDj52KK9oOjt4Z2kxqumSSHUINMsKugK6WI49djyPj3+gl78ilgDohS2n
X4WuEU63X1zqIwFF3hOH2UtvWmDN+0dIUtT4ggTCvTeToyn0ottFErdUzJX2/oWA
m6nENdszD6zJIkxqnA3rSHCslZK6fojptsI+71N9mHalMq0RXdvAIlXTEK3CVqnQ
BCtgZL140Tuv8uyIbxFJz6eLCaSkfbOI103jqz1DKHe1f06jUH/Zd1BzY/gTU/uP
T2x2T0Kq7iiqVd3C5wL1sHJzSBfoxocAtRjrJJxVguyvjEAidVEtpteR9vpz2taN
wy5CNLRmHTcikwIiVAlagv4mfBOvqvUjRJcnETLiavLHyZ7uEKcbpvSGXAVqu8za
MOTFeqmOKL6X+5sRDL9i8p7GIfYjmlkUnnJhCv9kfwTZkR6yH7BpBFv3vZz6qCiK
dg8LPRpkJ+MbHMDrPW1ipu7n1GcJQfIAoIp8LJwEx3VXtdj73dpKB1HDTt5FsQAl
BHRIuPQgDyHwzOG8kRqfpMuh3S2xb9p7g/yMEkrRcW+D/UnowZzI0n9ehixQHs5+
Dft2y639PzxPQEkqC8fYv35nlut132U7TpGm8KwAzl4E/oDuF3LF6xjWq1Sc+RX4
pKANGd/rQbq61Fe+HOvm55vxLuT3G2quHUx+XESu/5qd++v0NVm27v5r45udoCgR
85fUd2oerxk0uIyKty8zIFZQLFK3ZK+vVCcioQ2GN5XkAitOEwRdPPESRqw/4ZXe
/TnLVdDdhElQ6SgRGSKyFPT1irBktd/WzdUh+PRL3AKUZOQ2ceiRwQL2L2srMWjB
kDgvDP2dkjH5M2RdGP7W7TZWbWqhLfBLEDLLdNLaK82AMaPo9XYWRrj6zfNqAhkh
MlL+hNpWOOZ2NjIURTnsY0UEWrE37cuPyI+kltB3W8Yqnw5toNs+s4ok7C6fbV37
VG5tvHbpa0r11Xkf1hNTwjeyGuhER7iShxodbAZBMS1QQTzm6VpYSZdV5qPhWl7w
4oGF3RvhN1jkg/ecsKxSDEjfQGh6CwShSHdUSpjDsxAKl4SjwfJkvhmtit/cajiM
FcXuqrxutAJtb5VxPzJckKBprEbaL9S143z7K0owDHaelMuQay3GYUknqYPMEArP
YvHuurTdTiGnV/OotJVLb3SxjXzkJcBB3YT2VEQLNTsmey6fWhzhvqrYVgLX6HvM
aivDEplLbO0KqgWa5Q1ElUjVSq2JAd92vu9MdR4Bjqv86USNvV73OcoLEErAX2Tv
c4LZ+nes+0rDU3ewYP2SJgXRELs0JzGBBxCu79r9YIm5zJCmehaH3thPYkmK6F0N
PKV1b7mR+OZ46B5j4xjxkNBOojh4MLJeoJiPmn75zFgH7/0XoakWp2/I16jk8XEu
f6KRBm3YyCEUB2PJ9jv65QwLXDEG7pxPPFeWshH1eCkeoYtOLqhC3wR3TiXeUF3i
nb4w6nP7EOhxDY8F36cT3jgBScK30z3WbqDov0j9Gzgkm7vRajkACnRckYe9BpRa
cS1FAQ0uSZghxlpxb9b7a7zgdgv9u3bzgvXevQSYPi9Hra4Hk3WoRfL99kRnihLb
FFYjZgr4f8BfnejYlQzlLOD/OO6sTEhoX+PLaCs90s70tVGPgZ43rIyjL++8iJLT
lpVPle+arChZSmaMhoGvSAPOQW0ucA8oGwVOaE8MX6mMx2PGkRa+6ossBxIa278b
THjArFio/IEaTOqLaumz/vye2GqIxVZiKwnEAaBhFc4OewMcFSVRGLfd6aPeO1Xm
ep7Sx0LaRjHMjSXZPmRos/PXGXhFZVbLre8H/IBw0btXkJxoxGJTGtagUT0R3dxk
g2k8KIfT6vhT4B14eIbW3rxtZ+P2Aiq7tbgKrdzjeSl5Hxg9grRfh58yrn8oNFsy
NtJxuVuZlR46UNrSp4cTh+arV/Q13h+wl7OhaKOaL0zyzGHNJphEK4NKg5Ye0G+G
jOSkXQ14qFxjxNn8Lac9GCZl1nWVyNJGweLsBZooHpVcT0rKELbF0vG+DpKaCse8
IrZKP+8BkGVoh+7RZPQAu6YQm7j9fvDoWX2lI3WlN/viYTS9Ppn0BQ6nHEekFMDL
y7bT97F9sOhJkPUCvVYorW8gHTYzby/m72wdMKK7BN2hmEUNXHbbhV2ZYoxq5BjP
wbxciaHKFiJlK336jBXsyZR+kwKlCqhL7ZKNe5SReMuFjWNoI9JE8roJPtvGIG+1
rENjnGPoxwV/B38pP98XuBKM/dcIu7Ii3bRPKgkAwQzgp/VGemF1i3psZhBtJy0w
tCtWo7LWhqNte++KIEGvg+iYwf9Sj0vUwbL9DPYZa2KS2+KzPB0ysWViuzDG5/2g
fK7l0cbeS7l0L9eIr1ozks92R4rfLZJLoiO88UZ4Swan7S8GiBEMYK237VGK7mbs
YJMu+GhjQmHxcNPA6B/kogjA0JO+LgbhzvaoyA3LfAQhqhIo5Snm4jE4wRoU4GAx
tvd9P56vc746rENqQu8HwC8Z6YFSv3iyUKs1GQ6WusGW8Wg5JJbk5NBdiJdqoh6R
PQhud2TsDK0udBKJCLR3el9o4C30T9YXick6MimxcaffohAcpqjNyh9gW7Pv4mA5
E9hkk74H1nF3ZiaOfj7Q4AV33J5KwYOTCxNu70pr2PD/0nYTZvYzjF+A2rynhGPL
ypsnv/fTZC1bxFmA6Abfaex/t3l83lcYHkNfjZNTtfNSi9aRBINkZOSOU8omKaWB
KNMeAvq+MCjlGuM0B9+tCPfVLxymL0qMpzZ/CbJD+iJ4ashIxBFOqXGCLr9fXbHU
64/AHTwAOVqjzQJBAhcK3VFZl69PmIIClgMUTcJiNbg4hvGftijUj7bT6Dt07XWU
+jm+c/Q7bHiFrBhLZhugEROA7SoaIFz2uOR8y/b3jt3chHhcvUJtBqI4Wknpzf07
VcceTsDjnVsCw7W0gnQ6NGWIiXZzib6kavSMraU4MA0g7uasQSpuKBGsXqcDOAlo
4ZODG8xTcHVBrNgyWcrhTWhHWjnKCwC2hFDbin239rDzgRooMB5+N6KYxT4xsIYN
1R5HHCSTQnP6Hdvd8bPRr11s2ZK9IxquNvxo9ouU6V6imivPycDGKL/hNWSQLll0
t76QI5wHB5aklTQFyzaQVDRrxQW7CPLKbkFfQw5zf2/2dJZJT1d4WZJcCyo8lSi1
gYpGfU1LGJp9KK1uWiQ5X/xQ9fb/BABqkfPCDxZO0v7DR3A5Ai8DaJVww4/nSGZ4
jWisuO02Yg3LFLGif+QapCdIlbwGgQkla4/CdP+YDqOwuRi3LOonSQZ3iKW4eGj+
PT83RpMx833zITbZrogKcWWOB4KQ50UQpuMtykLmIdjIC0hn0FQZrS8LVOLujDbU
sSvH4QnlCQ8XTqHyloaPxKiEwA9PwzWPPXJ5qHttZBZu76ZDK/OoM/X4U+Ke29W/
TTk6fjwrp+PFQIwICLuPBF0AaUi1E2z51Z5PMrHlsPLpifz29f1mkKFtp7vRTquR
foJTe7YsWp7/h3cRA2iC2I40NBNJqSy2r3LpPrFShaeMymC+jO2g3ju5U0Ez4lUq
p0BXj3quV/78UZFWrzJjv6dufjw11ipc1RwjlHA95LbVYiizYYZUCG/hfyD3XZz0
tdqowu6AsftcmwmpglZu7Qdq7gQtIUNiv6TKDDd+hCiHE+Tp1wFW+z7YBMSY4cVF
aVxTRRk3gJ8FKu+Lij0N7W783ZkZbmx0Tlx1cQ//DG9owkoxrkHvnm2WeR59ekoz
ZSQzwq0DZd5boqiVGLOO8ZwpiFJ/2mC01N7t9W+NSiO0oVt+ohSddYGsl7MeBEkW
O1xxnpBn3PfJC5v6DM/1ircSy7YSetHVGxalUdtrL4OrheIh4lcrUQH/8n6cSzdz
NR5jozOiN0EaTNzM0dbzawLJbbw7JS5JiohtIdmhVDXW0vpKGgM5jM+SWkaKjKm+
GL8CoS4F0xi0vD/e/vu+W83t1LfU4uvJAp97jQUOLoeqK/P8+RcdCQOmm7l7m2k1
zJiHKRKIHrsdaECSNDTgU3LdXp1vRiU49UMxgmYXgXEBNnGDag+13jugkbPmbhAw
bGGoZmL/14QbXydiyfuFs48kX2eG/VWTJbYXqSef8/Trs9ekmPYL0uVVIwQKaCSI
CNoeLvhcTtxtEiRUWPIdssFi4eREu8ltTVRiuDZ8ad3HH1Zb0KwiB07Z1kEImn6B
MMvec1vDNz+GYMsQ075FP+32Z1RR3elXy+F/oma45SJ9GNPBSAP9BXlEOIpKvLug
19kfX7VmivoxEjRh8PJZpQtSR+lNzWHupYtiqoRoxtalfhIeLZXmu3Iape10KpIe
1+XZRFeBYFTrI5Tw1X+iQVCGnnypvY6Tx5tA6dEWs7wPFGNDjUjMKe5aCOFqlY4s
WNo9QQPbbq0Gy3qBKco+i88G/8h2LvUGCEJ3Zwnz82YM63tvIri5gwByPtiYg5GA
QvBrj1rxjMd2LBw7LjVI/H15Cf4og0fkjD6FEQmsenMmRHJnWmw6DEH9vNIUJ42X
C85Q1crtsDoA1ipPxtZDNmq1h9vTUDSNYMbpK+9J7Ee0HbhpvZHeuG9Nc77eokLm
SaqrnB3UgdtD39vVj9wXbdmAk+GK05K6UhosRy2dVrSK7NUDoLE0ULQLSzs64Gqh
MOKzWPnBdBZmnpeCiQUB+549c3v7eZ/y0NqIZWddr9TDIneDBTkdMFNFxwe6enF8
FJsGafwtP4Ncz1fcVcj42ojCahcFora+qHsC8KbViOqnW4P6+2tdx6cscAH5RUqG
Dlk3MUQrHY9Y7VUc4IANPlSnvpp92XDQXO9p1q33dwlCcGsQLaUP/QRIONuu5IDh
gqQFW5Ee7XBC1enkkymic80gLRtB/2uZAv3MIH9lGWoDlm1Fq3OAYSz5z2MFAZeo
JmHXuaV/XxqLy22xlbTZXijdXmJ1Zn/wgPzM3q2m3DvqJjib21Q1viho9D7igrKf
IHUxMTGePrH2Om1haRkdoj5DbhMcMHyGW8Jw5qge07Eo3je46mYr50RQTiq6xzc3
8c9L1d4ieCHIlXiFVzKoAOcXy6wQCQ7XIk85ndtxHbsXHVviLb5zvHel+g9bcjOj
WO8UZLpHCGTlbgzypFmmTGY3+1OHQwUN2I1t1GLw/eZ7o7pAO1ZTiFNFyT7qe+2E
L+HkYtu6YJO5kBq221kFBO6ocnzvI2U9Z4RgIZNN2E0GDFIMEMx+DF69LNZN/90L
iq+cCX316xYfzeXZpGt05F1lEh002ascqHlVk9vyfMxSBxBVZo78KURMery/2ZES
7IfyeDEleA0C9gfIbx/97bmL64J42vIJHUWVr0rpDVjRI7XBwoIsdmpOmgcHIs+h
pv0FPMWw0Gxg0chMdsdIxyS06arl/KHW4gK+8OPI8050vQz/xo/Pe9KjJ3kAFXdX
Z3SR889CbsTtDZ1NPn1j/36/nF32trTUjCQGmjs7dKENtSvk6+M1Data3GuGLYM9
TGE+rwkTxhlxjCXBSyRiRsq+vN0A+RHOjsmlAcu5bT+XJiMfU9Ntno6/ASTUa/uW
Sznek/khsyqBTv4j7QWQnKdIZu1U2/hfPyqFfWbQPatFFW7K9LhyzIiOaO+TlXfy
FebgcEStqxG5vmJr+P+JsSQNxtny3S8q6apzu9or3AI4KYJbVDwEZziWpc8ED04l
FirEYka80Q7LfFrhEaKynBAKpqJZpAjaF8KaC2DV5gvX2z4Qn4AqnAJV8ilNZT4F
gwHZm/P4XlvUo/ccvBkKyZuK9+SYQ9NLAx7EPXA09eRUJG4UMmM320taYSNfIjo3
eBOX20cS1hct644ibwLvBd4n2b5GBVIAvzYZcgKl5vf9dBqAn4iswT/Zc+zIu699
IMDEk7Reqgrr5OirTmonx2wgo8mmr+q3Ujum26sd90Rdo4U3VdKIYhHQ6je+BbZP
TwcLhzxEbYTF695dD78CsMAY047jhVqXXIf+xgVeCoPraBjW+9bukieEytC4CVyt
3n+77MN2zpKLPhGkmNNQ8Md1C6NebBtDp3N6I5DqDd3P1e+N13qaihFW65ZWfsoS
+CDGhKK6iRCGAseKhJt36epAmoVz1QQmGtqsJ+1iKYWbojEy57Y8F5it/ngBTq/2
qSnDp5JMgEwVos5gYFO1py3wg2hkpq7RNrwwGEWLZdoGEJCeJ7b41qjrEJl/evjB
tr0qwE0my2gP6LDXbIJgUQxNOo5EUnszNmIYZKuxMsOlKchrYmNiUZBswwF7G8/P
lv3flxLLXs740JmoAhhFzUxA66Ajhl95sUhKskun40fJBsDXYMob5DYlaKbwheZI
giHGRtAtLrQxF5JENtbp6HyLHgd7mph9oD969tN5hyj3TF5lGB1gRxOvpNGy9pVm
xrqG11W1eP206ZUYGL7LIW8BMoK794XfM3TrKMd5WgINu4E9HJRg31V5JvIeSgcn
xAY8hNUTyVq6CYVphH8Qwx0jj5cVizi/QkE2tUdaDYSFbnNPbM0nF0oz6pR6WuUX
BFnjQ3bMISbJFrPuPVfFcpCwxp7PCaNPTJy+tIMNpt0Xk+3IGGKmGf4/AOZU8q1s
NSo8Ib1CWWUdHa6QtiLgkupa3XLG07W1m3/dgHgUf93O2uEx+KueEjlftIL9pNFA
vC3kAxcUsUwp68aN5vlm54HGOOTWkMwnKXiuC86buQfNn+qqg/KIppdqB/MBuCm0
9rmBBT4xpDy171w/PTES9sCPB8X95o+6g2NPmovpDQkK30sRqP8sCtBoFNASOlW2
JyMmTY3QwGe6M7cAUj+N08NHFWztcWrzHVOOPTietOVM5bcs3W1gyhCLSyT8n6i4
Pckm7yw5b3vczvtFeo7paF822myzLvcFWqQ/jszi2VI2KRsD9gUuExOZl9YWQJii
43fEjYOijIE3XZpKpcsJDtSooCqvIoUs7HNGRHdVebFAQGk1CyCgJGrPRL6S/Nl1
wjymTxlC/LigYnQTqAqQheQ3hYh/43Yie2U+Fd87W96ahazAQzKlCmJVK4LDncrQ
GiwEF/itlhw6WfflhOQgwUCYGAFlYkfHuhkgazy/Os7KoZnICAZJYX6xT2EvfKKd
5w1QR8JclBJeyJVtMr51xbfXJhmHrrxqjHjbXdieWkogkBOnxun6KfXNm6QM4Enn
Rgx1XUXeErODCd5gcPschqHO77EQt5x0j5dYXeJ9RDhubrYXCPTlZAqYX1ax7vs9
jHmmKuYHFRyK0fPFJIylIVfRn5V5fB0kMpuC5DkZIRF4fd2hPkRSF/y/fwVjpGYs
p8I+4ew65OAcB8WESt5Y2VxpRvTBlK+Mk8tzUZak2JgChHrfcuqcq0ZmsC4Yb0t6
EMUn31lUZULZE607LNzVR91p5cA+wVyxcMz9bj8gfxKRRhuns4cPi7ZIzYWfNcpu
CxtEIYdKrHRY4vd8rNnzTQIpr+JmNqzO9C42YoYnareNXHXYdyKipIqyPFtKQ0xX
+77zgArAohNj4MgVPnzqn9Q4fkshoozW0Fwwj8VxsqrEkH99EjjSDeaYQO8ShEBu
ImDaoko0555Rvc4q2KIvJXPbRhvXom/GRGcVBoPVj1uHlivnHdVCTDIE8/JfE97a
S8lyo5TpezSsxKtRdlKqQYV/Yc3yRc9wD+xVic700KRQAMHAmG3BEgbwj/vPCuqH
lJT/sYSVOrCGj9SpnL/sqPbPm9z9b+Y2CDvVnpq2OZJrMREzLKvKtQLUS/TKJWtK
UPJPqcpYWie+JWJH5S01rSDclEFG5G7DzyDU1Ud3mtuXYdOw5zPKuGvXBYuy4pBH
ux+ad4/OWvEGQJuurXOdzZXbjUgfwmleTpJm4PCcCooKgAqjvwnUIxFJXljYiBPx
8BI/3vItksBDZBMsvD1WBqOWELkdjC+HaTmVszzYC37grNzjfaGCq87WoTk44ydC
hpivaZVW2kOlxoHms5c7WQCLzeuuitEBeWY6jm7RaJYyUXjUDCFPAVj1VBaxKNmi
OpGQq46JAdbpo6YSXNMSizevaJdjKTCnose04nQ7pVfofUzZ1vo2g4uWM2Q/eLio
hdaO+kIcjQTeBnoGQl1IAPF2VTGzbKp9TAKRRhgZ/l4DaAja+fmcPayj54U1mnGy
/8L0ba/2Zw/jQ14KLOEjHKRqEjP65LQ/kYTZRWXyzt3jmwZ9lIEO/Sago4OUoBEd
xvg5yRc+aRWrkp8kQEAWkgPSyltATlAC2AEOAfRhPkaWsqLByMzmTnu+nwgq0bDm
Pw242BQJht6iY1UOzZLhUTdJHEq5x34Lo0qxXuHnlIY2LwdRJ2vDkHV+TgjwHeOU
VAph0RlsnXKhGfczFPoIxSJJ+62g9mEKtEmS0s/ui+hr5eewmH0PY5Rg/ezuZduZ
aHw90XeznADv4jW3n8/FamuBNzINFjJgg1zpyLzbLyjHTPsaCuw26CKYQZfvJ2pB
jrF/8Iy+Mw12wnXTFr5RM7GK1fsWFAWgqWV7Ld7Ccv8rtSJC023Ht11JFfW5pvRZ
D6DSJWW/XSQwvKsShSxh+moKZFqvFQZ7Q6mqIUO3IHXPAQu66SoVRHfiSxOnYOHN
OYX7MY+GZ8oRFfx7lx6LyRdbW1WVuwZAbaFRP9LGslgg3S29oVV5HQjlxc3rSsJ+
uJrcLill74cVTeMDw/7x7CTxx9qnPc5wNnUB1fp9OMdaaESVp5XLpr5a+dUcB1a1
LFM36aOq+/UAnm7w+U9bdSKDCRAdJxgsq/hmDkqClPSllgOkPpRj5xzUYiK5aCEO
6qRf5rqQOy3iP+l+ur3uD6wYdUev8sv1McRdDJUUeor0nOsLpDPwhOHNUGz4HhyC
pIcqAKN6grp8eg8w5Y0lbIt/J33q4poybGq8ekRrrlutuojWO2HIfxT4LYRODFKM
3hmb+XRi64IBMdTV0YJzp5UXxl7KgLultRG8WLSiycGCyBwKgAvtXT89PW+r49Ze
ApvgyM4H0GkyWd1DWg7wpgkuRARHbjfIIqhY+0/DGml4d8MwI01kKyKLiXKJZPD6
xrlTEnBXgfQaPEf39QpJHyK7/OFeJ0WSoABNbmSPyz+L5BMWNiYO1eAH5DrU5b0U
XdOHP1I5TLl1/MPTAPh9ro9a+HYFUS0og/EOQz/3Topf2aqnGpOlBLuRceajUTA4
WHL63SYnGZrSrQzPvQg9Iq9eQQ5xGVC68WOb/hM/ufC9nUVFHuO29XutKcyZASFJ
YjbmWOX7riDXVjnGmlAlxoc3qFyFmrsPXtW4GT97qBBE/olQvJ7CsAyI87TzpF+y
ay15sd8MgVLx9vRdyHGF8BT3Q5tltDuuDeDDch+zbz01WjtK8hA3EjRt2vgHsT3F
EyiHNrNZJUyI9wR/SG3GA4u6eCg4beeZ56pd0eLGp58lYyeztejWz07ug/a1LHOs
ZjPs8aiZqwpgkFnhHmOAjzlGA1f+SB6oMEXeUhPWEXkMpkWawwq7Aua9UICcqi9U
jteRwAVxltmnha6ZDUhkg2RxuvO4CoYt+bl65bdztVBnReQDru8OX7GECRoHFink
omQuiOqCQrTKxUJGK619qHta0cnaBNq4U9zlRdi2kANFyp84fmcsi+Zw8f6zQLfo
nAM8mXKn8KTuQbp2tI8AwXcBOfOiHoWCVaMVIEoIBFpfA1M5AgDfhZ/DKIkBlrSY
osvL/UJRivHhTK7Xd4fFz0mDVxuTFLrkAQcFdFd1IF+f+OYjUXKzQtXA8Mm9eOi5
gm7UFFE/PQjOofLLO7YIeacMfCMEiYaP/PSPWAc5d1vaJrH2aWr9OQXkkO0LfPcW
KqBWv9Q9V/7G3LDNMiWVFFT/BMEqsC2L2ShQArzXS+fqySponiUzScJoFUPwW2Kl
uUz6+hVQJJ7x6tQj1lgUvxfccSo+SgPbWCkQ8vLvqIblLJ0QiT6lKC2boxPaI3x5
gAN2UJBVz5FKp4VMQ9uG9lVmEjvGnU6QS165FAZ+Izoghzp6L8rltutg72Bz+Xrl
gWZSODRrreZWPJlDqR0JV3lSTGxNID74LPh1HMKrxKjQVXb2VljPJ2PUFD1Wyk6a
tbvOdnjXkezPWzIdB6AmK0usEIcUOZ5G4NhIcnp4JuduKrGaPXgXt30lqXRB5OSO
8L0d1OjZH0Y3gOtvl7CXt6RhHdkksJXRW4wCPKhCDrX+bDetzy4i7w8DFPaSAKXq
VdwYMzuOaNQS04IYXed5gffNIPgWKhLiuYgTzhF8nTjWrzhZonSiWNesNyCicMYm
/Nv55yQaJkhpU4lwYMW7OmqBJcdP7kZKdhpxc7c5soV7fFN8DW3GYrPCRxAWcE32
r4PainNRGvXTOlMy064B6WkdF74A689pe8kueV4oiwiJNv0C7ZQFDgKRuaN9l7Sl
QrdGGuMGkQKnyQfn7PKfZ36Pro5ioanZsDPsz3ZHssY8EAz1vw9Jus/KK2LlADdV
usWoFJQNSPADI4Kzwd7Ddbu9zsus4EZDrhkbtGAhYiWfnMEOFIQD53j7aaERNFKH
xNFZ/MBTYvrAVjAxz1uLaGlKXCGQsRnbspJlIEVeA2ea6wx3GpLS1V4DkCycRB+X
d4O2RP63EKrovptCV5GTKnSDWpUGLZEY9NIMQGAmL8yoQ08YPIWIAXN+6tPTTjRg
06WJOUycHIVKXES0Yh2yJGjSg6xtmY76QLwv8wyumHjvL0r5fKbysxFSe+ljJTlZ
iQZbaSaoA8whAyllQ6/qvtkPpSE6lH3XwZ/ublHiUsTzxKsjzcYVpTVlBwrhGnK3
J05Jl6eRq2038RX3G5BaYfshaxecFkwpvdpXtNLOKIo0ESttXnjRP7O2OqvypuXV
RxVliC52swn/k/IXTwz7sOxm+a+cpUj3yyvKQ1GhrR86/6uRZmnKCwZSMbxpHfAb
pHE+ms/vRtmT1npxUGZBoK5gRqZzayJ8YLZAL4idkpnvpFTZLJuJYf1N4O99wcmG
3hJPW0i0cPhQDfUDIca9mYRpephNSVhfsgu2XiBQjx9k4bh6m/7pBAkAj6W4yqVj
LuQJsiMw6baQCwLD8s1noHvcMUBNuGb2x7pdS5JCKS7OEnzpnO1wyXCpxxYXmb5g
A6ddRkC29NvwfOYHUjGyrtWdtiIUjx3vydzaP9t5Rdggjk/UuTIjCE1XWFWPkG2h
gsYE+tswMy7I0TE3vZXWIuLMSthlCz6JcD44482QFs8ZxPF103uytKMveNL7+cVD
osfM4o1cYoaWQOc4mQ1XGTgGspkrMqle8X4yvV8QKbt124xIsS8PuK/bqYkETU/h
SH9MAvq6rt69WVLg3niO+2zMLG3JJjPwcZ2z1ni+P/+fLVqcDsrsHmYlvnzETdxS
rUjpYJyMMGfuzw7peF+IU05Xg5LBc1hArlcX+y/YBr4A3EK4tBm75WnLuGfYeRT6
2XVi4Yr51EPDV+Yh3Qr+YcZJHPEd6i8TPuftNxJd5KpvIdfjDqFKnAOaU2+Tx2x8
f8T6QQMnU5TgSABSmvVESv7XPTqvRP293c5kiphYB1gDb7Fh2GuroBuElIWgQUOK
AtBODLPG071sH1bbWbSgPsVjMSUfmdG/6OrFjrKw9mB9BghOfXA7HQp/+bwkyrHz
nObCJkwyk17bt1TJH06oQ/aJZ0mKFpPhMhzSochkhTlzavICCu3plgBTz0T17Z4M
Y9pAAB82aMLkJlxieY1ifpMxuyQAWQ4wDFckzdPudM1FlFFlXI06XaZiVnq2ueaB
8VGT/5qlEvJmTs6aqlSUJ0oNYnEM1uyPcF3jMQkj0KRtAHV4lMDwtSCnb9PIkjGo
uFoT6eRGJYtnvE5pTprmiETNDQHfqM0n+tvgX5K+tBHqqjMyr+2XTplP55BAZv7z
fsn/sKFTZaJgNkfhO5WjFlDEupEIvIuO2EdZ/eAEV1/WTuVzphi1DADXBaUgqjFS
V7rZns2x2y3F4y7FL/Kom9G4/41Oanh1AzjlZBB/BaDYmj+ZvSjygO1UISeo+b4I
Q84qWoNc0Mk2RjJKF4FZc+UL7DZOBlWzoiu6uYkjf3bd85hP8IH4qmylJkugVMTO
S/nptMNxHI0iLUaZAXe0SH5TDqG94YwpcpjEgQzNUh3pNEzAplTK1MjIWEC0rg8s
qSMASr/oac4hP5KmCwNtJaTTEO+6iYVrifBcdWi4LljdY0UV8WI4nl79llikAqvO
xtqobzzUo44oTU32RGQSH+cpuhAE6P75aU0rsGXeLknQT1BUIFfR5UFh/54JxSfJ
Rcv4w8Elz7LI80Z3eo6WvVMLuZ4nlJpTESO+nE6HOLtyABCDqAdNkPTZPgcKg31e
/FnNnlY/jSDNo+QSVRhmONkx5zbputfYzCKgJ498+eB7IquPiJ7NaEXfP9pDZ/yh
jkPzn6lOyizKN8/G+/gfjNaEfjspWrUcZK4wCm0tTFREMg2eOHCu8tm8ma54zlXq
6L1ldNaEQeWrLWf7gmNeClV53Fb/mi1cBCglo6qXbOobAGLBlNCdqbT0Gb63vCfx
H10c2D2e2NorvDNpIkVp9IcYhKkDLewhOEeLOg2SO+ZbebJTrPMVaCa/mAF2WfLj
TqQde8CQW/Of+dckaoZXMG0SQh3oGYDIci1FHoV/jH5Wa0cff3yi/Ad6Qf1MnrkC
6GrZbstrX2YKk0yozhL/A/E06rbfcot7sKrTBm1oOa+lOVCsxz475JcB7uZFKwQR
HkZFnTru+QjLtXmYgDcT4s5/ovnApYCOGd1wvdyXJuWpgtcevEt6z3YohT/Xvgmm
kcURPvgfqyfIWBxZE2sprOjubFqL+ZbuGjnHkiITGRwMvbHBZ9qpT8jGoyUn7tz9
DHH3tYRS2r0NA9iv/TvgOl7FijsXq55CvoFcBmF9Yp91kERhzLTiuyoOFxxe+9A5
krlgJBBrOtFrqxYSWzmPsOkk65cW+YE/aKO25ycOOCPUtONrMXHuaHIva43LZhlU
01oi1HNZuuDpTBxgRkKSSxqHAJB1GAeO/nZv8kdigkOUwIMhWykqsbk5wO82wXdQ
z1Q0f4xxxqUHVbz3zz/ZLvbkX0H455Mdk7XQzDZ0Ik9DkXfvW54iLbatiLB7p+06
7lbutONQo7PESQlSY4XHAcDZEWI5kYinWkJmkeY8c4giGR8l50AUvPQsvsdLVOzp
H+Lhu0i55YjKGGNrYjyTsoW/muaBZp82SXyrdsodgl86Eebyj8p3t/BqZBErjTZ4
PYGNV5XRvdp0GXhItidkrs70GeI6B2Uh8rKBQLz/jl+PmNYyTx35lrM2VhULbvlN
7EbApId1NIHewJXCyHHD+U/Sw9BNpdY6tGiKoAv8IiLGxuG51phPGZ/cdh0Ul766
3PGzrIJ8VIE/4BQybmcqJTH8whpaFd3GZL2qTU9jKiQeoz6ZVMF9Tr6L7eX+syby
frM2p6cx3qjwjkkTuNuaOC1r/J4qQ9V4LyXpwwBEFlSvCUCTXIDWjNToCDvWjtVK
Q8bcxieLbi+EWJxIpO+XZWCWYeXiCJjnIsmjI0Ni6shucnD5+O0M877PNOjotnY3
XI3KkeHMOzI0WBEXN0BG2g4fKAaLsxf29SUlB4zP8go9iZwpYsIKj2zpfPWZnADO
CookJUN3vs0I+1tsqlpp0YsW9P6KDxgIV6Q7S1ZBbWPAqcMj82r79u4qjSBzIA2B
w08eMfZTVh/6dihE/82231MUEaKs/EHskM3oFISiWCLCf741ayl3a/71h2tbcQs3
YKDEy6hk4QywbQDQ5GWTN32tPG7tsJnVNgMKkcemKfP6J3MCqFR2XM0oVDR1WpIJ
7kIsCm8E3EsiT229ckB8ODD5ArvjsoO+bHKbxldPUIsSNsgPap0K0CTROhWQUkAm
6ztq+HL475NFDB16mvDw/W2eC2AmTajKdExPgH6MBUt/wJClTSaVl1V1x+/toY+y
4MJC6lm1HGHns4RIVyL0mvzi6byJkbbOSdQ4I0uAhZP5souFvFHAeuuSWKzcFPdH
byKqiB1wP3fyO/SG7znvFqeuBdJhqarNB+YXqYYoW1XWxj0xIjq6NHLpruDi698S
tLaOrUTxMF7v/ogRM6EmUyPfy85meNduSLCcfHAILKRBm+3fxDdBnKZGtISpSkhP
TziOe76kORbzP2ui8IyJR00c2TTsBAPoASmSGxAsf+iRHwM5MPmXtTw85MM3hIkF
kGSjSMMgBOSNZ0feTPpGRdN9V2/yTa4Jg5ASSuBd6UKws8Cez5NETkpAY7+cWv75
5NMw8k46i8R1gQwnvRFwCGu3ZTnsGZ0vlbFCu7DCWVsDO1CWNO9gPbz62haXRXVy
q/ZzcF3zUSzkD9nHWfQt44L1thYK6DCJp3RJ5l0Yp3w5yImNQ77L473y6IHncUra
5EHS+e56Tx5UDxPwkwabLWYWmkEAjjGxdTfAwuLTwPA4omFm2ZOjf3TeGUIjpuox
oKjNwcmAKWXvQm3Ttlim79Qix9H2u/JgeolAB0w8faojH5yz28fSEds/TH2IA7Bj
2agq+gpKVr2vZTsOF/6KZItqNt/J5jW22LVuJSxSetPt2Dk3xfknEXs19yTeCCFp
sXy7QAhA21yd/fN7srnePMWfRIRvvVXn8/ME4W3lXOLkDed9t9B1Gz6l2HoGbB29
zEMDPwmyPT+znn4NhI2Xu8lbqjTM4icIiWyN3vWPg2gCxNYaaATB5Z+3RthW4JSm
xffRhtcwlPiHIgrzthRyZTLWH+h1OblNxghxk4Kb3lagBzSxk63c0kU4q1YLDcjN
Xrz5UPP/NXmiWNoHZKqtwPsRsCVwJ0PD/XPswBmXjD3/A6xjBdKc5BfOvXhWufHB
0OrLsFCV0y2K+7Kx7aFcqhKulNogIJZ1U1Dlg97utIE758vbaYotKk+aLpQ1L2Ey
STdu6+aNW+83BJUW0K5Uf32QCG3RFBBggpAXMmZmVbYXDXdBhKmhWgO+7R1/5op2
7AcqJ/2LoVncqBliY/HF8p1xFUJ4HUE9vD0NDWoebYPFuFoDrdKC9feD1925vock
ctGGhGoM62NNzM07DMibHPReULSZ1RuMk7m2VQE9NzPcnJYmn+QX4Jt/1GP/u7DN
LCG87CONr/X9eLQdvHqYiVfPOHC/QiP7WZK2KvCTpObMzs9NPNB2E260xzW3VY8H
2qeiJM5Z1QJ/qy9g4GhoiGJep0BZehoOtTubxwJJLg50SWe3Vh0Ru+ZS0Qd27irI
/ai5SFSYQ9pb5akxm/UOd1jFxojLRPCsfGjRcGsBjYuunyNWMsy0dKRtadD6gw35
1GbfAJhDh/0Sx3+XcWOE4qtOkPyzcGhT+9Uvt86U5xBynIqCt+Q/5DJwvxavZ32u
puO46E8U3xAjfqRHZeLBZB+EpkGE0nJc5zpUOjR9Oz203/O/usP5UYNoe2pxZU5o
cEPKaMhw0pWei8Sw6cpiW4goBCLa4rZkuNirJOSq5LqCgg7BOtmDloBB63e6Oq9z
A8euT5kg8jbCJEFrVy5kzDUeWmRdT7mndayBp+AssMJwjnShQkH37ZS/6OJHbN8I
ZkxAXYeQOefkQA2rGPiOP1FTGyDdUTD7g7dsi0UBJUDfrfqhH9swibq9havX5O3r
8wBYE/XhyA1/4u/vvNMFv38Cx6kbpT/kDeUEUBRiTmZ04iYfhY8Bn4JjOQaIm8pD
e7pv1okKcVZUJuWvVyCBQoaddQFBfo6v2puZRuXymz9FY3luHj+iGeS2+QkMs541
rtxohZgutfbZkz9H523oC+gTLoCcuTGOoB4Q0DJhS+d6Lv+E2L6IrxQGl5ovnjFl
xRtNPZhw3fmsxJPrTliLDLAQ6xE9bA4KgROwvOCfObXxfJR4iwTqGhzFct7Z7b3J
yO1P65j7fsDE/2xB1rKJDEwZAOneixQtRPRju1qXK6YwPOuMh/eo3LrXcKVFpPIE
XP9aMprxsZ5H1lFds6Dli6eCzCxu67pPmwWtByLVdFqJ+vArHtx0cahBGNntvYM0
QIjm3jxY/g4yzt/J4crShFqKtDfgL0eOpkGMEZju71vgUSjRM/gmU9QE4IopXkbR
eDpIg2gLXpISviIttzFJRJlfd7ayh3VRvK7c0Dstg5pzMdCpmOmAINFWzFHuTQtM
Ei+pIHmhpWdYn6qJ/l3t+Ta+fwt2O6hxGn9LjRffyAEjhe+zi1OnxCQDuiBk9Fr4
gQMRYDC6gKIUtRmiulPkhLt8pLTaKjqwcphGqHuNAF7Mukq7rQr9fktBdjPZl5FU
ay1dWKKEU5Ec/KVPG87iK1+UbQj/P5Fk3upgXzJaJrvKvzVuYE0L9bcJS5v6V/0l
50Aa13MPw0gSxX1/dXnuTmDlPmADToNsVd+2GmEsGJRus4RehpX+SveZ4Pwdb4mC
BRFnVbuXmbjEtamtb4G2Iz7ZtIex4J8Md6ATy0vj207uXsW8fYQtLznb3dNTTe01
K7dlAHA4+ys1e5Ix6S881Q/WzEIA1sqnn1a6iNzPIyliVX0kTZFBU4p1CKaxGXNT
Yev/ELCAbCwqUNog5/ZNoIeMDBl8z7OFI3K5QOdiXfymCgYav0f04Z9AUclMX/6W
2BTXoqdtk6zmwZ+upXmgV/Xl+syPxifTEXD6db67wvzEw2CwArszfKNAQi3OaFcX
XSsRNFlc4Fx/cNKwvvt3Tf7oua2Q6Nc6X/XV4ZXzs7i08kpjtFVw0LNU+Vx14R8D
7n2L3vWJvZB8bVTcwl3+H80pJPfWvT92Izbx2kJ0bTPi2oxgvnvaeu8pnopvi5IE
DSiZVjosXqchTYH5Ai2i6Ry554hl7inOYMUtp3QKVu4kfoKj7/WS/Vsl7VSQdgXC
jOvkA8iQKBkQC2xVsQ7KADifibKGXDZClNoHncbT+fC5QJov0GxC3CetN1fQw+Cv
ziLRWhgmrRfiQDyh+p9kfewT0vqKDTKPW/I6E6JxYfgXVoery34ZuDS9DvCX3eUD
ME9U1gjOWQyIfcYSDLSrK9TJdVbm8D227DVKxJ3w5DMkilHGsbyC5JFu/nWrruJi
4MLGo1xItvpc3BUgKlGfGUbM4XkwlQCjFusnI3jINCnr3vrxMF7rKolSzjpDBh36
Pj/rHAurTJENgWgErHRwUMtst+wrB4ZDDZIuw77xqUVm42NZUpExPjXQFh44VYnP
P3PMuaW9j5VvSrU15SEKsomyThGiyXwHrXvUo41VyNRqciVvvQdIu5eKjtYCd/Mt
vyk/rPfluCUO1+vNcskzTQ63k2jpgekcatuTKEBgqoLY4X6Y9j7XNNiRxD3jtaza
Jfctq0iH/FDIamZ9wBrmUEfqZQiZ0qMjZM6UDLpq44ZIrJilOEjWOwv5Zz/OaMqi
jwcWVB6RdBKHkIyuhtlWFnDF/L3/OBif1lpf1JjmTQC5rV+4RUfNoqx/28fzejHz
9zVcM5a54SB3E6Rh6VC3G94PTrM6w3cyCtJSTKTpHT/XPvk5MdtSF1cLvSmJsAtE
Oe3OxKE2YVdA+NXmxZ3VKNgBrD59bAT1TsL8LQXqquK0EMOwohn608HoPAar3wAA
L5WSOVYwsynj2wFb5B3rqtNqtqCb2V182o0edDVY5Tm8rVnhFvax/F9r7wxmtYLN
TBNtKZFunqybKheQcZGAuTcevaGQmv4U5QKW5SjAn4eiFjTaYMEXk4Seo1QrB6a/
1AUvdrEZBSwrK3Qz2aWGurMAuHbrKWdxwJvm89TE+uyy7uPKt98ecYgYZ6h0gJ3o
u+kDIDt6E4OmQqBrYbZ9AG/B2XZ5RXA/Wn2/MJ0XBl0/QFlUUVV2N+B754afEgVb
7Uu+zovKG4J2bayau8685o+XIESRb9GMmo28SXbVHlIhhVIWmi7r19LaR5iVP4Hq
DELN/0QWqcVLDnQONB7+Z0yj7fLK/eSM13Otnnbc8wRoXdtTBJvnJNJo7rYxeApW
hFOZTSXmRYfLmmsFqLytcrcVPExwYTbow6ezi5Ok1Dah4jE8fA5oCRKU7FKelQkF
gnuJ/Mt//s3WdFeDg40cWzwnmTyyErX5T0Wx3WoH371chWuo3JY7bTSvHjiVl1jY
okCkjLAhfKola1MeVG3I3C72cwIs6A65xl+QYEaFJ/wi9dLUtsxMCrPKRC7LCyTU
kCjS/UCu/rtd3MjJR8/2gYeOU70u59N9n6M4pUTJzs93qgBVQAOn2+sJXZTa1wic
9kaEp7CyquCB20UqwUcx0fVPOHHwZbAFVD1VzZc0hSwBz/xbEOGyIz+4976UIFdi
Ws6KhK98fXD7gCIJ8rSad0b3gul6hGyr6fI8lJIN7zN1TOsU/j79oGUH3xAr6hsn
sikUelB6mloVcMveX9J/Wl9TiPS97Dh+2YzkK4nvnikSTTDVYyHkBHqVQSRTjxsV
qxZAYWObXZ1m8RklAb0DSb2d/mFSz8yNOvuNrtvrlWhJLodu88EGf8Uh5/4FgE2q
pKBWQ4yLoQmUCNzjQZzrDGwtZN9s8nXt5gKjKBhXXxLE5lW0zyGbhlUDmGpv7UzD
QK8hWivvSRROt3f1AETB9V489OkFbcVqtTZMo8/AF36FVhBVGynsebqDmsJCghmm
J4LwrlbgsUKgS76Ht1pivw996Akr/Ti6DM+Q5c7QOmYfYnd6bIGeskzRAaG0moQV
8p51nBacERY6+udOJ4cOgmJWbMYEH+79SZQrLC663uPZL/LYl1mplojSdLiY/ANF
uS62EbKWb8KORVPhJKftO1jzYbxOpVA0XP1Im+izUasAVXsMlk2qh/Wsk/bdw2Sv
WDZ6ZvsnDkGkFwLp+lmf0I5XQuZvfwwmpx3H7LqF82PDxmCRs1r9R3WVIlMCLo4j
Zyz2eaYzfmUsQUl7JcEF9rtTKU/QHw4tz/ZqegNBPY3wpjKE9z5Jls9eLwnyMJTR
q2MAvF/nXTHjhfyNyg2kmVpiJdDrxoKMA+Bc6Ym0RVCXLkwxymoJ0yr0blXRqp69
QymTiLE7vjSQtI6/PVD4mO9vbuAkRVqaOOuN1QBPBxM0yqrNL6RPDhi2FeLnNpQp
gS0tD2za3e+yi05wK3QMD2nr8H2sRtoLOq1VEd+uRDm4IT3DxiF5tzGAlez19nYz
/oSUPcLYwxdDUj4IDBcKpcSaE8GPn1vUOSOMK724zX2q6M6Nb/y4IWiJ75nfYmF/
C9yEXY3WJ4OXq293LHWa7aml9g3G0DGI3+g1uiWDJci5+QJ2o4OoB1kiCA3tXdOY
APzcePC59uSuT8ruzrWho29oc0VYXOxH9cSG2c9AiYzZvx/415Js8rq1QzvYD8WO
Zdgy4o+v6oApXqJ2tPBhKyxCCFzENJqY4kOw0NFTxxl7pv9yeL/BXnz+hkazAaTU
ajmdVQNu/pL49tXuAS2s9EqADORcL85DiCCpkMJAiXA4KuIU8CP18RRXn1YfuO0e
42p7d4p7/CWROxniwFk0cf2nc3bJpR5ZnE0IW2Smr/vaKbLS8D2WCELGvsdpgrct
swQwS/tm5VcVXXX8rTcKkBOvZoCYLW/jyoxFFY8NstJRb1FsXXG7MAIP8Rm3JvH2
27x5riYNcCV3qIHjV1VQtB2VPYznW8UDYnxEnp3kET6XZR9Sovebp2O4vs4Js9Dd
E9FE0NS+rf8rqsmq4fh527xEQcI9P5AjkICfFXDqIdCLvUf5tL7iu5vngefzb3Zk
FNY0ZGeC1wJ3aeQCoPxbJuouPgQHOW3Iu+r7zIPmGQepUVkLNejUd5aflFyFuYUm
mdV3VQGWOa6RYlHfxvlnphc7FWp/ZZaxkILYyi2kmXBWpMfi9VaQ1pdUB4ATHsI7
UYWwyLBCWN9zkdZF1ICNDUMUwc4JUEXXJrO5XTpklvjHPV9RwyqPa++1ffe1ZqEE
5S+cJiLujvPUgxfyVtBkawH9/oOtYmYX3y+QbBW4S0ckVgFq1XgeAvOeSEVGS1jD
9CQHxglUYxwRD/yxEHzUV2Aq4LJoQlGB9ER7yePJeuDFANOPlObB8T0idda6lxND
yPR0kMKYwkHsSx+Wjuyfhj+/3CFw5+nb1MxOLswXO7/XcrigeZU56n43B2mAoXpx
XkdTNx4nHiO2o68zj43aWsrdiDLZys7p1x4gNMeCpSMwAXi/x3hs+IIg0QDwz83Y
+xFqwg4cUnxZ97WUqVoinRHfzRdVEg3onPyZi0svMBh96842U8u7HEjjJxf3Sdyk
a3hJxifNyTsec5/S+6TncGVmsQQU5Xz8Mtdef3/L398BfaUBf0bU63NQ6sm82CWO
XSDaQmQ2Izx48yrxtVF8rBP/oxTZ+PwijE24O16Raz0xr6aPUYyYrIqdKNOx+jj/
5xKaVf9bBlhf0Z08GhsNUOJdlajhx4KuX0c0v6zQv1+/DRhT/yZfAYrqcvXl29Pd
gqb1Yrzj5RuWqVG+tjq9JcbE4w0CeycNqiyYx6EME3udWi1yreQ/N06d17L1zzYn
R/I2y+BUxi++JzBQ/tsacNpewBGLhCF63xlPLX9jcOTdSBh2iEV19En71eYJ3ipi
2ArPIp8kHBkUcicEw/t41MeHJUTmuNoBuYMOFlqkQS3bNHdUk4btpd5p/SmZqoHh
f5mKa+OG4KNP/FXJ6eEclqEEUajgHNnNYC0qYijuopTU8P68FuKF8AnOf7y+Cv7Q
D48JN4xE9dPk4SVknQf5/UR398mHNwo+9vmea6J2jxuwLVm0xf1HBVrjjLr40VNb
7hjZQhUggKLH6VEsyZqKWj+3FvOykNK81gHC3Mptf2qaEFAc4NegthHdgZ4LZRyb
s/pDCCRFYS23xc4gyH20BE65AxDZNIsBYDN5Y8VMwkdk5eoB9nj3Lf27XPF4J4fc
RCKHcj0PwfzIWyaHojS8mSxqr3ZmoiOIzg5R9zDt+bj3QHsN3A0vfMv38crAThVN
eewH2ZqMgOF9vulpKaKXCCug46gxWhcvlbrP8yCVTpzvvbb83N8YoA9gJiQhp/0P
nTwJ5cnpl5CsT7AJFF9nMTWU3YUyqEvvxxHjapShcnXtsCfP5RE50B1Us8l1f9Zc
aCIdrLoPMYRO8tCuWZPO07UoJ6Yx33/5juNri22e8v/DvmkVHbajPVbEt11PnCZk
GB/g48Jbvh9L1dmJ2WJFId/qojBzKzVl79LiXTMSRu3QP8Gc7mRzL/PYp/wLrs2v
WPr+juAPwHSFtUxbghwkGmdkWrUiIBoLn02TgQfxGAHtKg5616S/ji8nDyYdDTKV
oGQptONXgwTxglhnadzv7PbbwAl/l3kMsc8Oy3OyxYOsPpNbkeBiq6MLD1LU5TW0
04B1FZU74QEhUb6FF6mY4uG7lwOAkusNNHEvj1RBp1EDm0QHsJx+YvsHvQNzWJvQ
C/6BTP9gZS4TH6lcVG7QYfD0UUvL2n6QTcXSkhOpodHfLs6VtbE1hSNlsDV7pCkQ
35Um423vrfOv9mrWm1PKhg8sKRPeaQcUxMU6dIrw3Mb0mODk0DpoNHlaLJY+qpe+
RkDQHKU6dcgt6+ntb37puM1LyXhIlKoAgkb+QMGn6XJvsu3OJNHJS6zyWd6+HHZU
Jy3vyO5MP2cRT5vqu+Duayz+ipCYwk7TCzLjt6TfS5b1MHZMD9sPxLvVTYFFCrY6
0ay4b2Y3whJoBJSm+vLdQCZ15UnOPTLt+e5945HvGBkxd3EYQPDFKHEB9TXmXDRv
/bicKfV9HV+9oj+AZQqPuMvVC8e0/jBeu4hmtY3du2ta241BV6B9uAwQxXoxwhjJ
zxnKt6l+vWM8BVEPPt5JjFQzCKEV0mT6qwW8k2mKwHKycYxl1a1Ky7Btx9sJz/jC
VVVpCIPV5uvZRiFE0Ha4TgImYleQwtfP0Fe200dbvh1XJPTazxo6mavAfAnxOmzl
dhgd3YrO/I2axmx4M/3iPYeXdSofLGE1EsrLvsrPJ6pmUo8D4FqQdGdv7wNpxiqU
jKTKC25W9vtgiUU7iG+QvIOUO3Vra7i/1YuoxfjxDvsFamOknfhAWONFCVbcaR2L
lxTFFUqak+qH3Tx5RQZEN0n01FOs9jUG4U5Fx1o4+4p5NmDI3+huqLcjuJOy50j6
2AgfU3UW5ttBhlbvL6RtT+Czls6jQ0UZOWHWS2v5j8i3irK/k+EWQJkgTclpauGS
m6/0m5zGKLjmC3MlcToiMBx/jJnERQDSMEokdHfiUbgEXsYc+zOQioNU/KxvTcKW
l51kVCcjjYvier7zZyLzIrN7O2Ngxfv+Aca9k9nYV0JSn1ZcfslLGMmdVs4xhtfv
pu0G1b3osLDwQCsQQMqQ8UANXg35ZbMkgF3KVt5LMSo3BTCnGbeNdxvwvNQzIAFl
b6EMm+is7JRVNseTpefiN41we3sX0VglIHfFe58AnREO6YwbgDFdxPsiAjx74w74
6VBB3bnwgEDRFKR3UJHRGuIUm8LMGRgjt3LQ/0Iij555wO3Nua1ig77Z6PNYJMgX
U1duWjLQsHLbwtDdR2rqCp+/RGHMp17X+GaTyGSfjke2Ohb0Opbec9cD5+TDPfet
EDaiKBrvwq6DFQum4aQlf0x8u5M448+Wz8KwnZ7SH16KLdZGJqV3a3d5MV9m9zlq
NxcKwXW8uOm3Ov/wfIRt0SZKiVKOZLAMU14WH6iyxIn89YTvn2X5yYPphwyu/bK1
NW9xJ0zSckmDNIjfvay5plp8CROkZcSJW7+S4KqEY+pixJJFoJBqfj7NPr2yk6Pt
+YSFNqbrWVv/TuYpYdX0O1p0VS3LdnAEa36adyvlzjFvIO9ZFppo6xPk0ew5wR8o
aDQAu8U1ZFC1//Rzga9drXaIkkb8CcwtANDIll+Ti2xyPQeByhFnwILscFuweYbR
7//t6i/4ETGKoX6bKgETL+MXxSj9CDCj0I+4YAM+pegR15Y1N+rhwJRg60km42UL
efhtpss26W6DodPL74pVOskb6ooVgWz95FxG+YYtzSXOcoivXo292OT11TMXB1C4
bzUl/jSpu3deukdsnttlWdRJBZmH0rYZC4kGOR0I5dQJ96sGdakVJy2Q3o0eMxie
EeVMwybSwejTvHvwcq+zE9mF71wEYuwac4GQz6JNnG/mpnk9xkGNNHpfvqtyKJYo
0S7HTGL/d5783zkDx5QnBknFgsJNYR0GnetCJw+83MLTcZf9nXwrQ2niuTwsgRhP
nS6W2Y29QBTy7wnlUuz4d2Zn/PDg8rDKBExdqA23FQpGR/5tJJfldMQ3JWwH2sZ1
zxtEJx0MWZu8QzhBPVlQWNTo/KPk3ezT5uIBXlB3GxdeTv0RCdG2LzkRTdtteSZg
XXXkzXYSI/m6djpKir2PvsrmhIzG2Fj8JzXCx+8I10wZOBwxI7mNrdWr5A4JM82J
Zk5WUQIEPqWrKPpB0yT5fOfX32+07K2BJ40FA0IZmguia5Th0CbZGflMVWpv2S/f
X5GIucxW6LxWm65UnW/zb4pYS6tVGBrPX1rXHZ3H+BjWwXPyVkx7hNT4rcCh741W
pS2XW9Ra3rMiLzTXosf8Fi1QUqnf84wdW5WlmM2Sodw1ykAOiwbgQGovxDk7rdkT
5XamgvZPsTTlQ3GWbWzu0fkbKI6w0WDH8j7gBfGu7O1mgKbeqo4tzegHyp8R5pd8
RvF8L5iGX6Co+CSDucHQbAc+nUSW+1m8lUstvTEDixa7QDMkeN45be63qftpkJza
9cFqZhLxFIGIK5NSB2YFB8lFx6YCDx0F3bkCCD3CzyiCrYDJ1aqkdA080sc3VZOQ
QnQ+cbYC4Mr21DBZrbflS+zUJRBUcAMSH+HlHS18iFTt0gRwV2yKK8fCMI/Xj7/3
mqsnRQueKU7LVJBNXQkBuzD2Wv1VGAs4LUK9V78V8lLzzYHom/IBIJ2yoANVE4JM
w00+OVX1y5F/nH6ouLuKi29w6OTHDq9CSURlaRFqpYeM0/8b+VGbXi6joHIOdqxZ
W0Zw7c7C2Ao9RR6613eiuz/7jlSmp5Uj9LhnphneVqRJAOxxh4TUzjo4mYyG6OgJ
gfP0oPC4QuSnvLr1GmMYFYje44aC3i790yK6JJXNPmugvn2k3Z/ydLuP/qS7cpb0
bWljYk3vb6E+lOyt9gBMf9FlDxthksx9FvS0WT9pEeE3wMK4zABBV2zcYm4BmAwa
OTK5rXhhlAUxePPwcCdMaH0YShGHeRpu7C1Y7t9Kg/Glz8G7FiYcJuOYOKC4Z7bP
Da68q89MbPNSP0aKjjBYJZvO4WgOfslO2kJFoNhLUsvqwDoF6xFUZbCyJRuW1vFo
c6eemE0A0onaWlXWdReD+ihTXvU1vDwe3I0MZdB2pCYFQIj5FpMTufqL4WoGCBad
l+lI6OZAkVlRlciid/Pkw6CLXEwGRSOwZwRWW4QXntjyNIEsMOFvc/W7FFNeEBGE
uq43oaZ9oNn058lEx7UCwCVTf0XVPlhz/aDFNfIqjaOnUpwadFFWTlLkzRVDJg0g
Z8492RKoCCvluWPNcR3OQ+r2e95HORa8yKgdE9QMpWReKRL8l3BiVgEoTIAnLmP3
5FpxI2CYCKc4RAyYl/gEYNJkTdoSCDX1Nb7cwjQirea6xkCCpfCdWptfq59WZhJH
73js5nEnP/Y0KE3GCflWhsoJ7635PvbcZ7WNC+eOC5HThDNQGJymkVkdKivNbn1w
DCb+G3Lzha69g5tKOpViYOo+SATYw9UH4QdkxOGIeJDc9otxIBdhFf92+5FFpNuf
XZbnteGRIwnOhJKnXDAHS3j/ztnWE0wUAeBeA4WQPSl65f40xs0UH7U04L+wPXPC
NJ+m8zwcWARrUDtnuizVeCu5idTFbx6bnVdVMov/kAja9nksz4fUGYC7h6HcrJpo
P9pca3cKSytepY5UBM67V4HwJ23gYWFQANJLoaQVJC6q9JGo406abL64jW9mXfBq
dWKqFRrYHd8MKqBq5om43KS6111jBjcN2hFTsp0XShPZwOq36qeswV8JfmNeUxs/
RQj070gnrCMN98zR+ehk2sbgYd8D5fd45UiN19499zRBdYN/vVgcMVE07l1Z+/Qr
VBed+2NvzEAj3bYvpfvYKtpmgjem8MAuAJvbNU/ikPCRTuhvWbzkdBS1ZXBB3tvn
Pg6xiLODTX48UclselLPB7UqP3rbwgUxBho8e8Lz0i+iSyN1SPLnIyuTDEtf8OWY
hnZ0qfWlScT1W6zPg4vfx5jM1IcBuzrbKLyWOTMJw186zuecSMncp10/yFAtqAik
med58An8TMnOgYgyse+I3DLaEXMQAZ5ip9CqbcM9904V0bxIMG8a/B4oUA9EG+mn
+CYhyZBa4NCPPQtVvlLJDDDB9FiN86WfQ2LTGy33ysry+aLrI85FH4AV+ey1Hp4D
J0ufaadcUPhdQV3HQau7EINliKPXLqZZXvAuILUbXdBC3CR5hDx1CM0o7tau3syf
ZVkyMRgrAlv108WUPfdb8+q66vNEgT/Q8MSzuFjtswEYEwgdzUDpmM6CLYJOi7WS
4daK+8LryNdTpfOk4vpvYoTnrLQVecA3uTcPLk5HV1y7EgPJNe3ADCCbwan1ptMT
Uhvdjqpi+ayp28dfy+VM57NQdR645Iaa6D849lcjaI2a2eP8Jh5K5KsJmT0KbEP8
9WhT2ZhNhtK/o3WvNaIH8gL6HvHBC5A+zjzJTiqNAXwtocwPbSm2QRjHCg3U4Ko1
+fxE+yLI4WV7cfpzAD+Tf429qzXY7HXw6a3QOU7W9ncHfq8LFJ86XoHK4hJA3IxQ
oQBVgzUGI/mJOo920T48Im3sxoCKX6BXi8meGENbICueDW/inY8VEHMiov9e5GBH
MehtzbGg0I+38pfumEeshG+pQda+/BRUfXGgLfn5Y+VMe9Fy2stlloL88W757wJr
PXAXPr+UOR/H/woHzDxDF1In9WqIqIInxnY/rYyQXv3DvSOLN85XpO9gA/l0dhKY
DLs5ZleuFAtWQ+B1XoBPZFIH4092hahyLhKOYSmxJwA/OJJdeyGsZNY8vrZKAv/b
oK64x30nAMfGUGTP0mAQ8Ff1lHCMflguKLsJq9NvJH4/pOXmje/QvkKrTxlxWTPz
XsNKG6CoV3KCsvov2C5uyzaRcBJ2fAXt6OJJ7n7gtbcOHnK+89AuWkuNg5GwEh3M
AUBV8NAkrwp7rc2wGzkfv/8OgkxnzMkDfrRRgtPxNMskCqJ9OV/Nb0ZBih6Jaa5t
sPu5o9VqUfvVIWntuyrXX3zaJT4VyiOgfSuSJIz0rcm9FwXiCMC5STWixLy2co0v
1fXzeuPSAZsi43tbWtJ7z0hcFULRVNLEQmgL4vNoDAAzkF6fGddrXx8wCr47UsEy
+0MaMpiLtb/7LK2mHmJuQYSwFKU4GqUSzbdR5gS3xTEmiUjkfSrMPSHVT6BaRlKG
MKa9RsitmgL4ujXppp8SiTeuXpkQfaLOvfWi+j8Os6l0AaMMebE5ewYgKxaNHTcN
4JeeqC3T+2tR5/0LPmOwqKF37gzYV39ser6AQtA2EOo73bArN+dxk6j1wT2MgbZj
/0MZU9xqtBx4dCX+ASbm6okFxxWTN0GdqC4vxhKRDTrDPBZIweSnFiWrsXeF89As
E9m7RakOP8xzRlOlnsZE6Rj2ByIl2Epg1dgJulQS/EfC+6I6EAEkyQILG7D2KhTv
GJOrnmMGls2P9hNCTdEXL4edbgf6GD71TNVRhljuwtWbfLyP18FK4zPua20G45EQ
UHdGZ1VpcYluuCNPz2V5DBiWIkia3RWk967pOzprszxk4f3P90EhlQUfc8xWEplF
AK0sZtrHgdF8IpkSaQaeNBH3VC1LfKKeroprnjovwplsZ1xC9Zhklln4/ArqcBsH
O3gnZRq2dTcrmhDkQgYFq0QkBuq/UW66Gx4IRvuZ0gLIZSXAeLK/3vK4nzKHlVxB
fJRKD6am2iNii0BeLyC9p/RzdLGfc2QEZHw9k0yL+s0rMmadyQn5koDgSnCf7Sm9
rH9sWU6YEz4BkBsZNxrOBYfDOgcfwjS7JDxtBwwAxFB+by3drSQZ3pjjosNrAMkM
jqM5qbjPJzz0dHKUrqOtzUZ6kCpjapE+tR3C1Bzfo/MBbSXR1IOwOqjH+wb91zdq
e4l0R/1KwPcNcmiMA+4G1MHZjd3ftDWhwS9bRE6iWR7E8yB5+FBWJ21/CanS2v3E
F74zll1nXlqvk49Nzjdh4Rw346b9XBVrfRyA4Ul0EyYCfv01NxL5gD1Nk4c6GSvD
ftRkIoeqFclntDziyrCRxsbcI7L6CYXcF/GZ9a8v0E4Sjow+LKgYPQi9SPFVgIv8
FQbnXg+6r462Q7gx5ckTGJeTbrZtdzHqsI9BCXxzoqsGN2v4OGeBhabEXvgpFkkQ
JR7qdvvY5YSrMonWQ0WY7xFC1W4rm2ZS8HpBzhVcvKkbEEqYMzLUZvJJBGqXuORn
z6n94LSGk8uJOT/FEAt2XXREe5SSJ0VHBgwaE8A8i5BdeSZm01tsZTeMQvwNGPNM
OgREfqesMx/SqfW3BOWn3cyqXyOaCqBCMrpmspULBZuTshqU6AkS8ck3O/lt69ah
uAdSBophe74FohMQZH9NTHDxANAITCS6NgQSXWD1nNbl4lc5RFuRX3/udNh6l+sU
mDUQbiT3TVWZALRypFTMppk8yO9h2yjR2K84IdfzgeIVdC8RLYlwkqUmf2Y5WMFW
C8j8FG0uivUw/RCG235DHdY6Wb44uTuqfLLadwcnwfybwvEgWjKXhbaSix6Bv5TR
Yy0gVwtE4iPehqDfPkxb7LVl9PKwbSaDIFeuIdRQBvNWSR79Q1PyM/j7fA1JJXj2
3t/V0gjngmU6QGfUmGkKcKhYVyGEyAHtto/yAXUuJEQyEzDNqRo/5zThzufHlWbm
lonl0+2xQwUYqbrONB3FqsxbeIBb8YhxxyzU65BYGY82kB17JJB88iWA/uxuC81V
ExUgd+u6qGQUr1A8mMs3gUd6bbFerBp/hZCypPIAlzN8ekLrXiMgSILsOe4BRiWx
B3b4/PcJDHKCc+Vh4+xkxDBaoamaDEMLp2S0koJ4k6rGuBHt7BR0TbYoSTXcNh7o
Sw/rw3piWbY1x1F4XAjJA6pqp4jP2Y5uekfDqUwfaCFi62PEI3ZU7Ew2NxatzmdP
DtziSRSu2lu8+CIWODwgX9LWjMq379r9JAdf9kqF8iFYFqqV3OH1C2G9wH3mG1yL
N8oIBll9tzTH+29hg1gZrODiCjUaHP8GcLTToh9CBjxKkwzzweLgp05QgrEnSFO+
lYWMZUKKaw4lK5g6znEbPU355mW4XcCUWfOqC+juu1C8oFOwVdC6BJOY2TRbzKgL
NmQNBYDUk2A64w4SqaAAcK5sUc4yEDakQHU8hh9RV5PBztkZKqlZ3d4CsAGWwEMY
/DIPoFo2Ayc6mq6rZs0jjzFDiBoHg+V0uC2WsAWwmcAycqSuFcoHOM6ILGAiWkCy
Yzft5zdJz4BPwmkfkTY4TeGl06ZjVlc0GntC9DQP85zw1fQUiHKHqR0Ucas7PeNn
DQkD8RC607SznMPtXycs8BcBY0bLJ/jcblOB73AJALK30QmEtTAwHp5wPBfquaDQ
Bqct2XFR+x1JdpSCOdRS0TcZOQzydTu67f/zdycd32l6Rcbw2WGXUjuMOtPgNwa4
27AMUv2p7y+SeJ6RI7qb/FUi2ffhxuDuTdGsJJfELeg3U78+kFIpl+Ym3lOU0aK1
sFAHr+vjtT36ichv6yjeyrPp8Wy5nvRfALri7oeok5UE5VRopL8vh4Y64Lbv+XIJ
WJKBr7cFMSWor/QD5CQ6C4VIbOl6d07CIVo57Hc84nprMd+Z+hNfhBe0d7pJvtff
DIJ9UGVWgJT5wD98Xo+ayRfi+4ATVMLlkEWTmMyxsnD1VMThg7rp0FxJqLWBnyL6
NMFwj4rR1AOrMoDsFZ5oRChtktk+QlgBnqHd7NIPgYy/dQJfPGBAtLomANsylEGH
Kvbrz5PkAvfKWTtNY6iUz8DpZ4ctofxHk4mqKS+aEdoF3Skzb5RTEHtM8G0vlkzq
+sRDEnhe2W4iuBt/Q97V1UQ9OolZ0xaaUM+UiJhdJ3/udM3JPBY5Z0HRslrQKxN+
xz+vfuz26j9ax0tvL8rkVtCNEsmO1ZAeo+vn3AqAfZl4/A6eHS8f/2VvaifDYJkx
/1sIclrhAHXESdDNxknqUUwznmVOWaieLbluymFt+HZcZajlxUqp2MiDl+IDHZqy
KgLwRuzLAxUpDAHqfDm75I2+/C4763azxrwmAWw1Fu93kzHNTwRfHxwf7XLqN5+Y
3lnNyLoMAB2Q1M86blbpUTcJ4N4HNIOQvyJYhsDFyIabe+VgaY2Pdat3XH7dGi/0
bsv03Ov2IOZHV142X0SndE8D6wmvY1RnY9kid/M/ylzo8dV620HR2+13nYcsIsig
EXJ/6f+6iqaQ6kuWgFeZTfsycXOPP1bQi12zNa9x24qJI4xZjYIutDEpob8Ok877
uxnVPANVImcTw19vi1ZPksgYNC/2ttx9Bkk2cON8KTCazKetPy8rNPr55XV+1q1a
t5NzZnCLlNvyWQiQ7XGtqYtbkcvxNQKMtXXnDi73FdaCslfYdZV7VPaVQVP02GwW
tBMeF6P6pbxGyO6vzOVEN9EWQSWqj61iPJiIXj1tGta481s9XjbF1RnmH+XGTBkz
y0PaiAoWGloeKBOMv2L/V8dIfQFu0eOCg+lhkiRL38LD5z49U7TQZHg4OaOO68bp
0C+es5h8oDu5mgpgxfVV164vvtJqcWDrmAOnOBHkYVupDWbzOx2D91i2VEqU65UZ
V/ntK6dXmS9zZP0eKVWTs70Ku3TQHvNnaLyKOC1aLFtqogzqSx/VVnIPqt5q8wfy
wwYnJ3T/QVqSWW1qW8mM0SH2b5eUMOuukWKpSph4H/UCAQ2W4FLpyNgahJNLSoIQ
02bFd6oCeC5DG7Or+6NO8gwj4l8ojJKRxfqsuGuZjkDWBuOXtpuXHa+0RucfHWle
JpJFV5LnzhLVm+wV7NKmrHq6sRx7SoxkwKmh9ejGqmhNqGcMujtlpsR8O7vBCSbe
dAsCqeQeAlgnfQSUwMTDIgTTte1mgn5lmXiZKBt6RNz06DNhTMPYBsrEK6OMOPyr
f1gQQWGM+YKZJnjUmtdi5NYuMPodZK7Qk9PavT7+FCxMFQXhmxje5ae/LZ7rRRlS
lENY3/PUtHisPNDljGdESRAVf6lFwf/s+wyKIv0/ZjVoJ2gZb1baji82wo42eHik
dql1nlJc3boPJU0e46ThKyz0HXERimpl96oIlU7pvWEgaYL1YP6YRKN/oTSvDAKF
X0onbWXHdivKeWz95B4cw3FwKV1lN6NfTGtkizMXZs1+UUatOK8FDrVzKtbhRm5u
odOcVNx3NacTzk0jckDAi3PMyIY//M0kwZVMP/BPDTWJJfHoOxGKnAG3b7C7WPMP
uDtPohnL625m+0wzOWnqejz8PaXpwukhUq1OUCd6mGySCTmXxudyxiTRi78WWRu0
5wK8lgo5deHuxWfCwLWqiRkAjx/MnMH+TogynzKyuHRRysCGvaMbRAyhnjAqXAhF
puqmjE6FLIqzqLMdbsvqFriBCO6e8SzAcSn5NTQVFi6TmGB4BjERh1zZiPa8TeRz
qIFFsyW/IOZrvSshzMo97p2lm/CGUXwENzKlB7RskGlbFEXuUNb1TG3U99yEACCv
WkDPbZzqSMoCvNaHGIET6sXngvvSNhS7tYmkAuJZzLR/H+KMGzHJHJ2KlEaXUgHs
UDeIoxzvMH2ivi5C5/JLC4FSJfm9pxOvHJYIrpSqiCYfduE1LiaIHOJAEdZppAV5
3TCv27TvFLYTUF+oHRK76AIBBD0gIM0C8MVczWbYjPcAz7cVrlsGizCK2pSGo0w9
csYvIkTOLuQMBMBEby5H5xn9rWiJJ0Q2NmtXyDVNchn2e/J2MK+wreyEVggLq6A6
AArr3wO11Lr4dRnHDGfQpTLU2MOCpbgTflUd8q49SM+ur29HnqE81sc2QCxT9iLJ
Pi2jFEQPC2TjlcLCiap7gwVl5ZfOdrYLPjBLNbbMW6/8cUFAddBhixM7dEUj/9Ct
ddYt/vZwfa8TsWREEE5Omazplojw89c2TA8N9JcXQENJ5xxELvdcSkK0rFuWI+dy
PKiGCcRccuXrWoEXsrzp69StTBRUpK583XuR+oi/O3qXo14J44UxiwZA4PGIyqF7
d7PuwXN2aeIAu+bhTfivDhAsaXAGjSQrQPA85xGHZpkfCJ0lz9/jd0WSzvlaMxpa
n/zbuwhLOBTGCccsePDyQeQ4ApIPY4RpCDWm5B/6q76uqApJLlZUS9lFFC7xJjsv
Uzn3Ww9joHWO36lfgI6sq5l037V6jIWuJPB2YedtvjlId1na4QyIJgf3BYz+6DQh
5w+LFBYYguj6jU3CCJiWWAjza3uloEgXzvZwm28YZyUbYMFPL0D/7n/TuaHadjM4
fkSr9zisOaMHnXDLSnH01eS+u//WSgO7QjhfE+4QQBgYVaUHMHM0KC4VqYuCcnPm
qmVfR9ItrC55TbBoBGwQY7thtG7BU3uaachXBuedgQ9pq0lzdrQr1cJYZat6X0N6
z4Snmjjityahmg2YJvtfk/cw12Pys3ch6r3jpzZwly3J/BU6ECDvtt8tL1rWGgkz
vzbOk5J1I5/radnejT7jpjBfYvgZKCZdXm0iDnB8+shfbi/hLbJd8Y4kYGdtK9ID
yO28H1LIBSvGiTns0KjWAJKVqnIC3hUYT1bho/z3wRQHVQGTB2IKqP1S/vGZFOFd
yQ2mIUheL4ptM5CFYZVMBYs32SNS8smu91v6UuUambmjunpIvivQppN/SSe2ofxX
KnGwgds+6Lfe6JuziCv+zsvEK4eP/+FO5bjgx+GdXY+LEIzdp5TRvOB/aSHYRiWU
YvmCOjgVssLUFywi6fP/Ha0xO2kZRWi16Ed8K+YkDS+Q5sZ0zNqu+f8eVHiwbFpb
RGdM9INk9nnYHvWeQLOjjF2S2NsrOZoOqfaw4tz5Jjk51j8JTavcQKM3N4CiyMdU
2WgxK/DSDUV1ozPDVrEYlStzkiHE9WbhWOu05xoBi7JcOoDq4h7tJE8HA2ivxYTN
WbS+krfhJcL1kHTOmhxGC30a/ye58opLxlZ1Sv7XmHb2EQEVVdQx9m9Vjaawy88s
ZBQLCTTBr0HU4XUYe7wCJ72bazpPdBObbvxmlRb0hyH/SbY7hMfLeYwlJKvw8GR6
mLtwO3UOuEX7CFelaA8ZrqYtOYx6AJ5CesZ8MaV316EQi6IXWCY7kHFcoiQFtOAt
/AM5fUIBWkpCW49ZcmhWpACrLrf4QwI/4981QpMzI9ALbhTYTTeG9teB/QoTENGN
w1mJ6HOLkHAodAHnHUBX6Xi3n6edxkmfMB8QvrD05xFltZrLztlFe/T9GRt3LaLU
6vytJTw8VprOiLhut3yy5lfaAeAA7Mndtz7FmFNctlwcolobzJRHuWyp2R+dVxB7
Z0EvMBu94+A5xDssyhha380Dlo62lPhr1dQtfGWIHcMgfwsYjsqeLFupSzTcu1gx
TCneBmWCv2F4vijTVGD2LH71Sz/7S20bRAAFqBDWR8IsjyviKWYti9DOZTlkPixB
eEvX4QdfsGvpvNRJDXaanRkKiaQ1FJzrw/klkAuudqPAt/HKk9CnYwNR3+bPVrCC
vAfDsVi/03JoyvGzqJpKqZuGjD7vuXYbN9lAeSQkwgdxIwXWDwTFp1vWqmWGi7Uk
mASMz2ma58tzIN1OtTokFxscoVWdBM76bM4HiOzeb7xZtRVCGwElKJsBsos4jSq9
XxV0uwBXCX2izo7nNv8MvZkJYYmPeysG8vtiu4CXnkFNyJwZxVas7Sg1nfbBpUqY
eqDy277BMM8I3kGn6zKGYNUEI2Gu0X48dO+K8zM+ohFbWdO3sH+Tnjv6h3ScUj0P
wtn8g5iPxE8bzHvmuG6x/KyeXirLlVzPHNGWvP9vjH475DN2gjC5wzOkJaUJAud3
tlrrE0gVmovIY7tgqrbzUjQaIHQBS/oyh9oHYXeBPSoSW4lkjIb/nLrZS3POj+lP
EwgQ1hPfBVSNIGL3QpkcEDaLHbGlATJuw5Zslq2lSMUZF/MflPqqCPh2ovVKjRqT
Z2pp5l1E97ReFdPv6ShkOAkoCEeN3ilBEtynZWuy33D7uZnfLunvMInWgMpl0IiS
jQ5q7FgTYnm5jsMQL8Vr9JaOlHvRhP9cB/5UX4lQm3alWwlJTvIKQ9EpF2r4BKjQ
ficyoK+ItVchcy3yam44J396SfnWrgDkL05zbaJ1KuYQS1XV88hN+UHWP21VIKpj
HKkX4fyuY9o8X0VOqs1uxjJFDBS58owT5tDOYBbaDCjJjZjQ9dIQHImcTEpvb9jh
BTeRNZ0Wc/ilbUH8ZbZfmiEeZI81CsLzSkVv/t3sKWPSEJsdm5RmidDw3nR4/bNW
/JMPDpsJBoyv9mYf1ANX8AWH/kRB+Bl8uQ80DbsXTvPR/R8QA46/n3XY1N6vD/fc
xSz88RU27alC3dCX37+JFERMYK45amzwxj/i+K8D8Rnixoh3RZYv/rtdAxlu+hvn
A3MK9jyeeD5wqsECEWwo+eMQtpGRLq8J2CUnmV512oxx1nDZJmrnqzgKfodec3Cy
HbYxRnJKMo/pysPBZqdK2zXDpTllPOocmj9bjjVYqU14q1wV7oAP1bwjn1qtwKNX
/gNSI0srEX6TlWBjmOYnpMdmoxvXp7JasBvjG8xO0aLKHj3nhM5mIwc/GbV/YIVp
eER3oCO6hTchWuYocP6CvcGX5uoF6vvYyvyyDfE8UBizTgtZdoiglb7peeZ+/1zy
tAzJpkiod9iXBRtfB5eKiIX2RLIuJ/kg3mGaBMqvdU9L9jY6njWprciIEYwkKPKM
gFc5v3aSht8wxQiaOiuup4efZkb3Jha95wjjecWxb0kKmURJRSanaDUgvbGEcslo
Ga1ZI4NwQEYGd7NjLnj7TWmeItetWVx+74tXFyvI3nk6sa1uSsGVqr2+VlaByfXa
QrSWF6QtJslm52394FiDjy2PzVJzTmNQlPb3ytzw916GsKb/yvI5UcqWEHVMurN1
uBNyhJq9xK9/zzV9fdF6bg0YCLV0BWVyWWxCSmr8pOaLHnVSdQW6ZFC0sZqU59qq
MHT1axaeQDi/oSkgl7R3oFlAYjB9Nsyr1zFiVMol97qT/p+8HA9uMNrRTpDHkPnh
5k/FHSQFXrF3LM5TxZc26eOECp2HDvBw/Sq5uLYjJnQ=
`pragma protect end_protected
