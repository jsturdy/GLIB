// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LvdJogw0ZORtyF4BfUqWdSEA6TVYC/lcIr5BUhoQ9DKPOG3xhxr/grXuuOVqzPIS
ZeE0uJk8RYYTRW2BeKxZzsQYiFn+yO9GyP/Txg6qy6w8vPt1+y0MpfLxcK7a9LmK
VD1H/a78U16qF5kInx0YJxKhiQigMxvdU6eM64UgSzw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 59184)
TpwJvbz2CceBqJ34O8yzp4S0Ajh3zH2uCklYQxlXFOT4D8otVtKqniwpxyleYHBq
IwmeA2mZE3CfRerhFr6yQw0zsFXNgXUUI8AgsU8VnwAAR9+KJsdAR3ZFvHWrW0Dr
pZ3XVtJbp985pgMEt7IJjTIU3K8WTisWS2Ih/tAmPoouPN3MCbHXffCTjLEvVY8F
cuFGHclkwlMEJclEg+hGPbm+b9TUc6ciIHNZMF7bwQV0zJYAcpWpr6PIUoaEJt4U
kqUK7xKO7MIr7/5scvad3kuXvOxjwGgKqw6V1wcDmeNHV5+7FKO+d5XEKSOsiyUb
dfgs3eCJdAVwcK6YjctfCiEzUfeN7agf8A86ka5AYUUJwc0IWdQVlciUwALwQQTG
kTo4Z7gHzl2yVTGec8nQ/DZFPUs0CqhuV8jkkxatqnJnXIYTQ0AUePJBoqDJRjeV
lYTtGHyuUGXazPXx2ollLqVV8PYktE8tL59lCJRpBTZj+j5cAvYKK9U5zUOU/itg
24VAhNFmullePzPz3e48A2RCOk/ztPR4TFc1+PS5otGtLvg/yTzL/D2iUg4zPPUS
JP5VYpMjiRgn8PCHMWG8daH/ClnaB1RZP5CkT3RAK86ulKP/JvgCpT2Mxe+qcZ2v
WRaVcpNLcbwoM6w73hELStRwo5vlj1wnK9g/BC6QpZKTErcq5u0pyfbqP7u3djnf
nCWwb4ohZkoaCShqpNkS710SiFEDxTmUJw08FnW970TJvkG43cEgXE+vyRnF2BpF
xTC7nd1jaDL2YcBglvQnLo/zuULHTEdjQ5Y7cR4Bhq7jA/vlEE1zJ0G6Qln3iNqq
A5z2sOjhVPZwbkSluPZ9ge49OxwJnAyq+oISRW7dkeOzkK9bYyjy6THOt53mYmj+
yjc5nHVQFPcG8ROLoAxoHgAQYpZdV6Kg2cTj3GJRVuWzDFHtuhICE5wPCDr5PAyD
r/7Vg2xUY+7l582LRe02B3RXXlDvxiydNjYKdfvf2g2On8FNj8brTMpsVEsjihp2
mg9zcFkVFpPo7NYBCZqoP9IqD0wwjuQs+Xx54vK6uptx+dbwHqLDG2L9c1untXdv
JwucW0rbFi+i62D7uafjnqzdhTW+nA2iOUkyQS1hNbkQkztxPttbTAC4QsP4NRa7
ky1N1m/cy47wtHi2GXqoCkC3MVL123oIDlzjKwKO3L7DJ8w9yQ+tyJbo0tld1Iy1
/z+sgmlL087Kbme75o6CzyvkwZbZmqrQJvOkwIgvLMcl37OEpVkFUHLR1JuuzvNZ
rDNQp8hIgFyFAqJMDitmzgTFmcwMoz3irNcLXNmW1TJy8tdg0cnwX8aDdBZSnvOo
Q59u+diQo7wXy3UAgSb3uk3ba+nLUx9+7F+IpRc/f7BvQZ3MdCCjVE1GDKO7TQ57
Cjq/EJ5PbbXU6N/VjoRBrgS3mf3z+Du47w6jBszrUeMXX+UO+VOhoyxCSgzoQ2n/
o4FOdihKEJoLq/uk95lbZTf2rPqbh9PEYa5hzsS8Ikoq8Cvf0I/hrAKZQhbMDcfF
IcucchFU5xPg0Qs6n+mTnB+7/ed4ueW+lzUJ/ukAgugxi3fkDzJtd2Trejud3w72
EK4gQTBEA0/wv/uEt3Xr2ZvEpwoK1rrtqwh5yNJOisIZCDwbos3OX7iReR2angBK
KRR/9mD6gxX4jqhjmzyEq/lMbt55CmEOO0aH55yj8IZ2OgD81pR5jgw2tfXW3Fzn
C6lWvrZSdv8UXjkIl1SY6diQYltKAUrfVmy2KkHsdQVEtBLaaSnXDUBJ5grNQbXB
LAcoWBn88XBXDp26tCUFz6OvprBiiMp60o8yYR9ajK7eabuGI6WzchLuJYl2YK/h
ow+tEQbPsATS4X08GoB80aJxxKJRk6U7kN3FrCPd+TbeXwbXnI9m6KngfeHWa6uI
IQG3Z2blSQtN/k1x28SR2Tt8HlgSmPa9gXlBpvgiRCJR9x8GdeJtPNb8TqysAG8M
5VpcqfAMys+AsJPxvrOVfkMbV0Uv37fPtmTwz69LAtRIOQohzXpqMxEsSatySS9m
WZuFLHVJsr9gy96I/fVb0jIr74aesewY19nECTVhB3ikEN08YemYdDqi+DCoLEJV
fVJ+HyH8ZJX8O4HvkVvRmW2zPyN3AbCehuyFloc3BOeJlJiuz8kahH9g9RkT08Hg
NnfNAtcutRrln3F6ERSYZstccXvPoIXB0Ubhow0Q9MnKdEv3JaFL6k62CFBvaY/j
TY8TUzyma7V7qu1JR6Kg9WPO004L1Ta2WToxXNZXolxgUBBUC2FUHqyAPOo0YngJ
KV2saysSCc5bY9MJ7uxZgnQAL0tLXUuS7KhjOat+g7nrI4IomlaFsbyJ9WoRj9m0
ZytR0sSbC+z7c1wasMgaiQvsdGgkI+VK240tighcbnEPCVLWOby97deq20Tis7Fs
O7mCLe/hE7byURwgZu1jP6CJpX3nlcu9WiDiqPYt8c8iOQ8vz5EYqqOFnPVxrhg1
VzirWo7wiwFXs6shXIhMN3dv+68MbB+StdLtcqwFXf91A5ABzesUsjc5s7RAq7gI
mlyVue6y9223s/o7uKDL1V0e7bSOyRRWvVFqc/iKb+hM3gpQIO0jA7d0hENplEMN
xD7TkT6zxYbUtlv185rVk6VLGXIkR5AP3HroVnx08AYnC/ixRk307EiRMWuo7K7s
07fLA7l598ypImfg2zNkbLU2BrPbVKJMG3aNnMj/Hb9WjssaqLYrVpt6ZbCnFURf
L7WBiR2iOgfmEhO9XFkhRXLN2ZK6cGZwMZPw0gJZlFy3GKKmUUtyhLT3aVNQHovm
vVIniGhRv3SrMk6yG//yndd2JLdl5zcpSQFyNHriLnDwfs+mv4z1c9fsKIpbl8tH
tEDoeAkktDxVmhQ9e17GvWcKepnL7z1JuE4xvTYCmnc2fVjdohiNHmQAgKWQxH2Q
zISXI2XA6ykUSCQKspP0iATrdinnaBr8k5ZUzJd+8dU9NZcKRelUqDkPi3UdrVW8
T5w5S+9J1j3cSKxrRfDz6ovDZ/3XeTY6OinuLd7MpaPwA+jF9TUOI60CUPKX+tav
R0aMYwdmEgQgZ8ByhpjmJkXE1llElq+BJVqKZdf91fKSaq8aHCmU3+1hLdivBhQ+
39vIzcc8LRo6sosIEwPhl8wDTzA8WbzB6l2hGKSSnyCj0q8kQzNDNU0u/sMTnDuu
ViyWEkcJkH9l+Lh/fmBWiiDIBoy1JrxH+FDHwTd+GcBYzYln9lo12+V4UI0cBr8f
OxRsl05XTG8F17EtZ5tmBSecn6sLi6LnNK6+TahGxMCZotJ7KC5Qqydo0uJAs42e
L7IRzpSHT+UFALnaf83GNRwevf86ec+nREjVGKygC/Zk1sRiAzsnqO6YSSUgRng/
9A+WX5wdk/vwVUk0wzGbS0tBB2x8zrrLWDgwvxAl2+ucawGo9tjJ7y/jIb1bihyi
a1ZJFzwHhItSSK7KFrF6rdNvzQbOKbmTyHJMEAhjg6KLuv0zC8rAkaZ/VlWncSRI
rqrjeoi8YtrD4sleHrqhpEgp1igh9tUGdGgE0jyZuNy7kRZ+3NiL2z3Lre0BG2Bd
p/zrzh5KSFo0dpFzhzU4tHa4lOOKaD17df0GqbieXhs88Bm8aTyp/B4tbTuRcgea
SLcUvcipTh2jzl4hOsbBQQ0qZeFte1P/77iGNEK7g3L1+zsvnWAEDdR4t2ONSxy9
1ZF6F1dxsgItB23FfVEYcjEI7qHb4lxWOFx4kOQ8Ed9Fq16K/QmkDC8qQqWjj3jO
N5FLerphFRk7gxizZesbeBvaj/dRViAierMu4uamU/93qaixb+PWMfxv3tGjzxza
1xAPghTUGuhroDirb6eq20P/5pCR5K44V/eLlPTbvxFGwHQnXUXPWePnIjKL63nX
pt1xLer6zdt6aBjIWPLzRp4a4a0E3VVtgwdcsICtDUbj3lkh4tMIzQZgyNzAJ5uL
MtGVZ7DxnG4/yFHXPuPmrmmvKRhpM+tr69n3BSZAhmlWydFc4jdyvDKWAkzKTy8/
REbAjtmpYno/t11FM1ju7J9Yo/stwoPCeVMM1yU7QaQxVV2pcxeNmjk3P32XgpSP
Nq9OZveHB42hb0DOwh6pjOvx750RzjMyuzgJXRud/4RqirLl/Ud7rfwjMURPXDY4
GeJokXn/rPRMl3e7/gdSKD1MfFJJZFcMOniXEfHJFVW/EufIZpBoStB3iRN4XuXT
XyBrG5sAR//k7cEda87zRRUrxWyr6tOSSyAkcYfxd9xBPN41n7zGRlwvtrToVwI0
XjjwCDIqI/pjVuJNeY2jA0q/49q/jK4h0amm0uD260HYWvjNCrFnu0ePVf8C5Xsb
Zq17f3MCKqcdS/kQrdLDKdJRUKLp+66PfvIzCgfbdmagFteWcJO0fuLv3G5Y2rQx
9s+Ma9QxJQwHSbbObtvcWLpmojzCVkY32n6H8X6gFCZSUygQdwyVD8cO7LQIc5Cd
EAX56HWRPZ40Epriey9LuneeXUyXEzWrnDW2eCvlGraBvsTnpGTjGT1pnNwKmM9J
dGO3kJ84DOrmrIqkC0WRN3/cAExr6+cnQdJQdX8+2/iBdWyHhyLu4Hpvxe68tDA8
AVXKV69DYL4KcGK/JkgwJOF67aJZvV786D3Y6ushydqUDBFA7DuXkiaXTzVqjnel
SZK7nAXl9EBKxFSHaibUNAT7Gl75FesNYcqgRmGMxEiWYhtEIO4RxQLhngLVBFv/
Kc2uK6I2pDLg9YXnv1kFDDX0o5qSRWO5fIo2qWnSn9oBySbBb5SxbRtaZnRLKMaz
/hvzd7q2DIF2oHbczzWpLFQ9ml1YpfNw5Oghyn3D2Loj3e7SKz2lT0s3h/aeCQ+j
fW4Fbj9sfP/CJobXkjIHecRVjR9M4oWThlFIsZZc4uvIyaJINVXlIPaTdLUDKvIR
8ghdKgPZpDpwJ38WytPAKcMOcM4d22ObW3LvU+grrNaetAX3RQzYV+gLrLVtFJ0I
o3Cq6qCppNFRpslyTPsnXUBkPAxoWZRTOlcPscwolzTFw+rdQE+WXIMvHRHzglF9
/q/za9XCHt6HAJNex7BF5pfdH9BFMzcaEwGWjA6KbpJodXfBlAGmpsRotO8QFSRn
bR11cKakVhoAOTQPB7ircVw1q31nPWOtCPxoa8Ugxfoq2V0FofCXXJf9xseWFv4c
KSQY5Vtuvss/VZHuYej9JI/Ge3js/kJIyC1UPKXl9vBjN6i90F3mieqWhNtzAdRE
aKCeTq20P/C/GbW8tSA8W4RY9UqLtsA/wgL16PyWaAwAyvaRKhjPc/oi6jhgPHUp
vfSGOrzNB+PT5AprFVUAagU7H22gYN2SaJTaKRiCOxqyyBlZPyc2N93CknBKa2QJ
yOag8XQ8zuWmpN/FH6AWSoTe7suGCthFX0feAJ33SbRSJ5lLJcNWH5g/J+U1mgt+
w1KBihXbo/cm1ahdtUciZ4X0aHWzGJPzGpOKHCX+qRAzANaPC9j8C8zeailPjhGq
5eQCfjdS4VapTeqd6bU6cjcm1EKBmbt+x35NLYUzkbHSdEZKe1rgTHsDJT6qmo3o
XzE0T8VqPSgBsvCRvVsM1HWdEPpJx/6+mM+trw/QvP0rZQqmzoM6Cpp/zg1iLOZO
KbxhrmFasH64+a/guJodofqgQEjb2Fv9sVw8X14y1na3Ziz/4fZ9PrRqHdihq8BX
wmLMr0b1Q4XxDJF6djnrfaG2bFUlMn52S4s4LEA3DM38XnHSe8Wda04PQxzYNfam
ZR3k5AajpBuLT8VzTQrj/miQfFBbefjs4ozdBxeoxDGsWdf4o6YRdvZaJeZBjG3L
Oq9WzV2MG1BBw0LhVLAc+CSjXXR4YvgOaFvi8uu6j5ixdujd0qCrI9Og8gPXxAwT
DHYXkrieorbUL2RrQCU8lTRMSZ5WtDEpB05TLAUZyDPLSCpMkxGiTHcvDzXN2IIL
gg7vRQQzRuFJg5aPSiXDkjWNQ5J3M5F6FQorhnLuTZQyP0SewfMgwzcwet1iJ4O+
p0SyQIyKPcEsfCTH7STTBcnMf/NhYgQq4TnIyC5yPGyw6Uh/TRneBkDlpzsM21cg
N0wvXZZak16RM+dkkhl7smjUgYpBNNFRPjKCn87M2RMTkVIdYVIQKlgAwaoj+PfQ
7HATdBBLUZos0TWibqz52FuRfUveFv5snFrrdXuwAryIL52iPuhJ5Z3an/ZLIdrv
mM/s5NSJuSmnyvmb9WmLzpO9cR3Ab6ya3qLhQShnCS8kCTN3RFczJLAj+CnHhZ6U
VBONOe9jmj5M6IVTqZq9xG5q083J8kKS8o5tWbYF7rUBS7LQvHB4/0XL3Eszth4A
RwviPVjS8J6DjJP8VZ+69R5wwmrWjdSD7god98OrbB+5g03hGkuA8tdVTXwHAYyH
OutmgZ/LQavi3fDGduaTrT3r5WzD+9jBEgTdQfJs4IzUD2lMQMXriLzMKUac/tI7
7a0Raw27oxVnj63mln1rOWwY4uOqd2/iMaAaZ6ujIxMFvWFddNDqxDkURUNdB9Et
uLjMy+Q65pMTt6yG3Xw30eiJKMyFxQJGPBDJVJPqkVvlsggxO6UiEwYlXcb/I8wi
4HmsMCvzZgFXC/57UFiLXhPJlLBNxKnERIgJotzZ91DunxqHhk5kKaKLMlphgO7G
5lFNPB0q5/CqI8fTkUBP0Bi0oTXmKTu4TCtGMwbldTjb1iYO6v2ZujduMvDt8+Sr
F1qPz/3KoSceb/6ivT8xYR3sKHlbrmgxRBYtmg8y5du/jBKVUdtGyUphNG+uKerj
f2cejXoehnlCJUG+Bdq5C+xjuu57xGPxBpRl/KML8+gHyR7EWLdsR6dEZ7VkWhPs
q5/2zMgycBwSUXFPhJ+42+QjdMk6O6UQBqLe7VRlQZuxYti7qmRno1Pvs4YdfKrn
NL2Cn5qRWjwKiKir7GY7OJR+JRMsZfKNjH0xTygZH77rxk7ankgjEyWwQrmnMEwp
9jthTLRNAKZIMuXd4Jw4ab9nRJPUMsJBpKeRIFIcZmVexPkLlmnttD2qhivjj4tX
/9w5F3GsfHXWD+qko2j9YA+sgU9OhjtR4YTanKK1QJoF7AiZXcVkZ2ounXmtrXip
B25P51g2nee5q00PqQTFs77FPomqB6Aq+hvl05Rfp5tohbmRqwvno8MzSC0GZuYW
mdnr++EfN1MLicxNUorzliYXd7liErk22kEEWF+UIRdek6m7joAg4saGJ2k/iREQ
XcLGdwwQ76LnablTQ0NnANG9gEX8TymSkdBpv0b+p1k7s+j8u4bvb0hsUs9+6JXL
pnZ8+Ne9UlHDwiwqCuR4yCOLGRaPy+d6CsaXkNbslTgz2jzGVfoyUyI+P2sm7Le4
9USID6BSm+gHanf00CCIXhCLsYIssvL5Q+D1GKQyUHebx7+OpDFZPKYa6i5jezDY
NIB0NKN/7n30UbAd8eShwdeUeLRlMbIMIRKSpwsIeuFTkD5paesOu7mgCJ95Xspy
YobUFWY2pEYl5Fd3H0oUR3GXtA/NyVvs8tVoe9NocJSYTV09tT54Is+TKbEnHSC6
ep0GHfVDqmFBze9fKqo7xolEH37T4Re1HhqgKec9g5Yjr84tMjgI1/bTDwtDc2Fm
GvQDoL0e2xy0M+b2/yRJu0EA+mJ8sTpIQA1TfFtbujZD/XXRVo+87rfkW1ZaRjDL
uTvBolAYq1PFKm8dSRBoeRkqOPxEUw0FjJfsN3yAR9rZAQMJdPz7vnMhydleBmFS
67Y9y8B35gB6WR6+Bbtxu3dDXaDqXUcZfe0Kj7gvOONgCpeL/V9rZ8hMuwQQc8Qm
5wXqTH4kp5RO3K9li85xNOdXLVJl2m2TwMoP1umxLKqEwhkU2E19Us25w7HQziak
FcfysaJfan5XP7mqFtgfC33oecY45JdjrzZA60j9wIclxgXieS6nC5UZLmOp452+
V3hX+27h/vym+w0uWC6ZtYE3YU0io0K3ibddHtcA9iIjqWab1QlgJvPlOS3qEYzk
L8wKvPQx/UV9doCo4KF6RxW5h3dCNJ7asBYQbr3YkFmcW/cYMAsCC+9ICcHTHCSz
FaDeGiyKeNj7EA6eqzB4PqVwbPRG0fq5qBZDqVl6v2zWb4VSp8oXt596Xz/Xjeef
tSQSnG8QOdinAKvSC+yC3+kQjsUSzZp5vtKZUtI1uQz/kdtXEV/wDGi1+DPwAHWC
ECxhAqG1StVr4nDV+4gCpldoG2ixu0Im4XSh2eTRxqDpQfmlm/oYGpJiFga+dHe4
EnrrPe8C6yN5U06w/4F38pF9lizghU86cWR0FUib8oLx0iw1LP43s66AuvhR9T6S
3hYLgo6H8zpqzfltQP8LTdvdFUunYY3d6jbN6GnJgkO+mrp8rGO+xGW98Qwsh5T2
8RRlLu4M0IlVui0nutflSpmNL6W0kcIW/WprGRjqObf45goPqNdG+wMl+MD6unNf
ZFsMHu1kAiquGh5BZ/RdtfMoJiaWRzu0MK+0EbwQ0ub2PWcVdygD7lI/dZd8Ud81
i/FE98iSyklYeBUR7PxaTi25owAzOtNh4QS5ZsSHJ4xbZ93GGMDNmFB0hDNgc2eX
VW+mHt55r1pqUe37R2t/jkmmcFNjj0brj4N5iu364CBUsJjtRq+kDblXXGdujUPw
+Y/zyWLlgawZCAa6jx69B+4WU1i1H79VRFkGWhK5WYx2ubWv8doV5quAFws8xbMv
v2epvY8rRh6wreZoR2GnZM3XJVwD0tokJeSrABu2Q7jCjzb7FVrPB9hIXLDjgoYW
mPwteGG/ATaXlR81KGZy9Rk7sQXnRZcRZRz0LrJFo2Zth1yUJ7pHOA/UnOvMgFCy
XmOuYHfcSitMvcNkY7sUjUpZi2WqN/SmWSRZg+kiALDydX8NlK77vyigjDrdgnDj
Hmg6lEwD4i3xzDspaMtYgj5JlhNnoUyxYqWZLPzPZwHn77r2D+NYXZwOLxwWuuTb
zZAlXByvYtKYNAqvzg40NhiM3YAZpGuZzcfks3sgkXvTE3rNrhqUO2zWeel6QQBu
16FESFlG+CQMivj7HtcY/MbGZ8QXrl9nwyLvAIIQvihjBO2QWj3KpoV2TtGCLRgr
9L6xnb/F5nS7r+9aGhCiE2nEzn2bvSqed7AAYtYmDLT7FNIncaCbOKShPqWWJ/Hd
eQeYwxEIDLrViUwxx5TquB+mr81/5Re4X8W8EuBPe9JEkxrUW34P+50P0iWwmHnD
AV9kMmpti1bY3HoCD/lis1vatzQrHSCWkkW4B+jcLNaug+Z/1wOxktD5nBhWhtHs
evUZaoH/gqAis6VnA6iJbNecUfqoF1nQL1nyI1ZuBUDXisueGA2dlA4w81smM+Q/
+meyfrEGJFbvDEu6PmWFxmBSfVMDxDy5WYsqH1ehB1XlY/ri9p0MGeN5kW+XhQwO
5kwgP4XDZ4sM1D0YQW9zQjV/HKp0QOLIuhI7AYxVM9l8450UN01/mb3hhbJfQFZa
oFKxCutQktog/gOiTCvLEQspUXnzNfDTHB9ivddacrv7Fw3ZpxAXm1b4hEdw9RhD
wEHIXUodCZFhcPnCIUK4WSptGXCvbOJaIxIYKNShvqxEshnFh8IsiUWdiC9F6+pc
O+dfdlc+DybGdYgvtnxeVyNoGSSIOdy8ku8PSfe679u4l+14eKN8KQpCDbHmiXTu
wLv+SM1uB0XU9Rb0USG0IQYNjShG+Qeni1KLskYB6noMu26AA0+eWR2LXC0EKLxJ
w0f2n5kufPKhWvHYZTU29WVisJbruc2KuWdRmT33l3d6FICHIRRGseX0CalHKThG
UMrOVLMonXyr3pHFjydR7cbtn7HXN+P2IDucBTTjl6JnqWa0nhv+ztx8AOns7eCT
57bDI7dadVbuXdcghnLTW3pgHR/OBEcsQ+nQM2m1AcgidR4WAIKlMVp3yyyKB0HU
1bhZfbQVJHV2i9BStUa9lFtKzHuEmfddTmWzSsyqrRLa0dHMv3Ovj/0GnsyYOeyN
VR99mFEm5pAP8avpDkMTTd16Gl5XT6vPKeR7oARhLwrN4HxU/+B7XoXHJWbzIO/Q
j28Mt0P4GOa0ByH0q/J3gEEZf94i85B6vpA6wvtZ8qegkj8/CJbKecD8Y+vwVc1w
xVhbkAy1NmsPY/W+GLFniPkkaH6Eb363hB8YaZ8X6VRDzbvCnRYvLESbTymag2fY
6/Mnv+ohp6wUFvxY49R8SejW6jS2mWQmlpPs+vFnHaj/5Bqfm6abgxOOgl8/eTSx
RIWHnNarUGY/zPYWUdBqSc4dc+6aS6/BeTwgoEa2QSKonjm+xhPr3F8UmeLf/zAr
g0EglzcfipW+M/B6bJ9ywTuRDBYKQ6+Fr7Jrl5pQfnnU/uLZY30MmlMNI6l3gXa0
OCgYjWV0iY2ENctzstH88s+qgeZJP0ExrSgnqzysfrzPl+OJcazyLouHyclZ1X3v
wQW0gcUZyTOR36NOEwsaBmK6Jzn+wpwk6NmZJBm9Giq1nt5yoSfa/GHuGi+lDWvK
y5njv/DYTYXV+FJeBmvInGp7rIkDqmnwTfDlJBSvIh0R1bIqKBTk3rZLORFCOhh9
PerU19y746tsj4c01BHa+VV8Nduo4Rv/LiqYOWgPD+/Pz02FV1sRvJ/Mdnj6WUT7
LdzL0MYgPEa8hPuS9nsdnGuNs1nxXetzhR7Ise/CntqeGY2e6xtwPNubjejW1dKU
5UFD7/37T+lLzYexkf067bzyjMpYq6BwfAGnaKbA9BY+GOjyuFcg0qEfDenmKTmW
khk98wWFI4quRCaPRAa9ETOVMKq8+tWfvCjVhS/SQQMkhMwfOpxctWAHZPfeTk5X
5h8CmTEs2IJELRxNr6KEZ1gehIFW5uRiHOB1C4CaVVV4gjBylNKj+0OELAAEbl2Z
5zKI9SWLspqWz49v95vzkgzTQ3i6D7oHRho6vEpQBYLskjgnxxlbMPMnSDEiqEVz
wmeGPeaCyVKkkRqqpxbZIk8HKc4s1Bc6oiDsxpthp8oJ4TI/Ki10nS+ewxte1KEc
Q560+Tb1hEln7DIweV0Ee0++fGmLB6G+mfyBatdzNWkMBMDpXuBMvt6MNyGiKd5G
N7vk7wvSaGLVrY4wrxzq968W5M0EsjzTyFMdSsSBtfaEBAMI3JrNjxsuJvlHsoi/
CDDsMnXFqOV0/Mh1VQKYvbRTSQ8gLV9FTqpYqALdrPfxL6c0q/F5k2YE5J80zFWx
vBqLlbti3TpeWzREC58MqbybreS1MvAnHgBJ1weo49ChivdObiODCFeOnZAZijaD
fW7aU8xv7/+sa29vc3YUOYEVeE/qJeUzn1H8m4BFiOc0vhpEb7xLSA4vfX6dQxk5
+teisvqvwP/OQjWZs8WdybmyttxyZr+8FTKINAcq/AYIVM3qvg0kB79RGA24BF5Q
LtfguIqtD5WjC6QNsq67rn8NO77s/CzNkEJJ+H5PC/0/3swUEThzsazAXM9moT06
C+mAKuF6mCS+Wi6nTHP1HJ85NDBQmU53m38xN393zvu3LXX6U4UGzRvh6oxYyXXD
9IKsCyo01GwaLQGlJ5abIvBMJG+nG3JuOnUs+++1hd5Tfqxv14B9EMrkD8lpWHy9
suO9mqS7XJO5URQn8tHOcIL+ptG4ecWNjdqrSc+zQkYmteU5Jwr6pzvKYqsyrccI
dUouTuYrj6yJaowxJpxOA4FINffq04rCssN/vPiAmjLIrPMSYKAakQEE5bmW2wIv
dAmfWaV5EMz8QO84f0xQjPbtFXrIUHxbfW3OFNmsMicFodVn2lP8+G5ZogzhJAYq
P5uoS+dy1A86a7WAFFBXdlmaV6V+TfPR6XOF8xyyMThrorGExgK2grNtbsUXfVhK
sEx256i75whSls5rfmvzjn/fgoCwYMsaC4HejqGBLiP5R31KEONtJEcqUIdGBnPB
K8am0fYBz3nplbC9aCarpwcZQztHk0HujIgJCtPzzjLiuxkXAuBs35BVNB9vN3+o
QU4e+gMeB/JboPbWnG4o0qw2XxLb7zuXcFIQsej2cRkddWhqIjd7d9B47KXEnTqf
TWYvapqfDhrDFTKG2MuWY2muvAbRi/3hkLBbquIxl+qGXNginKmo1jyr/vYbxVd9
DJG/HTL6AKDXqlkGVKqsQnyG8VYQrupP5cV7gWKLerDlee+Z1c2HInCAfd6MN8Zg
Acl1lSHcfWvVCdtGyolUml5dsQxwhnfGyynJ7ox2RKQt+Zn3HlniGTa0AXcVIWWg
EoDM69W2AD1LPD4S0u9TuznvWvk51dkpYFZqDh32HluReJaNxrV0JUawm+ufu4dR
WE8+HovfE6e4XfqwgvfLo5WmiZrsLZcI7ZcRJcHHnN4Hy6WVAbJSYu991U96ykO6
V4UdbZb7SJabAIbqsEhjMez1gJx/vFWXUc6tezKxlSDtAQPmuI9SDDlqvz+zKSTB
3fWP6WfE8qKUKMXSv6noI9u1UAWFMtGZzv8Qd2ZOd/P2GfoKTqXu33CWhZGODqiP
YDeRiMVADCUGX0FlIgfVoCZmpwdzpLmlOXpTKAKAbqbEBe2TBKwLTVk6DeD/Z/zG
JYtaKUjdA1w1N3frr+og7Bmf+/OPUbkXQyX9eOF0DeEykb4930/CzW2cAPvKWNAk
+6wEOe4gaORFMz1BDb4lB6APEITvlfoXdIOnqs29eU75b8z0xMZxHT5l/Ow2QZfE
IT3MeetHqSx6K93AB8JRCkL84j6i2eehmf8OSTZMlPikPFZMKdkDHWochZwh1AoB
ioccPQr05e1O6q7K4G7PqTFYFTPtCcRhjxE5SGVynuq6kp9xFjVQN0N0kCk/6RG5
NeTo2Z8kxlgFj4oyN12EZrZfaSrawW8H1FRvzTAL2jx1Lt5fjOb4gVlP9DouRcUe
7H5jGfP2IUxtorP8FlvP9rgEB/m0QdsXFBcw4MlhEbmxAOeJSJ47llr9JLn0pJpR
9flzv9vEttA33Il53PWXBQKmr0+K9lFZsssLeM6tRrLxgpeEXsZrGYUGVD4D2irJ
lzD1M4gBJ0o+3Jm6EKTQCaj1h7zPoDlUKWnfVvFPsF/RhLwsn/38auEvqRi75xuu
lxTVp2O63WhVfkOBXF5aGOXxWoeJLNnuWX+e+dP3Do0SK17sV6WocgLYZh/KdAEz
DQv/KXcKX6G5VRuykgB0mGpPtp04lLmUKPxKZJD3YoICiOt6Irq5e3leatHwIVI8
8vnIN3uwsvgPuq7MT7U8IAQzhjYltPdRdS81eN9MXkXgzxGnQNiO1NS16ViOQDRT
PVXZkLv+mANyvEz7tBlYQGqvnKEkYZA9TUuZn8y2cRaVBOi23tIGdec5ZJTzkcpJ
ISSnhZEQAfnjzXW4h6ACqpiUVGevc5iZdv6fdM45zCeLPKzooyotMDVEIiFf0t+9
5oDPeeTw1118bdHJAiPtDeV8JLK+Ci+VtEqLk0DhcHiRcZ1fQ3JpZi8+dl651AK7
vqFbjeuJSq6S2rTicftZ/8wktd1EWyQ9dTESe84wmKb5fMcT/ZZvhCimsAL+5uxX
fiWlTvIv6CfYJFUbvng+YRvPIQZynqhEjPnqX9PxXSuwUWC0+BMapJLMIM7GaXs2
xdelXVOf97TZcZgN69TnTPsSfQXY55D7AUUj6ZTKEt6kbxb10gce67OLgelCUcWq
OOUKtORjJlEQQHlUk8a/vibQl4CfqmdBPNAqb3HAXb6QcV5FrEKQ7mEQv7ULUqAO
SZOoDwP1zcjNRk+rcr+NHWgcyZvPGgAMHlcPuWWFbY9iMVe+U81QMGGpyhB/LMAQ
DWC21H2gG3RfzU8CdnDlwIZ9mmjuCGpf+DR1DFUen+I7PGxaTxfq1TDOHbOZES+f
QdmJU9DcIMi1nV0v/s/tYpyKqKNNOWC1ufxLwwCtR2k8H6/QhPeNL8YIvcFkbnwW
w5bpc+YC/zvVyFVi/zB/YR4LAQgp5UHIdMdclvNSFnAlRc/pTB5YW1q0TZ8w9Egc
TF35diUg85h+spmP8Mds1ozm1gPhQYJc5cgYS1rBRGlTioVS4S6FzlQJF6lVfg8Q
Cc8GWNp8WEzSAiG3oq3uQjgpgbiOyzBX8KznyWRP+RxXwieutPf+lqY0MkSj7bFG
o9730SAwSk/SHFhfQ1pxnTyRng3FURwhLftFemKJVUFunc13RqKq3d8uFNNL5ZA0
LUZ35FJfo67H7GoMPtuGPxn2qizBw7nSp4Uq/CJnaAqdL9EpRCXf/+UkLA4Azk9H
ViNKlRjdG+fY/S47XQIWlbFELygqZiGs6kZtiRvjgZQ6GEPg3TppxAbMvB1RfD9R
uNqcBaUnuAl4zaY+b4StPa2eM2pmoEEo2fyJaVkzL556L97lrJCGiEhoTj4VDv+Y
cp/OWWQHdcoBVNqXDjaRmxkuhEH5U2EBb7dF+GHqjE5zZet08+A7WyOPAi415lO2
R/5jn9lhUNPernxzUnIv3um0GqB/4B9MPibtL7/GnxGlusCxJkDTz/uXI/oOauFI
9xAMuLibVU2Oav5EiuyY1FrTMJfqxQ7fZH1IklSwmHLut2FFtnmhvvaNDAQvbQib
x53bOscSoL+XDJHA2vqxDt7fUArn/UZWy3hLfrTBoCWOE5yQ10UeqnQmHAgTtljn
J1+JwcPXqENAyxn2S5u4VDTs6iO/6Kgs5VO2uBvCYAvGkgL+4OSsSCZpvu2O0wL8
lNhcRC39pLxloeKfXm/c5YevlBWJYUMOXyWO6d9qiISdxOAWHYE4/ga7oqr5nwsc
0I24aQ7OFaAGx6y3VEqtNN1kZs2E3LU0YGimgL77LfJq+7rl3jdJD52QdaaYcCu0
aO6WmwHhOuvmzn0UJdZr9Y0iK3XUtUdoVG9X6tvmmLaYmdMEb6UDBmkD5fKJfc3r
PX0EGL8y3vEK3jdohmn0yP6JDj5wmiq7tWOnmHeFDTic/Vh0U/Stf7tN3suNpwRo
zKeWBegFWGZBzS9HE+rk8RR34XYWbl127EK+wEmEeCsNnZEdmwMtAGUNQd4HDOVf
p4PdLcYq39BJ98Gp/CX7fb6niDbNVYsq1kXzC5hlO5QfaDivXzlT8UoNqCHojmTA
RTSBQCeeYoxc9hR4jO4D7rZIdrO4ynUjjItVNB5Qvw5qndBM/542gEwze33J2xwx
9PGXS3ZbYrfMYpXkgVnY0iSUEIxSbp8Y80vgFq8P0lux3cpiXe+qYG10e40RC9e6
m7ilJqkQdWFBqW3Wu4vo+94Hc+Gdd8iPGHu5bglPg9hc7lo33S0WFD/zAievas5s
hJsOCTydoVQEYJXIPDuAw6rfI96ioPsDIFDHWfVJj4QVcr0HN+m/MAHOkmhejJJT
o2KpOOYdXmEyy5ffLegjUgg+6RxwxCZiJM8eDo7nu1dhHONvBP6+ILAFL+wnLPsN
vdMiL5syXv83q8f8NHzir5JQ3qyl+02s8D7sCwe65ISv/3M/PnFcfvLumaismbyL
qT1+eOVRq5Detn3E8IuO7Dpm5tZpjBBRfOSGQTUeGrnwYgmkAnelCzUuiBrxlnH4
9LeyHN2o1kIpttOWlYrZmf3H2WHIfgCRyT5RUlyVO6/aV/NFE8PausICbSwasWno
n+OU1mVhue2RSmiO3v2wHbGA3FIRrCC4ehWj8jNB6f2ITsIZXDnM46NpVH0dhgU4
oPe7smXLdu/mFJD9Jv+QfnERYi2gz3Ech1UTFxjr40cB/5us3ZNFXcU7TflcfV7E
nXEXDJQ+tdpFT9sAvycypHyoLJ/CAXpD8ewn+F2vOVTkThaeVzEusbEnhXlr/GkD
PSCr5r6SUqxKJkk+B+vLd9dXKjO+tkGzTVRI3+lRrBQl1bb4yiCTSIuRuK+G7Vxp
yVABBpeqAvLaH040NYjz/MLVufcNGm1/0bEXTF6RoK69DeGgBmmr8dWGOWNRqvR5
Dnort18b099kIPYMrhgV6XciAOZjVGnMn+PN0ZeiNE9b2yudw/VfpoYso12bqfVO
b8f+tzQtbgLGbkKSXu9bTH06DzMCWoU8YqZWNdVXbah10CwnwMW+HAiWkQizPu9P
YjDqq6mbnREwW7zqCRjwLbOBgNBxzGJX7Jyi4J1jMT3PN5zqFTENrvUKV9hjOLC4
huwXS4dbxej6jKptGaoFOhC/LIOwNnUoXTVHZSseTsNrgstTslBTIvztP+7rj6MJ
BwoD206iMCrBbwxxUQXjY7LOu3JhQ9slve59bwYYur3WWRMfgMWrM3BpiGfaXbwS
KsQ6FfMK51Bfq3T9K1Dy6lUWLpHoz5yv1R9QNrGxlqi0jtfBeEh5ga+zmIEgg1sd
IzxAR0YhNX34MLzSlgWrphwSaC3dnHa3yAZjNIIsmExCWB0Ak6KmWVv4oCtm18iY
BiY3JQLttT0crtl2bNyMubJSuTIneR87jCkwF51A8k94PhuBrHVL5n9Jag7YAL2N
f3EjraIqstEZ4OFmNa9v2Z5cmxn6ceTZknPAw/vgMHYF68+jFxl1iytK7YN2Qq/p
fdCvKG72YRfiAHzEpGxGwrsiZagOe0lFNzFlw6M00ST9Gb70wK7N6P3K8h3Mhg3K
KqFSt96PdkRXt5NWdXtX5eD69JRAF5/N3/zYyJTsUkzEFqbynebTL+4qrjRmK0FX
nF3HdKbwIi7AwuGdBoiO7AsWKoFEYegLHKmMFrhXKZUzPqraYEvVOrCN6uV++Ult
rH4EZH4UtPh9N5V9bjnOMTjyIipX0xZp97PWGq5e4lNeQ7onuWiLNjtalOGtZhao
6RqRrrxYrI/KChoLzMnrgBZiFWTTr4l1w8AnCwOWOpkAysXaRQkR1lTsUXOm/c3T
UUqsSDSoK6WgF4kREPtk5LeJfCJ5lgaOkM0VOiok+J2jxrYMzM9Hc1+uJfoYcP9G
aod3a5Hoj3JWL20c9gwTkLQ6na1HypHlbEA2Uqlan9MwndyUkKkP03VRk/H+GbUc
m75sb2YnbVrZmvjnZImYsWInQAXkC9YqUj6g4btFzj5cDIN7Za1PEfxXn4FVY4O2
bGjL4JgNatuzuAGdF5y7PRvhxhaeGIEFzOLAR0HJGHkPA+KkQBwuE3HfX1QmTpxW
cMProJpX6H2L34bso7kRsVWC8KKLizdTUkfpsWF2TfXIORBEv7APl4ixGiyDnXKt
tXYUtcsnrjBWgrHCVIVzgbECWqIR0xU4DMV9HN5wugbCS5lS/H2N8TmBFz7sgKXJ
KmyaboCOgasiZaeGUhoojX/Ctrh3prCrAD3DgMAduwxIYGLNq+V75OKX8YbIxiRT
vvCXtFSs97tLDHa+q/jPwodqxeVOVdlcFzpm567uthlDXvS11jQqry51KDhVMos/
hbHb9IdQdJ84FIUdGy4/uYKrJ/HCtyvlNjkyX7yDRvSzXnnSRpJBp8aZxcjgpXYa
7ceTbhgGgbQLpD/6j/U+Dz0uo3ya5a8iLzo4pPCNfLSxKjkuZpYbLqOGf8LNROwN
xj5nhEKXmU2w1o6MFnJeLD+s/IkRK6lipGCd6zUZ9m1jtPnkedJVU3lUex0nl1Pn
zxx9BALoGJyxogOHl3LqLC5Bpcy8/YlaMwgS1MuKZe55J6TBlvquRBTvXCNE7YdM
wxP+kHHb80AEB0Wg5seAy9mL1eK+R/mlq5AKRP8BvsXPO1PaUIwyKD3UxuOxV5ju
IInZyz33zJFQzyR+1EokfVFDghdQObka9Omgy9mUABixp87apU2i1Ry2/0RMHQMF
pN/JsEzhs9lnxiT6ilqn7yLRe3ulw3uw8MyqZAzGn/4n+l3CSDqqIX/mYWK5DlOS
gW0LFKHsdsHy0v0N0dvUpH9VTIgpCVjLB8PktLVmgsX1QM5ueIpCdq9DNAF5HU6e
pvir983Lq14GdkSg912DXTTMGZqr1t3eQdy0FPxheOYWQwH7M1dO2juOwzDNC5rk
KiUW3p2Qvr87rIWbZbkvLxb/oTXubnT8Ol8Qy59mtogZnAxBL0n7XF1YT/ceeKVk
2gSFantVAlXRiyV6WStsBPT1xSBWDvC81BMMMw1784OAXbX8XLCcHc/feMC3uyGd
GLFxBblbam2b7LS/eyjfdCo5iQp/0jG6myTjLtZT36E1ZCKSzuF29hnWLXJQ0S2t
SuEJkUjQi8PmS7gRYXiwAbnWdiR5VssGYZl+gjVTt/V2QYMXQ91eJy0W8YVRDFuF
zmwheruSAJZG4W6mRZjf+BBRZGgXjQSgIKAYJYp2N0rTqXs1QHhu3dWgVSpfovCj
uHiZ8LM/sLxYq6H+J/qDh1qHvidt8USIQOzIVgoq9+lOqfR01wIAMi07gofig75G
CydggZYI1dNRlbhkzPQ6kVxJBYJl1xuJ0DqzDPY2tBg3ecby4sP7g2nkqDaXuH3c
Aacu5YHhIZqwQ5PbW8d0TIgMdAGKk3phsjy6CTBqkpAdaGEaN9dUAvq77KjVyT+y
igAQw6BIzdPA8N51bsRgqKD2mwY/sXwek9ipcdq4a2LPLIVY0od5mLpmYobpNnvI
pDmT6l3kIJI1UwUfqM+R42lz5yD4T+6TcV+GawCwNbpq4L6eQKD1vSN46+vloJMy
vUUWdeNRJbw/JEUIRQt0j+vcvkcz65BGBxu5bU3ubOoatDid3vBlX8x9LjUUz8Sv
y9fB+mquglDm+jl59t1AgCVQedds4VkSpMr5E1QFa1lf14em35rZEKYXqQkAsRs0
kyqsgoDPy8NggeLP06LM9kX3gt7JyNxJ3JZzSgYay0BdlzQE+qn25yorfDH134su
HP3Rel8aikajhibTyeFN98JUtD5Wz5lVUgRu3MbSWogh9K5S4Bc1Z+cqSk2m2hm2
9NyXKJYKpT7df9oEjRInfP6jwbc0A1x2J9orpg2CiwlBgxYSnhsCUZiLPCF3sdtB
4au/cZCJ3mbhbbpmfQTwnt9YHE6YktVkaR1NP4QENf5HySWsgpqGtqFdkNhd3H4e
JkZ533zdgwMjco/WdRQY/bwmrJqU8jpPtJ9bod/xq8nCvUhDIr7msFT/qtFPk/Sj
D2r7Lqd7ErgU9h3iP62JpFdkAbXb6a9k4S2EMRccnkJdQCRjVVpho+Bzq888eeID
AHUnBGJN7HgWV6OueNzGr5vkwEFgIUpQB29Jkq3RFyc/pjEuGwGySbongNU/JoBb
yyPdBRBOB95ljt1fJgEFUO8S1sl9b0wVirITAlngR74vi5idNoRAv2p9btAMoG4E
IqWKGeCS6e8jbAIzPodQrLiNSSIUIOaePOlM+CQW8czQ+CoGEZ0P8jubRAyFtbeA
R8py/IhJRYIyVAbAE48wIOh/a7es1UTfRv/cON3ZLWHT/t0JMve8zqi0Lcg1Z5MW
A8HyJ6FQUbjChNhRk8j5uRyCJcVOCh/a7J06fXISkCdOvHEDT5jMSr9CtdI24MIM
5qQzEszrnInY93ud6bwpugH0fNtMcvclcnMb3TVuzCYlNpWY01T4Q3gYxDMRhlmL
nL2PmKqQST3UER3KwIW2vSlsIpA1jvr05u4evcnVFDv/uXi4W97HZMaD+5CjRC9h
UUu2gaxZYHU70rnYFx2AMu7ynep8X29r+5Snzc/wZY5oCSnA6mvROyzjHu03SDNF
Dv9bcJxNZJEBzYRtFG7/Lmx/3vhwG6OIsN8XsfBxO+gIECOmnJtkxXh/PnHuaE3T
PDNzqbkNeW1wGbn/L/vqOCaJZlXXqPlykPW7odFmjM+dr9/lJ5nNl3Y7TLPwTywR
uNJBjpOuTo85BOfUeOZzT4LFBshmgmzn3V3n1Hcl1ysQYxWZKSVKPIyHz5du5XDl
GsNH4gl+AaTj3er6x6NaDCBgAOrgDi3gS1uVha7ZLuueepSxn7SWYpVyUCZ8+w+U
qo1IKKNtuCnWK9EL6N3NhCTHFr1MnCdthdzUpKXl6FA9Lh9wyTR7c2RTf/4dqe2C
rs2ekKwTvxYSBxpw0FInwhSlozGcbMZ7tl3jgg10eii9FsQoap56YN0onZtNcTIS
9rXZxE23qsCk9rGG9hD1S3tHElY7bSHUwU1FedVUR89dh4GyQm60/bOAtUbJlmhz
d+AIfF2gufieQ+4NrUNnUtYld28aC/5J4P29Tst+ulk2M+9qCTijxBIibkLyFgro
AYgZIn01nYEMsFKQ1Rw4eDQJ0TOUdLtkK22XbY1vO3ezmX/Ah+qTuq0vnyDjgpWJ
jAxwaM2k8NRMHLDGcvIy8mmvKrCqu/MP3jLjDcYzirWzeIcrxTH7i3WzzxWMP/DN
sM2MByWdq7cdP0jevFKZM7wn4RVWL2ubcBINmMdFvK7lsD4ryrnD2DTj7j5HUfTS
Vyve4xhUISteqtATEVafeLpPJQ8OYHlkt/m5DpjJJnXqztkvz/mKBIPNIhc1v49Y
sWwWnKs1ccSohwBngYZHSR466EwkwlTd54w9rDfDE3FHMP/SNkzOfrR0X4NzBV8z
xKtuYYRHyuZBMNqZgQ9n4SNeY5QAHFMuCLCnoZoEinIywd/p9o1B9iFu/uO7CmSg
FGmUbCF51hTI8ypHyJ4KGa0k3+C1H4r8gs0Jufft8Seq/bimIiXAm0y3Tv3HCF5Q
WPUceony0MPPkTWB+0E9GRslTZmZJT6hJrg330mzNd5H7H1wuFkEHuxxzHPLvMJP
DP8hE6Pxaoo7+Y7bHneQVB+N7cW7oyFPh1diAssMFA13sdMSdkIqE/+I9R/YvjbW
8knZ/CThnCbrki1iMxa5EzxJd0s1IHus5q8d/rK1N/C4zB0MSN/ms+7q+OqLvkFm
pNOUgbiW2f7VVNu+sML5Y1+JXcfdVWEjcLdCFk4RQpPVf/Gl++LdFiS6NH+cmbTY
4QTKLfmBwjmlgAzGVWIjL99nqmaf85CS1CU6ucE0SxzKIuUL4Q9D30G0YuTZ772O
zCu42FN8ZTAn7DlB0R1GX+YYKfcu42qd0Cna65mDiBBeBat4odjzhz90hY3GaHZo
PS9YTzfxyOUzJnz2/DFQpBBWsC963cXr16YBykr5VSbqHVU9S58kVjHoEW/FoYah
1XLK8Gy+yIlNSyTH+3IFwGPrWVvIyoXrrDS8wpaWVP+aRtmfxWXWTDkGqWrrwgcy
u8nwgo9M5LVBIPJoTMIYd6OE8kydp4dbIv4SKAyGtcsMc7q3amSuRwYMb+D4P1o8
VdDG7wY6hVlH2UY8riPFdnCHmzBG1D9AYTCqgU+/P8s7IvWp80ERGnRaYvOUTzXU
VKnkVl5giC8+uHg2D/PBdcrCX6AGCUQqIkDgJ+jtB64lpeqxTYJAPvxECIRoGOUy
Tx6jEucEQPwzzUjlqwfXpUTlANpr8M893dktWKNdGfLOeP0rhGkt66o0BukAEtmt
bq3H4qRI0K+jF7aZ6T2/1W+maLJKm1MnlAmT5KL6DZXbtfuH2s+v8F147ZRJYz5s
afl+cUbsAYED0uDg0tiWmPi4LG3ftVE+K0tiA3QLZ4kdYWQ6rUKnr+xFALVq8QjQ
TolMTM4+VrbSIFAUTiBF3NaXhPNqfsS8gdJ8Wzn4Af7D3vXKVugAgsEceAThZmxL
S11lhtwNsqBoFfHuhX5sKNOaJnnT9c6SAUmBE+psCgNzQzKmTInRCrcmmUEyaj1+
j5rhO/4QJz32zhxt8DNqtOm/eSVBrRbILXshmxXU6lQhBDMZCxOQ9AFRZhgjP11T
Zn/y6u731peZvs0Mr/sbyms3FBH1uEds76IJcNRx/wPYUEcuJxOo8IofBfLhkMlx
Ek3lmZ34dgQN6Bd+sUGSPXu8tQEvz5LSZaXr/3idbGcacz6AfdIDCz5AqysPi+Ek
XEt7a1RnEjNwUSUXyENb8Suf8HxE6FK2K+cHAM3/55M0dssNr+GdZU+HdY6jtnjF
XKYnCjqq4rZrxSOE+TKUS6c3OkWg59/EaYJRONDblXRD1shdV+PWkshtQDykHwjI
bDTnYE/Ue19nG0TkWzrfz5JYu3m6F4Ys6bvibpaEejJBePFlgG1RYXcg5Wv6DvjQ
h4NufXAgLb4colXD7XSnbF47XqhcnZwcXjkZWJ18L3JlodrjiKpJECm+5bmDuuQH
EDH1GQ2vyRZv4j3RiQmezUNOP5o7nqF7F66GXhgWTI6bDeOvKOAy+STBTIGDGjbJ
D48/axmitLTBQ/3ld18DlgR0u++WI1gEFHnNJz36cOEQh0FWWLWpCb10wPblH2UX
TsjLgYYMq36SHhWXeAb7SdiZOxzunoAPxDjkFaiU8EBQu8hxvkY6POWrUzswTpuN
Zj/qvbI6EWSTYRCX2mMmMe40DrM6Jz46B8nqnloI9v9ycMqwPbGu84lsC4+6gVqq
vUYSX9K5IYz55dkfqD+Coogza9VqnHyeM8LbXVvgCr506HRyq/e0Lyp3XPqRwpex
61jxXjK1OsiQcofACFOfiV33g280wlum83/zeAruDwkv3A5yUDWnsfj8kGHb9mWs
kEmZv/o1sfUZe1yXHrmKcKekRAyylo5phnCGgPQ68ExAkFsCQ4rbimEM5DxnkqTs
FLVnbpL3ZqhRbnHOprxZZKGna0jfX4iaDg3+aqNWt/ig013ubK/RJpzLjyoPoUm4
XhEXVOqwhSOFsmGCtQaGIXpzljEfVFkl0hXJK1/fA8yOTQS46JdoQuj84WOavK5Y
RNRC3CP7ZNfSK6cjY4o6QwucY97Pw2i6QWkJDyglPJyUo7j8sE8Idp7ng+p59tx8
suoaoKanBLpDlGBqAUW6NWTe1z/uk/64ByYjRKj6h0lz7Fkk4+25hf6HesMe8nst
/oRs5a+GmAWq1WF4/jrwcIF6BLUjy0qAHnJPRlgSyV7ow12pKjAGw6GYLv9XEv/o
sZNAv8MTU9E+ouG5wG2YT4P+3OnxVwRZnzBbXnri/DV0jxtJcGvHexe95f/ZxAuv
kLsYpspmJ0oYRsxTZR1CylTDvp/BLK4i0DJAnzfQ/Wa17ff/p7JJleCVobAMpIps
YDg7JMB2vCGr3dBgm/zzxtyczDqprq0uAo/nEH1s0lEwd+9ShuIL74ZnZUvHX4jS
e0RypW101418d8U9glLvOvKO1BYWQoTzD+yy+K+jqrYOnb0rOJws7bPfQ84UGG3z
B53XBF/EJFlnO0+bgl3hBhLrjQxGSJ73ufgeHzlQdCKZaz8B73qClonPYuHfcbhz
ecWz23vsJt806vaNxqlQuZAOyGoTmXxP4i+hHJImVXVXc8Sr5p7Og2H9aWGPItsK
YxiP0/Bk0l/zBBkQVmPZEo0Z4wFiqIKABD+MMsljI/rI7TXsL4XSSM3VUad3FtOi
Xei6gOHIsOdkps09aN5Ldi/32UakG/JvN6FFbtdecdBOU0MqwT5dyDJz6Q9V3WSS
fDVJMzbIP5F/xjOul04lSV+az+X0dTRm7Use3kbangnZI1vjys9Jz2Nab/Ub+w59
zjehTvBgWc78vRbn3bK+133gIBIStivFog+LCy7dLStlO4dZAij8KWBxAE9IImn5
WoPd0ixNs2NSXTxveMq36RQi95OjgQYfbztTbNVcm73RRGJ4OiMh34GlKMfNryVO
mRt6IaeKdW0QJx+U8/TZM0ghwp66KBmwq0RimYwWG3+hodrTgp26y09lfV3+215y
x2myhmnWnD74ESA+fb8sCrWcmekjYsCpsEergH2qLca8mBC1GPRU3nRsmZ4vrUBu
c6JxbzwsoQwSr+zOVtEi0C5C2DukzJEgL9LIlms9xDlcC9V03G8Yj4mDHL2YciBt
YHSslR+lp3agT8oQhA4g1BSGZ3kMqUyjX4dTtpI38bZ3r4ShPvQhfK3gfbgqjH5E
LAcPUVG/bUI+AIdNKtuwSfS15UZz8AZYCjeVOQwRUhb5KFTwYs3NrHB2PwO1+KwU
D9mgTjJkaa1WQmExAeAO4b8yzZbPo2GWODJ8QCEMiW0WJcciuzFr11cMpqsw6NTz
kaR+7DJfT1pgvluAJYzLEkEVK1FPLq05OwR0V25hmKH+/0BZ/Cz0OYiKd2m6h69O
Mu6McZE4ubZyb9s5L49ZyCaRR72O5fqJO36/Z8CykDGOBx3PQUsHVeRpYRC84tfl
iznDB61XNIv5KT4NHMPleZNXvdG41aKBcpWmZKuM46BvmfwaYKbnQD4wguyh4D/x
u3CJ1hjsJ5EaaYNYbw08pcqSeHJSyEjrACBB3DUrWD4PD5XkkDTjgsTPPZKuKJPk
3EYPBMNFASlQ6CGPG+AvJYRfuKaJgANxkfGTSTu/mcoRj9y9j+gvA89wBV5PwAEx
+T9Vylz/vV0FFR3+JxhbUJPqOrFEb2dH+gGl4taSfmemjsPvzdkf0tDDXgqQLTG5
lAnEWxzZQ6+flAJYOmeoJUpsStI4TjmTvMdwHKJn4k2oHbzwRzwZeINoddoNKQ3I
fYRgeV4QqZeuR98RFrHdWrYsIgr993cNmQwdh/G1RyGAz82M2EhATWaN/8nBIWWC
ffrbTnMTYMvWo/OBGo672CUTqWOjiyb+2xP+u4R3dWRetUzQq3sjFdDNrNyILugG
eZCfp4ecqjseSCBbn+BXnkbXxgcSmvDe7oDLwWyOx4sJhzN7CCEfvspuquLqHBTJ
KpBskrP3Bh3MEsAEoxQTFZ7aB2v5N0p6cOCZ9I4Vw7jkjrq3fB2xF97ATtaipb49
Ez8ZX5fmg8dJ4VGeQ04FbFV4fEyj3sWxFtzps+IhTsAORBm7xvWxor4gDYjgIRnW
IZyZMy8t2lZ4tH/BnME5Wu4ghLHPRqjD3nH8mv2djWIfUiOrL6cSmaAkvPh6Saja
8q1MkoCDfjA1plsblP54TGtjyePcI6xSMms2uw2OS5nUlG3J4kOeX8kRYaI7CLDx
pZuBiwfDW/W5bKGfq6fV/okf5XwBaZbprMvJ+y5nL2arCmyTa8Cd1HSCvExrIy++
mZVc25MNXMv5Nz7WRkGp+eyn2KatZwiNZvqcTFNHpq5IFi8TK7j4h2toXGIW7oSS
RoYAkC8waHizC51v0/4Y9EkNbgwYX964AJZgdajMBNZKVGX0+JoozRtbaYpSazQs
GiJpvvNZOI2adK5EUscl/s+H0NBIki4tpCbNQ5vr3uOpXlIshVbUYOWAhEiaRV4V
pZyLZj5CWvie7B9up2I91OjXkb9TscYWG7M9vwv+89tf9Z1TiN9gYuL/M/D5bN9C
XkzMgoqF9tRny+ZWuBqMZy3KO8T2x4Rns2U4ZSE6TeQv7fxjcgP5r9/9mbhVhNJr
QshUohQHOTQcNVhFI1owIdi/kH5v/aW8OHJl7LpvUzEEPQOCx/JTvCIpH98cW25D
ypsFa0aKWE8fPsfmjHwRNCgYFjGOkomdhjdleLWIYdYHXet7HA5NiptyivrJPIEE
LdWXMJPnIRD4V1x6+gpLISr6yCWm7/zeexjeMv2WTr9g8zNQKjbDHZraT9H1YBT3
XY5qv2gZ8GQCTKiZp3bp9MW0zahMVURziFWDDUxtlb9agKehjmn43fB0P0S9KXbP
gJyIIOaariUdSHwcmoJJBBvkVXEo518fDkgDLKpp+Jkhklk7/ekAR9imVf2B6mq3
2m28E9WPilJnlnUlYCPeppP1alXYFYjaMZoj6MAiMHuBSQTkJwvJniiPQe4BCdPx
OsY+k2Y/E89NWLNHB9Fn7SDDFKky92eG8EGXhlowHqVHuKSGo6bLye5qvPMJVQUc
a15C/mAGp8xy45wIs21UVUjqzVnZ7+YZDGRU0q/d8a4cTFhWTc+8oPXDb+pCV4qX
rQr/w52/HVnZPKLfPA2CNdky6MgviIsHJaFF9FcI9Q7Gc2aGgz27XZoufkT/778m
H9n/sNQ3w8J0+m3l1my6p3oQWLTmdVMMzXlASrhF4TZKefJbsSCyPIBcpE2QLZg6
bmqQMjn6fYxekwOIeYge62pwZ74HrU7mB9FR9WACn2vk0nAa0OPqytW/7cdQHdEw
PPXJ3UJY+N7WqWOplxp9xXK7UGoehRH/HNC8uhhvOTdFuKfwfydzWqWbCNjqPK9+
ia6TpZHNX4WHK3XNdfRV1q/fYDjXaZfmNAPuPt/zG2Z+WW7BTwQudalgGSnH0s7k
hSckbRRerjFZlcUMc4gX1VG9enMQMKGMCCRH9eKGJqRQCbYTq9I/3LT58Pwn+ZbG
c8Zb2gsCDrJc3PGM1Yr1XdRyW6O/QZqDC8YCOpxMDBKIYEI3tUOqkAjspH+Ia61R
bo9jZatbvq4mivioSCq0ZFa49mROVis53iY8SBUpeoTWAnO5Rp4OZGMcRelBamg2
FgRCCfN+PnzytlDoVJt32Isi/s0FTw0clXrSI+VuDVWStX4fozGJsTy/LNQf5Wiu
uZSYn0RNXtAHbuSuO8HSxWSBa0nQKPDigVJtgOU6dfdCz1GsC2PDhWLIMbcMT5tQ
TGrHyqYmSvuBjokKsSm2ibGRF5ArmujA9FTgHnDKP7WVA68SycXBt9xwDAPZMkSj
ADmYbLfiCJjD5yqA/lKesvovG0JQxzKOYFuXf4dqI/YwySFVPnh+QNtLT2XKfLyp
zM+NBpIv3nKbr1VHkKJ7I+3dsYCe67oS3yQWL1x/yZTJsSm0z49ngslGfBFdMsqW
txipAVlkVG5PeCT3IRdgJCMtRlchf0GABF92y540ArBosQaY6mSdzA+5UC3HBE1H
hpzVDih0b5Oq3a6lPFgWLk7iU2BIgsD1MDCe2vPcl8hzbtXfWe6yEh+5T9Z2iv4p
+4lM1FNPlQKL/mVp2nJO1KjORVtOXGBvj77f2XyJ2KqA+G21o6yydQ0p4FqXsu5c
8HcbfuyFyII4cxyl8BKSkZDGb5QiQManWeJgg+eQEpW7OKsErPtFMcgQ36lWO1QL
PyVrdapzQ2zuPsgDlxT7nxGGJtOxsOVkrCB2obrpqHODs+V57mvl90BdYA6WUxOd
RREDCavayTx4zUndQZpwheXdECRtC+pWBpbQ27Zy9ngWvfvT1W54dwbmZKQwyH+j
50+1aD8w7yL4qxNV2HXYbzUrh0+Gq/9yucnbk4RK6bMHUlIpWjwz+5cIB8Di3FEN
VLQbNreaR3WbiwqsC2iHD6FseEo7OFBH12CIW4SgJVGeb+p2nV7wRBCUKrYlRpMK
hHPKV8W/LVbc30spp2r/h4yGtZJXzXdONzcxjszJcuXJJejvkty5Lzg2ioi2xulK
lU0kBigADHr/4GXr2729Q+E6iKE/GvB3UJpGhnLjohQZkF0bs5ZCH3WygsTt+Yc+
T5NtT8M+xbgTCBVeaz5BKslFqkiKMbCApujXeNdH9C/IMVZUr7USVaZg94L/8OxF
f3k5KoczuH6z7MbPgYDJAbQ/iSTRAs8pC5yRCrsU+yYYRAMpvWICLSKvVqeXmbR8
HJp37VN4lSJlnSEGYFOaRGPCMW3L1Fk/DzRfa62lgoaKokgpPEJbpQT1GQZii4qc
YQ3FWtHMJ6zaqQdrfJDKVMJN5H6R2+MqUCvjqULiC+/8yBYYL0AVJ252QlNlQpms
9SpqJ2KBMUn8zTY9z3T318+hHPGEaz21VvbsPnWt3O0HveNqTz+Pha2CDAvWmgsh
tY0fTDxP1VUuOt2jv6cmCvhVGvQww04Ea0yfR+4paaD0ZrPsZmH7tgYh8mGWRyNs
g/WxDWmkMepOlv86usNnufXKpSLNPSZQJgWeIeE48d0OV2JWfdNvUoVWsRs393bN
EeXjtepX0hmhHuWudYvd7c0+5i06vBW1jmxKBk0hZz3J9IOryy3WhsvQUfy/LBBW
YORrQhlvUoGcaUlBKb2U6o1iV1QpU7gkvUe8v+0J0ml2iEe8dFLvAgQXzPUOSsMA
M9CkyK6LV4Iu8dSnnLT4OgRzp0l4hYspay1Pfm6AUgcR6UiCZMr3MkzUpo8nOhR4
axRQ6e603srvvI47Pj/cv8tdrc5uTUtUVIO5u87zHF8t6ShHLS6X6NY5E2kkz0hj
nhybQoQs7Vot7ETRapg+xySfJ5ngzcFyvT8+Mu/VJax/P+LIcjkdLAdmw8uOXvYH
KQHb9Sp/gL1U9yxljAqcooQZLtG7C1KyW60x897JZVOkHCgdajw1n+zxACXSwNHa
qdQ32w6U2zLkVmBog1AURTc2AV0eew3qc01h+JAAJrmgZ3g5e/9F8NWPFfnfgDkr
+WDQBY7n33a6heoLZRsvacMw849PYXEJR+EZs4+ZTllOLsq8k9gA5e08Ajb4ka9w
Edm/2YSxyzT6Wm1pfP3iQnyFCl6Y9EQKGooh9lf639MfUNLY22Lfy885TOfxxdD2
/L6tolS9v0CVwxCVaDi2J2nMpoLsmZqV6cp8BOBeZpf3QkvACnNdbv8CxAQoioSu
uVChkEWhsnQawHPyJC/D9cVYtT0j5r7/VfgH+Hm9KLPCQHtqdAoLsCGXbRodHQiJ
RcDuvW/ZXu9dWrvrorbye8EnwlbUqV3wm1MJksjhEG87T66ES9aKOsIz+kDluaH2
WyntCkjgjwUhRUbadaR5Nv13zMneJogvwxwZ4bZhutJGj0OfdOhn16Yhd797b0yn
VkN1IPatE0EyWkHD7mx5fwPkRfSvvSL0tMUOJjnP7ehOwQ2UpAqSQXpEQcmvr2Ai
xFv6uc3gzfkwFJI0jT7lj+J4rt6ZaRgip6uwAZ+ooSpZksVGG0Ney5+PE2ctUC/Z
/h761B6ClQFOuKOxHyIu33Wimlx2GBgZrWa8/EteC1L3LrK4daS7Po36UQjAMU7K
gBnzCEFptsKgiPx0b94XlRdtThRwPf7yEwFdT8R2DB6B5ycrn54SSdZ/47k8vqmH
QHvDMz2REiMKd4S2FiWH2w4gaW0UVH0dULSN2WisHPCUxnZ6FI8/I/J155RhuoIS
pJMl9meWPIxzBoOny83CPEnolTw8rhVnAnv3MCGe1OAlgZnh0B5YRvAZyvrk2KgW
wb/d1B032GdHkCTw9kIdQsKhHj+raIj/PlqN9Gv7UhI7G6EzAR/wUnm4kL2Fp7rV
18ZrbBGXrA46qlqmcEN4RXykC0mNV1AE6j8K9L5aUWlcPv0Ybx14fBnJ+XwiNgzX
4TAZcg83B8plfu97od9Qu2YzIdNdx/5PWZtPUPeeZtO1NFrpe9iO6eRcEw82Gmsc
HM72dGkg6dvHklis0KRWzS4JobCxtfeCAiU1rgtySiETLbOz/NRbq3q+vXPokGQm
qBW3sIwoq/ZibgMjFDdByZabmS+dnBbmmURw5ZfkEvEmMqk0MVLOt9tvDfkmSLaU
PfkjFZGz+jCmQeggfUqF27DqwLryEF3ZAmXy01FYSNo4lDKrZROUlzoipTAwxMEU
fGI0gGCLdAEBDerNA4qfL1o8MfBnfjo8rDcSVcC6mZoIM9uF+EjO9pKSuNz9BusO
FVwWxLSO+fxnOMM4wwTVMyUtaQachZncXMgmrtlrTD4PUixGwVIk2CG3ngitmy84
9WHQnBY6E1ndlRXxIOmoWxZczfCOZcb9DWj10mkBzC4Z0HV6YerxAopaG2i9tybW
EKYWzbhH2hy05qcB8Zh33GKTZgrxRl0P5+TaCZz6t8UOByV5XrA/hT0TSoGWCk0D
jzCWaltNMoxzH4Q5EokZk32OP6CLRgA7nrD/sJEEZ44+MpV49AC3SokmhDhJKC/J
wSF3hLKXGRAgLYMphsJNBsoCeXEzaGnaGFtlAgCHtacc8c68bE29LQ0+i9s1Kgvm
F/FuJXklCYm0SK5ySvFAApB8PrG+rJ4b/s8Y0uNoMZuA4UiW37a4furtgUu/qzEc
dCSqamm8Vtorv2DYq5KQcMnTTP0EHrZiU3qvt/JhYHcZvRq2enURo9k4jGV3hHyr
28BzhWzb/UQQNzkxOTJLlN99VUyJDmhh09noGAQ2cBRBVx4Q1shvsonekHRWY1lE
Tli+CF8LjzGd7fZNGV1Y+hzpqVCD6rrQ3owB7mV1r97tjlsFzLeLRNWu0/gLIGm5
rns563BKqeS0fHlbbe2mzKazcpswA6OwQO9gtHYXj28AtpoZfzyR3viUl3ejzRwr
FrK1wzODU3/UUoUj9dl3JqSMMliayaaedEIAOjKDnZwKNBLqWXce32qtcwLfPPHZ
8+pHwVsOQo/XKLYT5Egbd3rDXfLEosaYjLaptB0Wt9KgXsA7vspznNxiPe2g4rH7
QK3IkUdO8GS6mrX32UnxcatrpGm9JlTiVwU9re/YrHWDlNI44JMqkaynjuXgC8P+
olWZyKD8SaiY7NI+hlfHCElkaZReZB6o5pTiDClZN2jsMiuzRVlMEZWgN3YfDFtM
XE86uR5P5oTJ9qLp5Dd0HxKBCDqSiGb/Rm91sSq05Krz1Rm+ZA9iS9iT0P4V6xRd
a44mF27X8d6+xuCmEyalC+F2oFrxXIj/FCxoj/sH6Gs74k6uxnRx3S8prZ4f3ypo
sBz8wuKSW9fcl0ZAnDcxybIO6DBs+dYNezTY2c12vrch2PcM6FZwsXoaelWe2PxX
d91bkneHsmWy3aTQwwLEc9m1BBukXhORUYlWvQFnf4vuYXHxTHlMNtKb0f7Iw2A3
2Ct449CO5OgwRCBlKJPgLy/O8/I/iKRSn1bw8RiKNaJX8qqYEaGTrI/53m1o+yrY
cmUdFMu0ZHcfGxNBeeFlcbfestofcKjKbki+2rBWJwb4AKJLbSoBj9u3uyViXfRJ
k3dPSJZxMu7JSQXUsr+ezCs6b/4YuO8zEY9pAdkYwPVE7anRHLBIXN4E/iMh3veF
xvPmqyAuYwqUkXqnJ2Zwo91rId8/uLyzKQmuhxVdA5cFXqHOwfEHYTLvr7dlPXRQ
dFxkgtWWa4SZRsSiwSYs2Z2jN9OcAyne0g5KzQKKWbf49Gphv4NG8PxTUpo/nils
0tY5gw49rgnHlrzQWPAwMfpr4Hlpm5mOEpdpByXecftba18LTDSFvB1aJQ4ISE9t
fH5Z4VP1/4ejS3Od8GkVKfSUE1fOzhi4LJC/PjyJx7sFVUQ4Os+QfP3koD4DSvt+
LoQ1bPHsk9tjculkykMNJj3dXwBbXSfgW3SFOwc4N45x62S0ITrSxbfTcqvu4awQ
ca5N52Wn94PFkR8jze1X+vBSjR8hMwKscu++51VxYvLuHBt46DFKWBQGJ8OFOCwp
AhD23LSLm/XtemfkVpmgxi4v9tTRDb8OAF33/SEVT9nYzqMRwdMrOQBnQKZhpvI/
8XAQv5jVl0AnAKkVdhG6/nWhoaX/3Nt9ADxRcHrE98ro6QEsLomCR176EAzP4nR+
yQU3MX6rEKRx38obF27JtQSBiHDJizn7E6Ql9OoLLtREpQ61oByEyp4oG6fO2llP
xDoKJFt2RlUC4yyyVnE2ou3RLPOEBL/aj5WLzF3fI0FaRWZF9LncWCGxviJo6K8x
BOJkJCLXt+7Iua8iv0P6jkDGWGeHNLiOs7lIGWcwrGRc0SeKf3P7DQEPBE5BAYUf
u0Tb9kRemcQdFW4e4Cjd1dLzzIu3DXOBOdh5ozlkT7PvbZ1SDB2HMbNdwf0sRmtD
FcPP8KiBxqeOEeQiZFnskBtwC4CkLzI5DZgAfgeLOr4DMM+Kjy6WkVrZ0j1/AD9Y
gGjjDuGp4EFW4nppQtgiDZ0kIUYeE7FD3CSfuW2CIx9kLG0i1yRdKo9jLb4NDE0Z
NOYPQWSLf61khX7SShlnhmEiyvjxSmn+xrmrGoFvLtVqj5ACDLPSZ6Gv/cA7bgyD
744TbHmAUB/17CuFBkmutqTUdf8slNYihc82cXZ9DG5caULWYdlbDO5b2lhylN08
xam4dCJnfNSVCzFdBeArwlAzMKF5Lr3jZ6TT6/Y7GkShwTZ0JPOD9lPAhbpDKQiZ
+RirZqMXHuNKEiJwMybfKP7tMWdXNubaEsnBzlUneM92l/3wBQqssC6JkM4Nt5wZ
DKCX28HnBxrpkfPvxleBOmSWDcD+M/lKKfrNe5D3fFZ87Y/8rf+s5IUYHbSAT3Pk
PgVl8iCL9k/WSiIsUkXOhHVqBenqCDK5Yqq0Ei2z0omfyfoFaDIcjfO5UTSDmN2v
sb5/nYwkZ33+6IvRBs7ShmdHKwvyPbIFNTvfHlBZBSo/nX/mE6wKbjakwm6KCB/J
utd4rA9q35mPtzG9uYDtMYpq6kII+EbHijRQaHJy3luJnsglz9l7NQ0WXcRVKwmc
3TCH88LCYLC9M1zn961mCNVpNQOaJ8RwV6DAgsyPpPDgv3wzr6UeO/Zo45gbTswa
rYYlB1gBOBlsLwHWB9i12kEO4ey4SRZc19ZrVYy/MwtuH9qrVaT4o4QlRxdYkcEA
ylBVPAdb1DizYpkd0TXc/mGwp66RAqwFBG+jH73H7S/CEACekXR9KsSA1yMhz+4q
bd87NqZzPj0GroLU3VfouPn6ShTfYtURdxP3ndu0XTzDwnMtMICQsaHhdMrGEV5g
wJYBBDtTfKseEHvXtjRp7YDFX5b0i4ob/7Y1gq4tZXKp5ggiKio2prih+/xSE70g
RS7KjG29S7jXX9zjjPNuBUaaUv3kyt3hhU+IHpWYrq1CrAKzT6xjrQioZhf5IE2V
UEYMVVn0IIUVy38FhPEJqoefi0b2N/IFn2nxmQIe4x5YwfOIXZY5NVjK5BQdtQN3
YrzdF33z1WHt6eobZB9mqjsW7ZQG4serdjbgb2naKNmIdTUG5c0b7ET3P3sJGsdN
A9q/I7/daFq7v9feQGW5DFi11PkTkncX62Zk0hF386+XwiBihZ3carP6SyHbHehF
ZyUePGyM57tjaD87xea/E5gBvXQvAFr7aBuxW9s4lmo0eU6ABWcMNSmK682PmuTz
eRH1Y2hAE6OW8X7SVKd+osrHsylyb7pcOeh24wRQF73hGDNqqnKpKCo5ewkz8wVK
C0A8ybxJ9WUa9D+1AVEOrSitAVZTc0yT4QGM2uUK4FU3sKH5X9YfmTWyYVNoNEVu
MJoA0EppwFg7ekJdxkOgmTAFIMa5vSs+W2W302WkN6mQeT/dFjF69h/W5KKMA76Y
DWVmcmu4+u3FV1tpaK0d/PpYqeTZlklMMd8332SrwLIO8C4/unfCTBEZO5fCiOPc
HQPLiK/uAn12Y+JrlmV3Yf2P93KiAmKp4cbHRh4vMbRmv4EoMcd5wqVykaR3QRdg
sUskaLkOMrCms1dDLPtPk0k1tjNYkQ3wNsJ6zToxKDAXDv6Df7h3ZPAaJU20Nu0N
Se8Uek9BKHRiZf7auaWmk/NAQKht2czmzQv8PQ0CdrvPV1wbjXjky8NpFKcahKce
dG6w1ys/8S9dDkdKBU6Zc3YnXx01+xqk+v7HmDFgIeCyl0+nj7/TWUifeIZlSFD5
ABy+GXwjvsR/R2MNk2mhjtWOqjLakuluZfGCuZFJ5jWGOuxukRhnt28acCMV8eZ7
huxzXO/ndAesiPRVW3M71xp+JlWdSXon1mHl3cHmgaFyOFnvwd7ZR54IeHIiDeDi
QA9kfLBHtqXGGc+sg5CONKpIO7rhaHH13TmuscF1itcTIZSgaDjbHGK+CY7r6pVV
XvEcj9TkvM1mLoAqEG8Cu3JzLhTWaoBKk+fRVIp67FfZ8eR20wDvN7pM8osRxVmc
I3srUyq5Qh3wu1GP2w3uonXAMYHJwM2O9X1JOJ05RCIj76tKUrgHoNUNAEOzdFzM
pKKAH8/p50TV6pAis4iVq38h0Ojj9ja9LD6CohQAcAubvN/e8gt1WrqvfBTdTaUb
djoNSNt2sounm4yGkVnuhPJkhBcuR/ThDenyPCguEVQ1FPAlQbXlab3S5+pAyfu5
bJRZYAAL8Fzuz4pInb3qtR4/wnbC4L/PMQF0g9Ql3WlURFZntC4FBjDjQAI00g4d
5eXpui6F64P0hX+ZcQtBr5feLgvrCzGWUgEU+3sGN6e29E0xq8UwdSztyMlz0+SH
jSONl1JCrJCiND+b1dr+4pmqoHrSfmEqoIdnqjbvwnDCenkbfsUxE8JzfHfFF6CE
QZIVPTY8fAv28ILEigTKoBjD7JfkfjAPpXzR6lQNBZSUSKOdpCh501/l8IfJ3rv4
tp+3AsMoEiuaI9NPDjqeWas6npGAlq8DsA1pDm7im2mxlLsexsluyPJHXFOGcN/w
HhEJSvV6eh7kKRp2gpzuEA2JMyAIWL90Plz07vHNRHxA/4BBbJ2mqQW8eH1HYeEt
/zzLbfmOJPdwmbf2Is3LZtce1flSFyPpGFBuC+rLclRtJi2rTC7vrEGv8U5C4Zb0
oCJj0j43QOa+/wAR1lvB7jX/CmJakRt/2HnrqAJr98lNquVce4SP5eziR8oPKj6A
UTdbciItvgjrqJ1S/h4PBbmsc9u197mwXPg9FFdJ7I5u2NQJnrb4fBgLO+Gxodj7
tIBBoBux0nuiXLyJKCk7CCwSF47w/vYz+QTQ2vBvasnWuo6zNLYIvlmVwT3agzjZ
FyEKN9K9LXIh6zCYWIZiuxmADK29bwzF913jCps+cYoNcve2MpTZjIOVf04WCfSi
sC/61x8pfG6tKaUOFlZ6OnEnmKhWq/wGQJS+hbvwa5BfiS7+U+Wbtt6xah9rj4lr
fPL1hMxtrkuJyR/NmZDPCCClxoubm0J6H8/ZfoSgxOkNetnMBRzPK+6uFRPTKne1
gofAZMqV1uIcQMoo2zT112QYdmUdRdfUJ1+iRFAOovDqusp5fIeodyu+3fN1WWGI
8F0449k+yuFc+ggF2RqX2WdV4jl1ITymqh2DmYGIlTixv7BNHUoKXTHWDd8KYAzJ
Ght2O43hXuUWvIVsym0Gkx4nNIZud3ebqRsywzvE8fiJc7fIA9YqnrW/jCmS2Uts
mDuK4pSAdQXcZ1tzK/34Dzmd3TobBvOflth/9wzdovK3jRsodz2zN6CXVGO9dLuG
hUQ4/yyDBG0P9EOQ1Ti+/W1TiBf8NV0TqTWV+7sVLU7JBLQ009eQYvN4X40UwQp5
gmoK1hxBPVvnYRjMWtKfmi54zAty40h1hC9hbQFGkZBhLvontB4BO4TU7I9Lmvag
J8pXIe2XwNJ6wJMcoa4aqp8eqbrMLySSoAlkHkVG/au1Y2i6PtwJvS924yQ9E5pm
3gNDKLWqCbnPwwihHejoQjJlOZzChdqoj0lLlcEkR/4yKjBHuhkqk4Mgp+kYv97I
d7etArIeFPQE6xr1BKHKGEGv0hqlGzhlTL2WKcsxr53oTMLurwDv0BX/L5pXU8wV
U33FzItrVqp7TkzhKQJsJR9ts8hue1RsBqOErcLFW3owZQpAakdB3RMQbBqZ0xQ8
kqAi33YVrSAbT6o2ECe1IoAgUsUNJJpFimfXL8NhO/GT3rP+nVTyGgJ69amM03dd
m6A7XAl9Hgqb2emU0ICUlfJ62h+JM6yuOW2xf8CEp563TMonWUbld5kDIL7GFiEj
+R6sZeAtIXaqX2K6A/KhOVtu2zVk6zp78hsVqaj0LAKKcKJWd4rCHVfsh+y7pVCx
fWaLAcAWOJZyxyOiCMmMeteFgcA+XbvvDan4/5hkY9lHc1Qg5tvgtu4VEjwP6ea3
pEOSD4x3g71bHxE5WwuqS/go3aNSW0v2pmiEAgRQm9vIEFswkIct4HQRLQworesm
VsnqJfde2+uJkYR/2jCXpOLgUna/GhsgBw+kf2HgsRc97gfeUlRUz7HSoYqaFAnz
OTGU7wwjq2Uga770en6XWIS7t0dmG1qXa0/5lJY/zKKqO6ufAC0EZAkdXpe8yIYW
9GKA0TGpBq0iZW4M9BDnpmsEMLn8HeNF5P8eC5rTc0GekLoiUuLUyLqEjOraXKk9
/868hnGOnTDISb3zEbGmm3Jb4k6ZUrFoUbusH3t6qRj839OWQVRQTdypJQQXIdnQ
VW47tdTd5cTOQ/X5FqvfvdPF1p0NOnEiIori4D/NOXeK2xkb4PHxyYKjtRrlJriw
JEetgsMMDvaWYzsLdc4vvi0kb9A2p4+tD/mLRFowbuTsOHFCP8+/5Ic0HBQu5ddX
UnO0oJUx5QfuGVzgtUD6aIhzP6f8hJtTiOvlOmVafJEX/xeokMLpQmr16h57JAnF
DUBSf7I9S+/ybciF6mcWpB9nRKCCg93HSohf4z+x0EKJSnCe8tQ6SQ7nWuDw5BMO
fQpL0PwnXclZe2nOC1vjIo9xs+Cb+imELHDsjKOco7WmpRS0IvxIJLYLeMnfmrKp
sSMFdINGMFINkJFqeRR8uP7fmZQ+ptkqMnkAcV/mUqwzdo35QIFHmj088RS8NpjB
WpMQXJz1B45806VAa0WkFLgW4wXjjVkpH8YySuVjlWViP4nECN9ClZYWqSFforRW
hGxB3A6aZ+PVDJY0XsUerCmBkSmqBr7XilYTKdu52IAF4upSBGtgO/VcShS/HhEr
v7fuZ5ysfhbB6r+fw2bfne7R/hZrbWTfN8K4M73Jj6zLcrZ6adGPPw9P59AYxlag
qiRP2H4Yn+nSGIEkQWikWWts036O9TTAFnMnF3BTnuDgADOBQrj4WdC/io+dPmMG
tC3RznQn17Secvp4B9vWabVhLLNemwKoxNW5ol263lAvCv7WXt69tnMnDURB72x7
ir4+A836yopU+Zp3MFXLMVE3xYUKFv2W+SpYqoKJzCJa68upO9QiPpFNy7rLGZxO
J7qclHqowa+YQom4N8w+1kN+Sub278wZjLFoMxpkLc1pBCCeyuYJYs5Y6utc0PmM
heYkmxeQynREaBHhQ4lxgdTX4uzpcn94Repn1h9T1mcWPktU5V3BzCaFMz6rrCD/
UMf1GsMAji/CRdpQE1f6hEeAN5Nyz0iOohGlbmsVD9t562+dtHLHEJbfDkCWmwWF
SPuIRgCuLD0lAgH3UBIpdq7JLizPAycQB91hj7qdSPqLZuz7bz9MnB7dv94iZQ7Q
CitFBqpZDCYbp2v59wzd7jbwDfldR9lMWhhbsGOS6HDwAsvD2iVSQjZkjMvkinGa
g6Q5e0o6Uey/Aue9XbfdraXdyp1+f8wAupHtjSAGkIMK6aPEiDp2AaruGkdAosJY
ctobXNponjv7cgjabYqE0gvW2mwTrwejx/pBaf01j+LNJR4arWnLubvYwdNy7kWB
BSWJYoNZokhpKi/hKfi+AZmvMTa0Aq8OaJGo2+1ojFzx5Q5TaLDUMhcuKWwv6QsC
/D33zzB+CbJzCCp/L+TJpfbNswxjsLen+iVre6RhjM30x5nLN0D5zM2q2AODwRgD
u9dX/P8zK6XdC5MJ1BlraqiwMJdNEfjkzywgy2/pTW8Pqa8Bllt/AquFA2FAhk5U
oLTnVCto9HHij4qfFu+zbz9Uop6fo06pkylRCtC7BWdjF647fCvd5IeU96PfyW9h
W4kB2MoAkHsUB3fRLzZt2Gep/NZ+6AdI2V6AjhEOZX9nygq7W5vOkB2ZWOPjL7vt
tTHAlBCaoBpXfGQo9zHhiIUHc80MPUlemlJDMiBgN1+70uQNTU0fORGuF9xAkiBk
KZ4x5rzIoZN/AOjO4uXLmUBOtCLohjW+k2Qt/Os1AxfYG8Lt4fVWuSENFgINPJrk
y247t+3rTdZB18xfSzmhtjI2B+MGehRgf3zFsQpeY+VQBh4RidcwGUjLrEC2iEsV
m7I2rblmLLcEGd8aDh+lDHi1/pVo6CMCRJ2s9SLlr4f69FiaiTBxol7iQuh04+zL
6TSpCc9Eddlm+Fmys5svn5ZAnVmS5rFN/wXPtNVSepTmNr1icsEgSObkv6dBODpP
IaO6BmXSMD0UrayEHLn90BJnfIKS/sp/Z/ONxZzwsjyAmHJI8Alodw9JvYdRsO3x
thtcI1fStesCtFbOT0XNingBJkIWps+PlzubXObsyJ37mVVEHfE+Yy0lWsLSjPc9
4YSQHfD4c5pRHyMFmvzw7GtbhYI+Cj3kcZBD/DLhG+Nt11l0C5AXTor3C6iRoWR4
HwrjhRGs/GUvcBG35NXfFTM58DUc/5n47HLuXfDLSobkTj9SJXjzYg7QDAKP2m5o
E961dmzhpKqzLTZz+ISlAekU132D99Dd0PiWcOmShsGYd/J1cVwwkmoJCl4lzljF
uoDVCuXSfuhvt5dvD2Q5OYlWmlELdbLaxNqcIY70KEX4qpEyY8DPCnM53KErf3Sv
h3aHRfjE+FaJ878KDi+r4hvrroBlkpElOkmDK6R61BeVQ5pcBsijdGurKP5JUDG1
6QMDB7Z3PbF+aZd0NGCJauw4gW1OPfw9ZAJGpNm0FLrVXrXFHH1B7paD6f7f3hYb
Uz1MRNiv7k0ESeYOlwGWFA6ab0+pIbw0MrddqeWXlXBxKluVF+YIWyNWDv+mvivT
LZ9w65HOGfuJB9sEL4G6Mhs+piSlSG/b3hIEtS6M39WfdrczpB9A1YvCLGxuYM4B
GVtnv0PsNo4L3FXRxkszXk5O4khV135T0nj5dUFRzTZu7Ydq9JlnOIjySPeAyb+F
Z9jexEHSblgtHOVkCiOYqzVWcTiIHqh4vVXbfyCuuee+JUoV4EInGcwVbyk5alDx
en5wrvJecs0AL6ByGJHsYstAD2lN8UecZL2XT2WJoqU46ubKIu36Cza7B+H4m2lG
1FhwOpUcQVA9P/u23m/HRZSR0NJ+0o0LxJFpnTRz2ndSxnfRYH/CNRgxjgAdG1aS
5r2wXz0aHSTHA8hHFQTGdT8qqmkFHiwWvAk0daXQwKi7Y56spCGiRBsVF+XLNnEh
Q58DBxTM9r/V1wj7Ho74MQz/LGXSWbMrnN5bhuKtafEc1dfcx/c576H1dFzfOtxD
Hrv40wR0rVK3dTuBRhZNCYZElrJJE/ZPYwQvk+eGiJQ3JjokCB3gar/EcnVXKN22
DmXXb8iQ8p3ocuCJfXhM6urr/nFVPISybXVccmBS/t4/5iusaNitfoZoRG+cDd1l
9L/PfORpCvg9wea9bU0g4GBcUrh6w4yX/TzGwfh+K/KbXsNzqvfVeheUXsRXSluj
Y5eGhM3CLTdqy2ZDLbLK0MmnAtCMAgUK7wgSe2H3GdpRypmtXQm29v3nX02Ujthp
tIr0UYEJSm2jQraaFgOflRfY0J/nq1/+rKBg9+fUbJuhS+ih6lgk0XO7iNmX20q6
NA6mNigCvQkn2MyR+MqzWksGACOMoqNnV/ewS/mg+8DutfnhV6qgjtuUi5ECJzzg
xZHZ2/pnFVPs+FW4HIkoq60Qu6pHaF2tI0GVoIzYFSDkWDHOsPdk6JAKYuBaIfz5
3lqu27B+DM0woedIgAlmglD9ZPld7h3KHr3dLz1aEr2wYRm/es8ObiejPd8Aysvf
bsxJNihPPmdJqU1tMmH7EFgk2plQsgEY1pm1HVvIpRYsfgMKdZ3GNfbq2EBnUlDq
bmmMaOG6AntQhg23koUV3fdBoJBGIhC2V6UjPSx2/pTLE3KiC9wIg2F+6GN2DM6S
XO74ZCb3BFakvI05FW2H2CKXehrI7xzzTdBck8ivawX0CLI+AY9Xrj3NXLQoJNUO
DYgRhFfQKqIS9BhC4WZiDsHLpaxwsCgS6w1LH7B9d4GvVuLMqCk5VPuVl/EKmcpo
bOwG5tVW3qpnFIRiQk96U+BeSv0QgDG9fQOQmR9YwvOEvkdi0tHRIoz0ym0x+OoU
G4ljZ6Prt9Pm8jxJQp2RlHO1wUbMoh1D9aCtqk8IqSJPSWx8Mb+dzGlPO0CN6ymB
IGjkbsnWYTZi1DMpHnM40vImYVEt66zRhx8be+jKRfL63K58gWvw8Cs6xapbPdH/
x5T9fguZr99szl0KhKEQMDh8KcMrtneu7xNgZ+3oUZhsM1soNcrWX+XfQ4ZsrZb+
JfFwh8X8hT4lJ9ODfiYvA+KLvf+c8RloCfv5vMipbtQ2c7nCWle6TtPva/XzRaZ5
VR7tYbWsRPsTG8pIkNQUEzoGpnKIk/jaGH0qa1knPBDcT1wvpmLighaRaktWy+f3
W7qP2CZSlAD2CURMgfL+CW5c3GeZTjID9FLadVwX7p5zs5ANdhsbgtPBnsWAgNpD
rpIQ8lSSS6oPBAUHCaWE53rw+UugEtDR3FU9E9KAqMd75eDAZ9DDsmiLK0nFgY00
6xyC4PHABWOyc3Ig9RoiKyl2hSJnz2pHKRDDo6R0RXb7xU8BcoqbJjWNFqSj1IUl
iUt+mCVh/eNjyl/xDfjAV/H/HvkR6pbFlfIvJPFsg7Y0W3/ugPUR4IpiPMob9d+t
/MI8fi/2mi2Bnsox/Lt9+cSFeZxanbY1FzEliAPg6yAK1KMx0G4gNOdDU4AfltRd
dWL+J1QYzuJXpHca0mubhnrMRnYXFrk25Rrmrl+ety8LL5ofUMY65MrPAgNU4P3/
H7mW/yC1IUUjWkOsiTczpWV+snpSzbHMzmKoK4h/RLoBGmWweEePvRY2T3Xa0SJL
EdQoHped/Y4il9aFTpBALSSjvykqNw7RmtxWk+qz836gQUqftUiCY2LOWSHrvLI5
iK0hhTLQmNfYWg5bV0j+9waVBL06Lk6lLPkN9+Oov2eG5JWJOy1Oa/cb3/Ma83gc
8Pkob2fPwHvzUH6M6oSXelet2p1Z7nWLtJXjTaqSrhKqVbV3R5XTObWEc10eBm74
fKtODpjlamrDUA5SfIM6bofyadaDeSUpapQvlfeQ00j83bXuY1/dHRIueY7p3/Z1
3wk18vGaulcN3BDMEthdZ+K4skyuV205KkeywhqK71QnWRw/2pNZxTTwadrxGQvs
vM1TQgyRK2yrp9iNcIFSi1BVQuNZ0sRTlG/IRDj/jGY5iSDVS0stzL4f3ecdT8IN
0NNd7331sVfEDF6DyxyOugWqUivd32mJDv7L8tEdmMY4vtTdojyyUNLf6lAi2EfX
P3VTN74DobJJjdE6iJC20s9o0YJDJbAFAUdfCFUPeKAuWgr8kBHcXcOlruKzb4vq
saKn4Ni+VDAD1yRPr6mcH4AIoAcxRKK6ezIArcbAzbhEt2zD45xMxzMdtwBMMPi4
dx9pDoRRkJsVuPtGuDFpKhuKM82M8lYpYWCjkcGrGALwODChUP0UkVVsFMNl00Xa
hOyDCv+hf9vxIgcDZmbJFw+kmB8reLzoBcqBZA+qL/UZBxo0yHkOStsuWuftWVvH
LzTbIcn8NjV9G70m/DaevzIMea0+Oqt5H8OhKkZNV1rgDtxb6/EwPL/1q4snyC0i
+QHJDxl1Xai6bI/g7E8DaxmBwzn+HcHtUA48srVUs12LlD99eDgimhFlrY6ZsHMA
0TMd6T2EgFN88SSQEYqfd8c7Yt8eNBYEx9y5B9cue9Bi6q1X6+l62yIVY5MMPXC5
qg/vAROMD7i/YIhtZl0OU/BlsMMxOUCASAEY2Mnqg441pKv0XCCZydPMZuVJMCzU
e563WZVlM76Ze8rSqa8lliOzIUJOXUc7HH4xgdTOMm5At+J18s9JvJxQ218VTgM/
uglV4MegEcsPjFFE6VtVlj22/liT/sOsvmaoAQFDLnZu/r61OCTpsWqdabM/Cu29
w2QWBBhwtbSdnW+5zt2kasvOu44cm7MZwej3imkwlm9uz/GbUOkt5HbL3UWkIfds
Q2Mj7bpezab0Qyh4hVn52/TfsshgrK5Jx29NrE4+zgnS59EJf/lkhxLSQssj3lY1
mYhre4jk2oYBn9I4WX4sBIgWIKJzciSrP9al3tHPr8RL3O2GhWvz+aj+VHHvUJ1C
mRWR9TL6yupSGSe+huTNLrIF7X2UOL45wTrHV3AEfZ0MqzncumJ7aik03i7yxts1
+VuEaJc+Cie/Dv60AFZCAKmiJ/K8pBUJNLMfvNKNda7SBfZfNX0nhDlsEgF2tqK0
FbVtve2iDELTWlS03xeqYw3zgX9nEha701kiEZX+xe5BHyb0Je78qD9fSzSIwoco
rSn97x64SQ/0ozrdhL4VMedOJOflwOL2isIz+YQKAiqHNRPAQ80ef8A2YXm8yJYj
w6BYIFnH5uyqOTm1o1OiFos3Z5IjoKJJ0QWNjQcQCmLpg0FU/y6UW+j//rKvGxTL
6gbFzkjX7xDkg6vYHghYuLoObsma7Z1pWGebFfMC7oGGfsa9YRN3eQZmeP4qAE9l
HvqepsuF+5/y18HZZ3O0SYt6UsRBb2vYfZR39+C/wz3laHxI/0tNhhyavnPFeE08
K4t7AjdocNFoYDarAZGrawj3vtj7ZhxNtwqO8btizvmdge5Gyn7DKS5oXTYwYq6E
MZt9miXbHzCuwbQPfeFLq1tvDM8g4QZjnZ6VLSXfQRuy5fpAFuASplXjyR678gf+
asjK7n+jfJoovwavXgW2ljvtuMfujNuzqo+Sg0eok4G3aPbhsZNyNl15RSufIYt0
GntdgUuto3NJFQkA/Qbpl3+9hUNIY7IiYP34QeWKrUy3nnp0emNio8CNuFWyseNz
tMimzsba5YajYMfePSGuF5FysC7TCyVSrzlPTsBQuMeQI83rByN7Q90+uD4LFHwX
Wl1SUbTbrG0mox30iRlUztUVnyTsssmT3Avgzg48GeZVOzqQkcoKRHf0JCIKeyAG
XupoCBqE68FAdnTjV/6rrlxbGwBqTsf3461GYq6+bsZYI5l+SBSrCknTsY1eWWpu
woWUMhSOtfdprutHg3287WB2JKBkEVUnnsOj9W6rKyt19Hjab/RBtAvrNzmynWKT
g1snrCFus9sfdUXWd+gReCbP3fJNmCZOBmZQyCe2Q6+wV/KYRswL5spUYocTJrF7
uXmbZwc0+UCKmMZ9OBYre57G6OwFKIlF6gG0GdDpLW/vyXShN6+ArhA8ohUrzcz+
Z+n9AobrBMXayxg14aOkJgWVXLdKLda0SyqJrD5nbYZ9Xc4H+HkA6k+K5o1E8nqE
RZvgRq14CFBMslmHQz+yAr4OKKBnyfRIEZptXTt5NRi5Qaq7VoL+sdpgJiPgP18D
Hx3MaDQ14ma4uT6vHbWx32ZxaWCY0eBZl/8U7Mv+dF2r0SjM6b+WSam1aryf+iU1
G5z/oKneF5sAnG+/P+E0gsEqGzcTzZZUoogXBJ6HWwA2hfLvidCx6c0hFlc0dpxr
6AyexjCIvyveM2Va+0PlvXddMMRP8FQBfOhe90dJZe6mIMIUp+UK2CTKUXVcx+Ws
ILTm4+6/FLDEIqr8Yx++w4nJSNEeGHdI67d7rvxvDCTj9qr/hixyIQ9SN5bv5yDp
QyKHOmv8us7MEGA6L0GsVIrMfCcyKFomTEvK9QHrSwe/V3zaQjgkEDvBqX9LnrG6
Zc37VRfbF6htSowe4jU4DbZ2WjzzdaSpObd+/c4sZFI8LO7jiue/T9+gw7D0qKud
e90QJA9RQiF2v51KrEPgC4h8hnSIbqECYb0CgwWFnxe4VMg63fCV6sbH6wwTnoZ6
AY1I58WUYHC/F31d06N7fzFESxCgm26QH4pxtJxEP8F/NWla6mqodKK6OjOyAuQL
hRMw3RpcTmjJmmgSsuJB8Mu94o3KtILjhyKYOsi8tQs/j0hXaLcpZ5AZv3+T6yTm
mES7rJ3iuHL2Izd5155LHGEZ4J4ml62yHT1Iaa9WNv7GSA88FGoh0sQzSM/qYehd
jR7w3eAIacw+y7UfQKOHix3VTrT//xHP8AvdlGFpxjWC8LotF6S6GUdYxtxKhnQM
cRtoJi68PhmXzT7xxtE8edbXjJ104HI8Ip6VFtcLMhbfHkMCH+fU+kLCUnjH6UbE
1QLc77Rq53Px+fLMhKSMawLy2R5CVLJl7OnESzhr2xqaNJNzzXTcPHWODbTYPN6M
wJy7M6Rz4YmWfG0GC368tl8hMS2eKl4uGdWnI406S+h7VvDsVdiCUe6/gUk0cVS/
NLUmDywwgD+Avaw7bItYVaQhkYqbiTiKCWNX0qSKFiWraISwo755AJyc7d/28xY7
pPEDWyUfWc8dwF9ca4875bsJ4U5BV8xS/Pl7H2NkRIfY49+ITUfRp3UT5jIjsgHm
0vkNPKViMVvMQckLkliygPR5YC+IfrKDNfpgDnhOZfxcPCr7RWT+XYRgLgXQrtbV
vxHajQXhIlF7hLIUg/+0KjDf2ZVHgVzGawIFOZlhj90zA5DEOLAp2pVBOyTbkN0Y
DnvrPgLbIdw/Lsed7LARW2bqijvH3h3i3zHgaSRfktEeBpdNoOoY6eOy3wOWBkiV
EZG3NlOwWr7pa/CQNHTXqsH+YixBNYeZa4CjCJxNo4Ny2xwWxQTaDuEp0w7WLPdO
JFH97cy1VvfZCSmrKv40SFTTyYNtlUghOBfFueRP7P/b0wAKso+TkqV7djauZTaW
Dm+dEOxGx2EVwhTIl7bo5iyD5vKsYLuS3rKnFts0TIURaen8UHuBj5mtWe4Nzmnl
xo7JQ1YB3pu4F4wgRVYD1KY1NQ5sM6nViirkKmMN1dEVu4HQZiH22ushNaiJQltN
Vhj4Jp/3t/q2O57TkBp1DbM0d3EmDslwfhUElC4ruDQbWfSs0KbGcSVgdfsBCsFx
m/Vw3tgN5aNVC5W0aLsmaAWLk7igjPM1KvClsDso4D3bYwwtsQ6vyvQ+irzrgf30
Dk3q5oc0/HgTTsy3xnLcgJzD/xnz/G65NDAnmHhfvW9+k0tmTEeKtBDmXI5Nox2m
wcqkinMCM0F1ORaPGhYGbjZ8GtYDJLUy9hgQ9oN9uerejGuPvoykSPjNhpvZG/C9
Y2DVPut/OudHhh3hTY8DejWjdrZ0YeyQqQCrJZA2qIEFB5Crwbo/ZpX6Dfd5kc9e
74ATOtzKWZsgk+0vaFYB8oxdnumG1j8RiY2UOpKxmMau8+5ixvcBr652zg4957vI
AeDiIuFVzj/CNIKH4X6B9fdHDzT5mqqVlQYTXkF7ppU+gwptkHe0kFI/yvOY4kZ8
wldwrFJzsXsg+reoIsEv2bgqba52Uja794V71wXRQasv+HAv9JR6K6uVDf10VCWw
i9yno7F8tWG0cq8NJWEp5cnxrU99ZMl2VZTGIGicgJYbu9zjhxLi2ev+1zftFl3P
bHeDJhYa3AdxXpJYwP7LnOLukPFFcCMRgRYudSrO1PXLsMkMPdfpV3/PLjbgPVyZ
Od8HfW3knZpTMXblJDRlaZeRXv9/avuH7m2vvbIz+y7QekfA+P7wFC2hWZ719iPg
sRWLB4LMnTNNtqIs27A0iOd2YNewD6+EyCiJu8qSxRb0hu/IiMEUMPmNq1s1hNOA
NgdKkJ+O42vgbtBHHhFZ7Q42/A/rA30ioXIZlawp6NUw3FPoH2UCZim8MQDNoPIq
QhQpZgrS1GD5RiNKH+Nk4POnGErVCkiQ/vEPGpF53ioGR8ITgl2hvSgE3CnIFQ5p
6e4bpTWNe/OCnOYLDWJYW772HcOgs8Miy957rS8CFlG1qE0AiLqcRg72m+4RUwNK
XWZIsqBWBK/Orb6mA3ZNH8US9qYbpizkZGTh9MlS4zsiaUl4rkzU0GfhKN62+r/N
CrK7bBPSleWybJ/z3uhrht5O7zvF4w9K+I72blaMhDYOvY5KJH3urwQysgrxEDfV
5MPWlUMrxAV6BFJeSshxUWfsuEQd5lcHlUAedO0L72ykrHH1QK4BF3bhbksrRuZ2
NVhMe6HjGSK7chInxhvs5oAdJ5ZvJ65MacUWHqIJK3w50wqaQ2MOIcU+C7UZWbFm
ccZ68NEZmIovf0BuvJ4x8OePCXyUv1PFJuC8R6zrROe4gf+lcxTHhk5v4wn7wfZV
1/HGWNEph+K7zbSpeM9pz1tjBoRTUKNoDf/RExYdek8dCP5NvO6LAerUyORViEe1
1P/8oclEDal609wfUB6mup5FVdIzLtiZT4nR3twyRbpxx5KWMQg08LFlr6mxBppa
1FcUCw4xQRRq/zIw26TCGvzHqLlslNcOnaCe/ST2d/QdAigDbot0xMa1AxWZo1Zf
taTc/FTyvWSescae4ZEee2pkv5TWHSOqa24LggjNfsmLrH49A/CDXJCwty6KKbmy
KvoN6P93mUPGPOgB0QOPqYk7dzCRcM/78WmpvoVOMo8/wg5jjZSxMxONcDMlp/PD
LMuOQ3RX4fhdW5xN+touwVV/SP+ddq3C2NphY5W/XY9Ql9ypDLhBte1E+hm1WEye
x13ptc41LQ5LwTDfzyESGrpGgAQzNOGhB43sEvjl5Q2iJEVyVH2j5XpEQFFVmW8i
4+CzJm1WooIM4vYd+LIrSWg5zz+0VsyV3XQNSfBR92F3RSfsYSUZ8fcW09hCz8FQ
rJO9TGwKIvWy9eJ2n5iMEM5qYMPeOxq2fQhA5rpoBviNkh4Tzcybnv1/P8a6nB5h
oyFWzMwLJ3CGvglHL/kHzt/76RCekOxx89zi0gKvwKupTScYXsZgp5ZXivb1t2Vr
UfF2nnR4TJl56SBeRzzJvweBmkbVE5To3D0EPJ8aYeLYgxb/8EVmR6Kf0WoST8UY
yK+rSb/xtfckQkwJstNJuNBg3uJuY/HUhwXwnZsOGkNunWktz0bQRLIgHT04a1/H
d63Kh0bHYldASrFo/voOqvTo+G4zHv0b0u+k654SQ/2lFkt4ryEpK7N/IysCQMAI
lHLLiH2NNbO0ySYVP74UZ6e/ZUnpUXeQsbMNMA9JegUQj+NYOxJB/7tIA+awIX7b
j9W90NiDm2E+21m1mXp9bPKjGFDuqGUxu3jnN6DkvpzETE50YUg/NYeyXCAFgxlN
iaJMf7zzu5iGxqYootmQzb5AutWV8PVyTZU+3AeyauxRJydjhk6SCVMKLwq42pER
t9iCApS3LvC2KF6tRxLdBz1fPzJxrSC+QOxOYCez6V7zAus10pXfEI07Om0eE0Hl
XDRsZewLl//SbksLBiAYiifLMHAABnQYPSANBUp5grJqJb/emBshMkd65oY/ENNU
W2Xp0uCBHYJfptQqhXZvIN9aZXxSVzwXYLXAn+b2umy6h5w97NL1+1NxSUi3d7jz
ZJ0T8GhBy1yYIkqGrXSyvjEvlhsx+0UqDTPnis269V1T9ceFVpZzIfUr86kVI7uA
MaUyCniSnVEQgTY5kZFgNhCzfaYqZITfEh8MTpZyT88mtRmEyOdJ9V4m9M/9pUKu
dVhXJtVWudJZquzRfWKG+1/qIoX2qqL9s1TQNwY099YDvj0UfdACucheudnTqWzw
nGt57dJR5z2kPinDhSCyCZZSY9Z03qQSd4g9NfFfE9UAUjn8JWgaDaXyZWSbyZgW
saVPd+FcptNUf8SRyFSjNXt7SkaV8TCkvJIp9PqkfWjS+RncfUKUbPzHPDjLbjo1
r7dzsbAu4HgDPp8UU/RYeXZpiILjIx1X2d8H5UyCrBQ8Vha10viIYkf35rfmVSxs
hd7eG25VJi+VI+tZqew2FFhf2jI3mv2Pr3fiYSC4Bwrlqhl/MqRxTGU4VsOmCXTd
QmwWi1S+31wLWC+OB53nj3q3L58/lQqsGzUVRCLNEOxozoI9EL/BijVaTzr2nruD
+4r+Zqhxm6TTseki7BzQe5FukaJYLLNMhGtX5qKQXGk7nkWxuBPiS1JwEe6uy302
AZfpBfw9QIOvor4GN+37GC75enaJytrAebz7/tZcdm7iZJHbTJGznsWht4JeyxV8
CJPfdEir3S705ZNpiwWo6NbJ1jeo63OxgFeQRPQNkyPNZx67HbxxRQamGn5um2sx
4eJ7rrWnsQ5eXihmTQaa3M7ZvhjNC+9m6nv+v1O1bq7hPh1Rg5MUDp4f/zJzDoBI
DhGmnL4Q9x1QoA1zd3/DEUfKx3WHzA7ZquA0qh3FpncUdNC5qLutjylaEbdyx4hz
s/hTGEcURJT0EQ9Qa7b8rMVgTv4S9kzRNx9Mc598dDffC8JYQBtMNy55Y0vqW+Pn
q7HeU1Hur/cMWPk3A2a4DPyEF9gGTQkanvTsJdHobuodGFRDfo27totvu3Eh/u/U
cA1W78c3x5s+j42kHqjWJLOUZZ2eNZfu5REv8rH8UwwQIUDonk7LFJJ9E60uova/
QYDsZ1NfuGnRXeO7pcMzfj3Bj4BfU3pHKs83irPGq8A7H4GMLaYIE8dTU4hndtk1
XTUCSK9ebw/sJ8wlg/IphCii50eXP8YdxhCVMRz8mddWvwfIhQK8w0PHL9Z2KVkv
0grdBDo1owdNoiQykAYss1AOXywgX4OA83ohO5xzFwFSBrmQatMFp0Upc4RXhrTg
yzSQWEBj9qtg4/km9u/YYr4OB2LgQsj9QUBkuAPkMqY3buMDKG6wL0wUgyihTZeW
Z+tN53wiUIheF4YvxDLJiMvjL2SZ6mj7Sl+voo5WteZQv7ARre2StEgxwZ+vYf5r
uWSeXS+exruwZorofc9vJ5wJx++qyDcX6Y+epJmncLFdeZ870ad/4ZAmTLm/ntq9
3ceg4+TDKhkASifXVRm7B3D+FxAQB6EqA7prmFq8WDf+ZjHZI2FYRtFL68/MJ7rV
3OU9jLRX7eHI/35GaUDWLoLrlxYomwWJVpjh0oCN8DaeN4TAHgrmBl5Xhu42QxvZ
3sK1C5c/58hpnrv4ZBvYBdjhFGVU8XLiVSllFBCxjAS6YBnqrrmRtvlm7mbYbkXN
mhSLjPVfKq3LhzM8scqGUTrvbbj60VuNIs5E/oiqf31+GGhsrAS+8EbOpo6YbUC9
wKB9t9KnBe95jnVUUrHw6f1G2iI8jmgUH/y3uGO0vwPJHKq47DwgPCDm4vjG6Ivo
im2PdeDaEz84ioSGN2c9mL+a7R+Ksa4/fK0/XoZtEJX+DVj+3d4JEMzUNh38ycn4
cLbDErwdjTB0b4K6//PSb7pPrLCZKfn7qaXikLKEqPz7tUbia9Nn8N2pgskeDmlr
NunpatwO3jmZh7xELMxuPwmJJ1Re2SpQ1ahvcnM7ta+QsTVK6bD86aODKtAZosjs
wxH2f3komeXBQj4Skox9ro60Tw4qRNySSKHDrLqOrIfIv+DGt3QVNHDNBKRtotLI
PKen1z1wZ+xs6cHN0p6MgPI9S1/HetkQG4+qkyBAIfHgXAGNqNiFAbSbeDLZuBGG
4mXyK/V0CWRt/K6DH2d7lBljIjtwWII0k9PGy61GtsdXhd7hratI0rttr4QlaQgP
xasxU91PXRuB6aC7NnzJTklrvdOiyHQcmOfCRJzZz2KLGRlG9mpgQPYnUCDlvLKs
qW5HJGiPFhefea8w8S0zGdi7xnPnLYSme6n4cs+ZQ1vzEdZCfZSUjNBaEYsa2tL2
VnKr3pEYRIb3NTDvrd6rp4LnZwm7sBnyamgvvre6A8GOICNv7LyqqNALOTc+ncEd
q/ImbruPdXqDxNU7K9krgveHDFHZk3l24F6NDoZ0ppYOd5BMkqxcPo9XYh7NcGw/
4NDkwhpCkn3ZplJrILGRLAayD8rCA+Q/4uqro895PI5eJISfW8E/5PWvC9O6WnAN
jm007dObH5ckxt0mIvX/OX4nxd/3AvzI7YPe38op1cVlLtI4bNMEWjrY6mviLZoo
muAu8u0k3ENAAdg2yxd3fVCNsePF6b0xyPwvKJGblEX+i4e6trHIXjeV3yenzAxF
K9x2r2+zYAgJIomvONT0Ft9S5exP5f4IS5HZ67UwpMyZbqWTzi0qjnRpZldk395F
DnJLIRF0C0L+oIuM5u0iD1tzDAmKqhj68gDADLLHskmdA2KtR8JZNIFTfuySZspZ
PL3+BringSEnPsp9QGNwND8gDcE4xvjEXSyFj5MTwBA5qMiJQOZ41zn2tAQtYyIT
tJJ/0ZfO5/p+5RJXKx1UYnDTaHZGRo08MZw5P57vxtgwLOiRCYFcg5IDuE+Kvl47
YWjhKP/A9A5BqbtX7RL2U2uQDfjgFBeSFtxW7yrlIm9pnByFbEDysYG+NutGMz8D
s9tV21L1qg58j+c94Jw3Wywrt+GvIRzg/SPU8a3qGZt23CYCDuXJ6WDzX4OIqnnT
ro5l19Y4MQqaU4YRaXsevYA4Rco2Ot3lGgm/6tDH30MAV0EjvwJ998QdFlBrO8fh
6Jv+d4FvNS/s7K1q5UKI7GW5FWgMc0I7Mu6ji/6ANUqFDEU3GQqO8Ine/TZTrens
RLUDQ0V+zLxlNwwUICpR2we0g1yeOXBsQaYvLURAlgw9XUr/kQu2QvEVPym13TMO
PYxySa3BfCEMo+HBP4CC1wWndNOrCOagK0LZXQZVAv5gZZcUl1+cRWdePszpHBv1
pCGunautmNHEZ/lDxolSDRgFnJQsPNxJHaQUrXaZJh7Du0H71jlqa4Rh9bbdW0gc
YTTvuqj6SaHJ5HEDPAhQpzcKlvO/NS+ka2tpEcAKp3egZ//f3JOHtbOGcDdIjyjH
d4xCVDoOlDzhGWuPYlZ4MKwvqEtNaiML3VHdLD2WFSt+yAUJSfoMr9x1p9qmG0lj
kwXzWoc5JYXrfITfPCffLJHLkHBO4N2aBpGYd67SH0jMitzEr4md/kxdMRnALPZj
Mqut5373mhNvSkxlkwklESjbuaLzkR5LDBf/g3e0dWWoX3Dd8T1nnNguFgdyqTcP
CSvzNMe9N6R3+JYG5STS8mK63TfA/QzGWjEDYyItInc3pENEdm1DJVfQlaq2hBGe
rDdp+sox1FWyz9jxI7JShDyhOlqs9QoVEqLt+syhU7LbfccV/6G9WYA8Wzpg2uKM
wJ/87UO5oR3mMX74NWoO6mp7ceXBbcpo/VGds3wIAgYj3Ud+kBDm/OXki8DDjW/K
RCsptnugUuRI1XsdO2o3o9lH7VcGACLRpjZj/A8th5Lv9kGXTw1VNsGFfGrbjSFe
9QSanQXzTvr9C/McbqHEKAqOJucXCqS2R8KFPhmTgcEqPq2lH/moNNIR1t6Dj10X
7IJV1zv9sU+MAzwGqRMeL2Hhnhf2Z3YTe7dYTpj5dj7sj2vLXGhyjq8p3p9eLWQk
g2yCnzkjISbIqGhReXXZOETxlhtTP6f8ycHqUwkop08JBEm6Z9eqVuVwQnwSvlMe
I1W6XEGicm2IcRy0Op3shBk5ttpmzxCeKQBoojh9H8UWrdDcJgpEEdyAxeAG03Wa
sVDSrbiURKeXTLsottxB8AthMeYKbAO1MRew+tbogA/fY+IaBI1J6uF9mPIVufcb
r71Danj2kjHFpbV86cTgF511Wj6fU08Q/DFHQQQtTEVUbkhjcPC+BYRwIHEia/5A
A2gdlSw5L8oNt3PgrA9ote8YodtpEjmy1ObUI9VSpL4pdLELSstfeJLrtmpDg/oW
PTngS7NbYGtjdTknahbUnrv9W/N1js3glJ8l4wOEH9LZAleW4e9G92XJZd0En1Wz
yieNNg4xSDQpdciZE7Y2O8Z8VFw2rfvfI/xuqg9F19+7jS/aN5ISJEm4eqUfY+gi
BesATdGMbiaC4+OjAbPYYP1hamRYnj4zUe7/PAl/c8dTDLcyi7dYioC1Mdx++0C+
QG5+XZLM0uoo3lsQ5A/eNX0xl/ztq8+0KgBHfzimBhXCmhsgX8ayvz7qpvMlIz4I
1nhIEWikjaA//x04ohzod3C++COwzY5J8twcqoFZpu1LjN3JuvhtyvHZSoBBb1nU
EOFLI9N/zh6NR4bFV6lydhpWq5VKAlNCKdxgi/hkuWUgwatDMS0ayNl/3CyEoRZo
n7C2fwGRK47F36Zxlef7IyFHErCGv9wQF438QZFFuM8VK9dmCoKxU2A3dx7dEHMf
7087Bc5YYwr5/vzS95WT29LbJqgQv+3nFOnboNmnu3WWgNjqdx/TdUZlrSdFM5do
+EJwiFTXGw+aww6iLKDNe3xKoofBTg16xDErMzgLTj4CE12nv4gWB1d6MD2dH0RO
GsQrgDWG46eWEaNTlsodK8O02vkeGToWTU+b9kBCHgH9wX/c3SdZl+km+Agwfgj1
3Xp+owop+7EiAjr0uciDCmSeRzw54tFfXujrSiFhgccHZ0Qpgp5EezzmtNYJQTZq
839RJzXWearvDQs6INKuWxu+beSxZya42cCdq73e0+HqVH6GSuAN7xR8/FrXFtdy
XswpMQZc97LpRJQPlIF4vnLFq9F9Cy+d5ztiOeQoVbgI/XvBR3sMH4KCNizq5/rn
wYTOsRPgnLCwl3XdqaQFqGs5SwJpWSkpn3wtE/WM6w4ZXHLiAow8bQNl7ILGq3dW
XOcrkPlRU6S9COmWwwZXJ3lEgNicuOLoJTSc5eGImo/1vkrmaU9is4Lv6lS5rzbf
iMelRRRsJCaPwpDt1Q56rQkeKOut9wIxacQ5Q77lb/goxCQCcPyeYUxiEgvWUk0u
m0NmrJ8D2BzpGJcmd1GtNHgaYBtrPS08E+GHpxLaQh0oWI1buh7w7rb6PpwFdkiO
xTOVD/8uKWKL/zsxlBY7RlvpXChQpwmXKn9SAE2qgIP8JKyCLN8LKcxwDmJK8ijP
Kq5PyWyGZJaCaGvA+bJGsdb/HHnC3uHVIZ+NDTa3Y8O4XhtDsHvtsBy5SF4CtqGp
yWPURebUJEPhkxaTRcWQ9A9G/k7DF76uSnCaTpb0ujUJ6Wl3yaKKD2RB80d8ZIF/
YGewQXTrWnu7OKbrneJ5QqDsAvTY2hHH5MZq3hznbxLiRBpAGF2qP/wJORWCJSqL
DRjVmjZFxOaWEuL5fHIXhcBTeTXmykHEGVIYVqS7EtwsTE8ofPfH8z+tBkfLqroj
PjRnVgKfUjdNpi9KTyOuOTb0yo7onTMozhXfkep++rafZMSP93ZPxzUAiwx0dii6
Qewi/hyiIiDeppHumAMFfcKLy0OAgEUVpeF+lYswYrs5v+Bh3MaEw9CRVSpmUEoh
PksVKebm5soyXUbVOgqV6AjPYxAectSKoyTMI56zrowwvVEjMDhq8nYFjctQrtwm
+1e+wVhPpbnLL2Y9gb9LKENPe/LqnCy4a7cxGzu0kqakzJDDywaoiy6DVBQJJ1EF
vuLoG3thlW1FOMs/sSr51af3hcCS3HO0TivoEpT6kcJmATnGKhu8ap4Tq7vuHPN5
RLkSjuMrntlyqA3J97d0pf//AZLxaPhYRPWsMWjLtjLHkC8dx4hCaFJYHYdbSDXQ
vDuhBzI5PjQR0yk3uOR9TihiptCGLAXFLSM2dtspJBBVOSOTi1n/mcF4G+MlRyp/
MNbW6dDZDM3NfPNyvj08O+x/PZzMx/S2EGAXvomV0ZhG53SGvIT96m1QgUXZm9nv
BDeRlnvX5BeOsm2DsdEcS0rbMoekiyxttZGMzAcOZKCE3lWcvZ3ei0k3T5WNjHYy
m+4tsi2k8IRHyl6//0STGoNjQsBmGPDgVq7Ll/rZ0UnaEn/rFJ7pKBzik7vOOWDC
iuVNhBuZ+upjLHO1mN6alEIm0NaKr9dkP67X4/QMH2URYchFVQ1hWiDTpCFn3P0g
TRQDvir+rNRwttkJFFwnkM2dqtyT6P6GGCWiOKr0stjp2saFaFUMbcGEAACBBaj6
sICIDCFjznFR4t7tAp6AKWYOoWyPOoj3hWMkil5XDQazRr1OFDPNCVsDd6ZEfB5L
J4zw0rEaWs3XRqLrlfgJQjUItj64GmjV2/i2q2WxAE1cnUhLkkqk5SWmHmecKNBA
aZ8KFb7eih8bPG5zvyIUb78EzhS1x7tPaIZFZpUeKtty2zUAKBnD0Lnsw5DDPojz
cpNR0Ct/3Uk79y+9nuWkIu0Yx8Ui+PAS2d5uy7PGu9RSOC+ljrqETEtGbAY47qb2
QOMIayUa1ljPCOkjm2xXRjjAdpCa03kkO+YhmB8Dm/X34r323+2g9cr+zEW5ixpS
h4c50r6b5MYISZdSwtPL2OlQATCEMIXEmU+RAXx1NCHneag9P4qrvKQWbxNMIh5A
2daShvU1bCtvThbYwO/LK4agr8HazhfxD03aK0krPZs1t6XZOaCNmF9t9LD5FpaU
VrWxGuEmeTJv7jfroqx98+J5mO0uIngLmX/FpIohvieHlyV0pDQTz3HksrSOVruY
wfCibtevzwmZmPwN0dj0z+o8Mj76crWmOMOmcamsrFfREpAjyCye04V5+sQz08TG
ftvmhFYEGQ8VX7KzEJgzOcWkRbKFn92ab3p+y77ov+/zyFDQcocWLCGEwm9VBv9s
vTBiqh/ZMszmt3kovCLvjoRHfRZffLV3U14KspggiiE1AbGjKk2ZSukcVsX4INL9
SXKtTFyFU3X92tTfakS4HLnYWjWHXLp/Gqe73JChFQh1PqT8Fv81liW1I9CVSAgl
rSpCU+5HL2cyjwyIxATTj9G4GKbx6n5d71sAPo+11nr5EcUNy2AJLtnZnY+CLAAY
vEDEgkxw3DXsic0DY2asGFkXIUrPCTl4eodSK4E2DHdZPa9H+nSCF1gz4F6Kaa01
rqhCG9ITS5iEAr40149Si3/nfxD+nxBXuIhLc+LbNBq6T+q6E6Wcd/6u5lk9xf9O
6szc/FuFw9f2T6ZGOVQwu7sutjxCe/jFOTZZY4+eWHJT2SCAS5vaTbsuwvpLNgBA
V+BPFMzLIqpSOXUX6Tu5HxNIPPnIUiHPP4kl6z8L+BnXlrNgnmIoTA8v63SYFCFA
15h9fMV2JdbkFg+twZGe5xM+52SCkPjYzKEERwuZzUTMKuhbxmXHKMF3Xf2eLlsQ
h4sVv6iSXPFa8dA9X90FVuW8qwYwfk8AhxSp2j8iilLXe2C04Wo5QVHWBYPk/BV8
7Y3lL+ABkls9+jRYGFTYN/C7XuTy7hEz1S0QNHnVarpWt9w/oXdI2Qq0CnvijmcR
90QcRlGRzWaVZzQi5rT5Ek9NK+MWAQc99ImJ7tO87CoQyX4EcgkCA2vDF8Wz0a1v
qz1Ep77q0ZL5bqK+Cd2PiEsN4KGhiOPkNEPZ5L3a24raj3XK2V6vQQo13BVKGMgO
slBHHn2d3D3rCOpVCkEn0Syw/UvT1gRHA0DWOtJZ8cOd+qgPTUE+KRNsO9D4AdqB
L/ZZp6j9WxYi1Tp1lsTCo4OxSlkXkq4Qt3VAT9QsZ1YAWChZMJWrXfwtzEWcAUtI
uXMYr6kdBarOOxuPyhj2g/UDhBtbtHAfemeNbH13KVQh7KJRj2v25p5c36TWewCL
VXQ9F0ei8gVHW+EH7BZdkWCDCS1oF9wIXhSFTcJzyYeswkAW/h39KpF/WKnGew9T
EYlmWsbUguYMskP35wvIsAqeKMrlswoe5hra0czkN3oWkPIQWXY+cGbiz2r0doHP
NsL1uCoxqWWRiUgHpjAICOvcXFMKNqEDxM22WCpLgsJD4t+R8hm8yHvsRJtNkx+8
fUNfNEVOVS8/lPoSWb6nTbOVFpCAfQYyYKXFIg4KlQleixexYYENScASxZJgTLhs
8YSn+39gspIdnrFrc8MV+Eh0FsNDx/xFGLVMNZHY81abngW5V1Je5ttggHpcnZzY
RTfP52aqiYnfHzbI59Cv6ZN57V7PHpw5rFJNuJ9runJbvqnT2a+dv/9DFpL40b8C
citX7bowlQ6+od5bIGm13pI1z29zlAinbacIwFzNVLxz+2TTlPQj97xyE/c4ApTb
Z1kZ1ZGKtw5igl2zSmiNIFlGkOnwKNdxb1WP28xkmEC9STuxk4C83tc/hniXC8eW
fIGq3Yb1yhHk4YPkOjpJx+4C3T34+I7VKcB2Vck25UDX9c5WnSceL5xQ6wTsykTk
0oGj9f/FrHq9ekk4J2z+XT71ahmcqZ2cqGXPYovq7SSpOecZsuR4DO4ykfe7QLiE
VeQ7AgFFJx32tGSG4SU76DHXa7OfHJWy8hIHGxepaiwq5KkbDIQAsfBu4e/S2I2v
YC/IDVedxle5Sq9AaND8xMyEXOrvIBIYNYg5EMYshURKswTWqHlEEcwYQCmCM6LA
RVX7al8JvuwqQvnHeCABhFoSS1gMmCTBEPGlrVPkt7F5XNGyoA6keoG+PInaceit
2TXPMzDILjen7PyguCHGl680yRs0E750ODeCWadQ2taZojqNS5si63zGQzAzjvJ7
84oM1AgzHkyiVIHVr8mN20KeeNjorTlSPMPoB4mbZmVI+pabg7tzYIfWdNBRIKcU
X7ZaDrxd6zpOJ1y2821KzqfgSsRB0Lb6okYvG+0zosJOHFx20E9IfEPJuo3Orypx
jgMvdWkGElbTjMt71KL0dqeKztFoAdQt3qEMcshsHwspFAZwcw1xGJF60135e4Et
0TXYypVy5gI3QFcFmm8mWm9mvGGJerVhwmxk8BcydSZIqhcKsJrfUZ+Njk64qiqd
UoeLHr38kFrvGk+Z3aaPHuE98U/X7lczXXx7+BVMUnL91Y1DdnNWkpkrs/G1NSD5
Wwq734aysLhkke78hp1rwmLh71Yvs8iahsjdEjqPieNhBTdRDf5TB/gt0UrcTh74
a+qUebBgg32+45qE7TVJXoFSbqs3YsOh3XDtIuB0c7SzqUMRV48Fg5ViDQ7vtxO3
Pm555Y4cVE43QhvivK5AjaV3bcYzMJnj7+BP1vziioNyYxZQ0hcfChLQ2Vv34HJN
E+rW4N2KdUanX659HhYctk+ApOpMR9TQ1SRaEtfSpTb7vGYkUpJymmb42M7vces6
4z3LeOT2hxJnb1XiTeiAN+v1+PZYkXz4gIgdOpBXMrkutJk2W+ehMll+flHsWYCQ
/FdVwVM3a8mQV6HrJ7NWfE2lyDDd8eqSvAaH/vcewzfYwbzsd7CJQX5/n6Emug19
K9hssQseQtAPFBb99qS5ZtWiyPAVXhQmKYMu46g1en7w4uC5rfi9paqoqgOn/XTL
6mrh+eAtAyaX/Tqdgcb3Qn2nDWuLAX9EOUu7qRy2LoRBOuA4FhyJ+rbn25hytglK
6g5CZUdBH6Umd93NSJunwDOiOppcLIeWpBuhiQ+gmuTOBPndWdPaA8O+CWZljgma
qHKQnfj/fJAAFwaj+qGsuMlZD8BmTnqUYcrMKC6Z9UvHej+qV2WzQQPDxT7jS8/V
ypgH49MSbBGCl9bCbja+vlsGUwwGfY7cdN6i1Tw/QJ+qZGeiaBqQ/HIqLDqZnAcf
gpqWMuvH4mJ7U1xh0Nw9+M3lwMq3dxS0bB9+C+qfk/hiyp+wT2CEXkUDlMBrydDb
UvNCDeQ9LS5fZ80abvYPW92m0alu5h3SIJ5TvCyLNK+1gooH+wZWUMZIIoA5vI/T
DYP5dnSl5Ja+h74YibpTUIEN8b7g5Yt7h9FWI/YSf713Pp8hoEA/zJ42L2kXNzO1
VXsfj5ler+3D6lub7VkvQVr68JGW6I1u9MWueE1ETC9CV6CC1BrnzN14ih3Rt1QN
vyPObxE+k19/PkX61UNs6pU6rKi5xGeUXAqfB6wxcQosKnTycib+BJLU1Ts6SAbA
b5X76jYEHHGVtNSOfkqNzp2enLnr5ScVZt4645gS112YxCtHshOdNGDaBSiH5y4W
dCUN0oGN+olAaxcKG66mVGKBWw5oWxNA9KXRxe1UeCpg1Mmv5VLsconQsC4l7fvz
JP/HdJeKWF6tns6AuYkEeomBGkfwdfjTjJpMHIMXJ27MAFQDnvbjsmrxP7ZEeDSR
LCvuwYSk0mMQu2I8ZL3Ck8SEInR1bWkXfJVLtfAnglX7mT1ts0iYH3blnx85Sgq7
T0Pe2vkssmv8aqDwI8LYeY3tGdwtOhldTf/FChZaYREAS2Dyq7y3k4CFSbZGpV3s
JVrnCeTLRYH833mb62xOMHc4SqEj/8hN9mrEPoDf0PP/nJMxlZ1bNUCP6/VrIaNE
1PjJcL27/ZuaTVQS94cJQ7eRrqKM18GM18im8NT0FClti9XtCrA/EBsz/FHSXkXw
U1urM2dLx33VTvNJnrCgGwPXviKvA2whPZT7UskVnBSvVwMBODxe2ogxOjCVXLPV
/oVYkx1DW8tjmZKVAr0otdsSLl/sUTyfblmh7qSGrFPIWqwcZ9KQrJStAYGQlbCP
XDDcFXKSiI2pu9+1/baDAOObPy8C7uNhR73LpAk6lWrUETowYN9asWYP+NzQnjrw
oc7j91bTC+aQVlfTx2Ix+tkckUnmCZGRUZlI35sgfyFIDUcKlnltafXxU6+VqDbC
bI+8hIIR7Tkd4CUByK2wYV5YZm8qHnjKkl/pDgHjr3bzBCTYJ7280pXT9iAwrrjy
6wjUMXSN1SNsTMsp4iI9CkIEZRRvrALPCDGv8l3uKq0HcIfi2Qsu07gb8zjRyE5v
8vj70YE/t8zXqFH8YSFeoJV9BxXOAudtZii7BhLpMKTp/166ke/ZeHMt4JD4TKBw
b5HekBYKaWpfD0Y1A/ZUe1Giscxg8Y02YrcKZs+IAgpyWQwMuNxogaqgFOrpTdLS
9jsu6jUYJ3RtQ31798tQC4+kJIlCCTtDBsJYbkz5dR9nirvXGeFewl+DIzSt5bu5
p8SV7iqjgdFJtZ/gaF/Yu7DCeLUL7bCDEg6XnMnDV9zC3I/grP0NONLsPbKpIYrW
yOCeftcevZVUjQpT5qyvn26RIxqHaHRLqZnno61/bNmyU44zqyxmSZMKYyE6uxQX
zQBjjxlAjnkjt8AetGupcuOMTanDixW+URyRq4VKQIFC1RbdsuUcbPDlOAyFLwBQ
ViuoaROnrKIc0reYiq/DULJePXlS8ohFcXgVBr8tz41F1/khJ1c1q+YabxyAisS1
GZVby4qDkGWW+5A9cMh7bve7H4YjrCK2oCnG+X3IZeuEiSoVYzATG20eWzXQ3eH0
WOIqIlNKqAucDjUY+ao6wYPeMOb1zbT/cpIxST48SOVu+s4XjFVBM4REjCgb7kdg
teYt9ozLZ9aMG8CsIp6cfLHTcd2O5HOzWE/PSmlFocZ6mCkmUbkYOa0a7oif5db1
cqX6hlb41AIO5e8PRfzIoHtK7DaN2ZaOxEZLaHhRkP8GrMvi/D7cu0P9VBmuK+xX
xajKEaoQZFxFY8anduLxilJ5wNYAiF9HDl4jKSV34dZ5og7R2wfGkryVCgn/VZTc
6rZgx3PK8YLvGxfFGbw61gVtgfpaa81xdJtneB5mRpxf5avCxA+Ppb3JeWCoeSFp
bNKEHsfWU/OLxvda9sd9sEB+oO84dii/Vswb8n8lGSp8SW0C+aeIrNp+9DNxqgiK
pfwHWpnpUHY7vyWfESEBxo2rgHOmMRVLMIND4u6VTYSRXtA4ti7j34SZlao+YDOa
J11ae5WvGrxPKxHvh8Ny3Wc7II9hwKv5Z3cpUGke8pjB0owb5ce6mVNxWjhF8DIg
dDFCcgvaddCXqdIFs/nOxRUWYeNhwPqZf5CsKbwVg4DnxQmGsScKzUqZjNWMckTb
DU7l/iom8p0zpIpU/qgNJ5SExv1ZWb6/UXabN1TIq2Jd93TbLMXwbPKKRdAcPKCG
/KYYNY8vlNjh+pHlHFuN61eofN9CWp+tPz7Jq+uQUMPA2dAZp8ec44a28RF7zATE
03jhl0p2fhCugjYXCcsYsAQfoF5IbooCKw1OyY/46NdTvA67PsR7wFQz99RxXq2B
WxRw5T8lGDSnlNanJqbFILE2H3D1lnRH3gGKPWUWR10h7ZEJvA/U8q2P1CGpsRdt
DsIDaRpkqI8/Oz2paS+oKWUO3V41o5hII5PBuYsdyl1xyyLLp7UJLa50AIhJTImv
migGB6gWWuibCnkMEBrBjN2OAa0J8+l6ItYBzV76b6nDwBjlFpdDcjip+QM2V+yj
dJhdh1oIOIulPxHO4jQfXK+TCxUinPB4UBMZT+nTbAcmCbtdyvm5nsfk99jrAqwF
7KZ0fhwSaJyFc6xEg3pg9NcoJw2zEGX/AhjJM+Vop4f/nivws0q7uav6HPvKkjsi
yPu6VirtOxWYG2dzcBMRB/ijQfVWmVZnN0TqL7lnLeAAgfS1b1lIZXTr/p4sWR6o
3itGuy3iF4yKpAoNaznnmteqqjWHpldQWUL2x+EiLQTh+CNHsbVZHsizwusrHAOs
/I9SwFINhHgLJBpYlH91M8QL1Zi1ST/Jb83Rsmhfwg9WYD6mxBnOk+uXmJbI2S23
YNhxktf+GOAR+eiyMwCRG3OtXJaX6TavQwGk9VB59JDgti3nnnQMPBcUmnNd/+lI
42829qcS9IZPOWxleYKtnp9BDsO9Ds+6ZS3nvqQXsuN29yRE4K58mtEg4Sj+kpu2
fhB5PAiY6CVlBfjAZkGvLvDFcHfka2NFftGtyBnYanvT50xk+TRUdFLpRNdfFCL6
enyjPUYXAVGXcvzX4Y/UCGuh3HUcCnI0HQFSAkmB17fg/7XUmslroDKEmCi3/jdq
0s8376giA7xI+YU043D9uxbggbNwPN7T4FplK1q353/pBDcz7GLXKUpd7uC6N001
r7SYNixb+RzoClYAil5OiIL1nVuk+iovDeqHskGWrY8ehBu/9wbXk1tSY2qwotqm
K7eWnyMoCGE6B3e1TlXMVwv67LrhjfKP5XgbQpzxrY51kuv9L7uxue/wpHNA6jlq
nqihR/cpLo9LhCorFJRbN8IqI/EeN4AvXvOtHDeR/ryu9EkNYRusVz3gWKo7A0Ub
YJkyr6Mi4xr15nKyCzTtpolN+nkLSUzaRkuLBVcoGkWgHbQRcHDK+2FrlzbAxuVY
BuikUWOFQpvGSmUoTCkYmpgLtGpLctNQ60dlt4B6xgKTQAY8bYpBqsWuQLjM7DTg
9l6uyRWf7dEaMjsChwjFnIOCAgTBDgtlOMnL4NOr1qnQwuNsuHXwh99vewz2YC3h
46QFP7J1VUa77gjow0gmXsokDpi0kIAUiQp9+b1ijUzotpbTzVaNnluhJfAWnv1a
yLQyMyurHdbVyvwqRLihRw7VsYL3TccN5O20DwApd3Iz6aI57otjLfWJoEPwz57o
Ki2SAeSG4wsVq0FSTtZF/uv70nDqajKLnV/x+sidoGeZffq1z3dPl4PhAojhiA2z
P54eBl6B7Q+Z295kee0APe2rd90amv7i57h/V9MhP4adn9klpC1ML57JK8sEEU1Y
k28lrSbiqoie3cthe+HHtQt3wV3SaiYxk7iuX3HaZHLXeG2r+JXATeYqCHry/qus
13+wCrPRxZbb67pdaDf6XNUKSPnl3ii4Oz8fYbDN36vgiXBoBt0DD4HdggTzsaoP
v0crvULTkJrBLxE/p1tHZQZL0ZvIb9r4vIy74W8UrFRxTRvhmKCzTbMovgk9khSP
GoqYDzHHLRCRRxifoqz8mgWWaZv8nw3/FtcMO1RXs8VmflYUlRi3maUb7Df/Q/y3
BamjTXlI6PLJk9zKsUnU+or7O9tVl3B+RRDn+6q0LNS++v0809qUNi2xPiKXJMl8
T0hg5bPFXArEpaxbLvH/5wIxOl7QoHzq4gm62QObyjeYO5Oj/wwiDYFNv3ESxuh+
n6U/GBeGIsRftF3AmPIZOAp606dZK0SwiNWXA5FMq7etBQIRER74FM9HuV1/qXOW
3mPhxH4Z4pswjjHEPI7yjHmGiDQoRjfUQByOlB6Kmm94hp4Pcy0HqMfDeMyarYg/
V35+tCsAk0ELKsEsy8waLGV0i6tRWyhqnN21vkg4KrUezDVvJtv5ea5Yv3jNY9pw
BtusPnpeV4pjcVIdUTiSc0lzIUtc5SiP0REWjtNMS9TZyXGlnIz0xM6pI6FMvdtl
/RdMbxiFkmhqFlvCjZfhHO7shlwXp1YJbm3a4JaBISP1PfwEFZy/fVxa3Cs0C980
Y1sWSLrwxzHOROUbLLs7d9S/yy3UPpTOBYljnoAg2pK8+VuOwrLbwze/01jfdNF2
Q0NNYKTDi4rnWy5mopRNVpH5GyOcoSVMX6Eev96x89aZM2yjA+qqSwQGb+JaYbqQ
a0NTD2nnSmbwe6YAh2NSIRoQE6draoa5WS6jV+t9ykz+ABiVfBR00gpTlaMG+bhF
P296ZcjOLiLgSqyWIFyxxTh2fdz01O4tyukBho308rORAhUDQzWmHr2wh8KrsZWd
XdUbbBzaIoCXblm9T7q1j/ZDb/W052btiWy6xA5gIs1FTi1jbioax81KymzwBCeI
KvigirzWGR7aB0fJsEyfBBLSONJngs12a4D/x1YidgKycQgBhfAlTi5Y/RIAzdXI
UQloSGTOQBnLiGw356kHNob60jCGuXU8/CpuF3Ez94qoUuKrK9AlPjcwrZCRFSKi
jjgsxmlgsDVmsyj6RE7Doe8kOhlmCdyQQHpcgyQF/G5nZzJPegHS7XsLqzeJFh6Z
dLV6k8F3XMfx8A5q4O91uKpY5vj06aqmsQvi4VaLbqQwSRvLnK3EB+IZwYTVvP7f
v3H5R/eGGX4UxwZolKxLuWoBeoSBZBA7GGRDLVFKuCTKrkeS2WclA1GnW8QA/VwD
0EBKCDjAL0nHOSKWgLjXCKq33vrfXx9jtESmM2jDqF0U0GRonBOp14H7lKzZDjK8
LoCDMfb7tzQqky+Jkzbu53xNf7bFjR3esAUSviwUtXDrqkOpwITcbO/0GMY5mI+K
SNLuY0otIwnOzCerMWrMDvVUG/R3vZPFP06HI6HX/klKf5u2EORoj99yhbA4QLKb
PTCtViVPngJW32WyrxZxdpaqYiSPHsfOvJaR/3DNhNoVgw1FTwzNt8/mGTiLgGd8
Mrx24Nnj4vBKt54n4jVSj5loz8f5n4bv9AEoASDyxzNLzGwotUZTvISBR27c3KqX
+il/Be3RujjMM49AJ9VyRniamBAiAzs5FZAPXboUZglYAZc6kvk5xrAjYdo/k8QX
ej1XC6qY+gqy/j3ayUrVp8ARvlV4ru7OjUnH4SA4I2NBo0Z+KZYh/xhqOZohlLyu
T0oxbsTJJka6T4ZcDE0FSWzLIlgPbxqwXCSPHMDMhA4OXLrVhuGuC47LYBTzH5+M
u5yfKuiUoVhTUrHwaEMgTy9Ra7ImumU34b9PG0W8G5euvFY1dW4ZlpO3L7AMIA0v
Wh9F/zIygnwl6G5INknDVTpcyiausnRlltw1hnSBZqSiM2Xy7VJpKLavwL6E0TT4
aXO6Gn+WSl2vKaCzBpc4rzMSrazUJJImsWtkxEOwnmox7+0JhbcM7MKxavhsprBH
Bw/HtnGof+cvd3vLjnFPnL2AlBvqQEsD6fRAl78BMAsQ4ZRwGjZd3XIfydtknkpI
SkmHow/NQBAPhxKSuVJdDtDrsA4XGwyVHfu9NFKEgIPZJFcU/nmgcECMlCv8CRdS
xKnfzx1awfytax/tkhvOzQARcUfuRDsPuRYNJ/nyqLHpPFqZ8T3V989T5LPAdrcj
L/XRL21QDpWijDjtuHTv6arm6s216RPnw9LGgLYKYAJKBzRRwAxzII+NyA9TzjC8
vQy47BsoaSJG9PeWWhGGeSu+FCB2I9GGiC249qkn5rChGpzgE1F6SrPjDjXtIz0+
X4215wh5wG9j4XK3DKNeEYYzBnpSZXKWnzvztTYdPD1HxgquBBVx93vexpO9De0b
+cHUeUqu8l+Jb+zWXW09rkoYahwPfQv5BlIFL/FHf5Di7Pk24F+O5Z2ZOiSkSx6Y
dz2sVei5rO/o9UYi+w0hhRtxcPH0vF3dzxS3VvYJvGsK7W+z6fCxazgXu7/LQWFU
13vqovc1ihnjW/nBzpcv8Ti6FG3Sv10TSALdiETrvg2/TISus+/2CCzpPi1X9Or8
jLqZD+3g3jnYDtFI4j93a7ucH5a4/UvcZQcTon7J67lU/U4sonOqsmgvqvGtPuU8
GZqq5g7pd9wRI4M6yX3jWhW9wpWbqPezGYdPlFyKAiwoIbbSu+s9I+RCKzbooZZ6
20s2h9fX06R2rQNo35lRIZx5vcCkplAl+kpnEbygGEIYKvHytiNJm/Gmk5PDaB71
tidOYcTndeutWsFWBCsMVi2fL7kp/9igmjXm+dT7AoVjdBW8c53gaT+rsHGq7aCG
4EGkkJGm+Ev8Qp4q4jAuDjT+OAAe8Y65kbrSnNsODsgj3rfd61Nh4yn+fO2kuIyG
A9Izl0hIM3d598J03zvCKhJJCOD+dXyQKjawd5Qaxtif/10YCAqGZoxZnrZR+v5/
96QcypKTV1EuQe9xOBK4qUxZAKZecRD322jUUEc/GGy1NRF/XUiBqeHhBgdOv3Ho
gzVPSbUMCKCYGlpzui1afTxBrJKGu4UamITX9wMPBuIm8popNP5wxMIAI+7QadzW
x/ncz8rkfnRDS7VO8q0wD+y+oK7ptRt2Y19TOl+PRJ92+645Db/5x0viYOdfK4xT
H/AHgfkznAVacYxYyRTURe5imS3Bm7ZsyzaJ24reShNYfTqRTxoGlnp7jeI5Y7fO
iG+b9vvsPU7N97+DNDvY3wCiumUu2MFkUtN11HPaos+YbPz0xoPmiNgNWM2RR1Jm
NdTiC2on3qzi+b3mdFrXQ1JjGneaG8W3ZND/FJuJTGJbIp09XmWsJs+SRoxARV3H
YFlF+Tp0S+T6fXD1A+EhFGgAhgQqqe9Qm8Y9bt0OIL27AnMP936BxELV+4OoAO3A
dCzS1UvQZ3BFqwmUtgRD6tLrj3pp2nCZaEg5FIk7KU+ofz1WIAx0I3t8oUFR/GiR
MKSpUHQq8x/V3id5DLeZQtbSFrMctTqwkEK1WEYkORyDXcHvy/jOvT5GsfvrxgDq
fccbQW/XP2Hi4Z/R+oDmPGkv3hL3tZKr47715E+KNuQ7LGGcEnqR2zqTgP2xX9C9
hbOtq/qZSf/u7Vi7u7lPMEKjR5sakX1yrJj8ug6IplnyYhlxU4A37nNmnJxfIMU9
SelBwUMVIWCHZJPThFE+S389lJegaa097njv4y7ZAlMfP9SN4CVeA56MejglV/kQ
terM/s3rjQLJbGmtSpy/98TmxdlckZtrZ+oTGWe71XA7N72Otcd3cPP/Do046vST
68hjL09wayYJXA0Gy4FGtGr7vZ8IvKU+deQQh4VP1ODw0yVrVk9X3GTT/4Ju+qY3
BifMai6h0IZWQ/FjglagX4wijUBDEN2lRyqg3v8lUBuyAt4sU4OyUqc/u4N1jD1D
biaZJwAj3BazpoHvmuAP4YRNJSRiXVlAo6Z3QQKg12pfnweZomMe8qNHywvLI7CR
b34BQvIfw8fI3s82Z4FOe03mFL6/dmZKznNvhmNpMR5lsX6q0fYhqdkVaWnEnYUs
rxUzlwUTeh5CeRc/cz6V8zLKcBt5Go+SvKFC6J73mACNoyQKTfkEBGuiDt6lsrCS
MLw5bRwxUJB+KUX3w2LOUUA6ahtHKknY1e0Izp4GDTSR3cR8eYMJokkq1myD3zfH
Lh+NRVYaL2LlBf3xj8f6cTjbT6xWDI1FFk3fBiOpbGc3dJ8ru3OaTYSS6Wvl1olF
EiQ9ZVQG97ShRWlBEkNbA1z/qLT/tkeyKijjR+PoBp01evj+kptzfnq7tobo1pq8
q80f+DQ+DHhU1AhtctsXg97lBWglF5iTaX2m6anrey1/oK8ZAQda7yHRn5zVug9E
epdYdkdZXGUH0WPEyk7hvxEW8ECrMbuDwL5+W0536TdKQ81SdesbJNfprphUkDKd
745XtWvXM/Shb3xIefvDxbbBsZ8mfEU7eGwt0MUGOkrwTZg96j3v6MalWIbuZgIM
Nn9Oww2kzJMIGUCltw8AMj44/+p30D8L/qlX15Nv5QRYtbwSiz/aJ0t7Uf52tCme
ByhhDrZO4vUSJLtckQG+vi1RnFjPhEFMHLrSDSzI1A8tE0ujZTsEkumGsfIZIiHd
fKAbmnlt8Axlu0hoIP7MDv+K2J8hhCSGYjLIU/01uCVr6AIY0UffxTFTjEjwwX6J
aj3lf1lKlFuEh+OYhhHXw6JiQQJcsLtlkMEerb2UTNbUG5vcuMC6sy/7On15P19r
mfzASMOsO8aSZWR6r6DTj7tVqYk4XilhOlrE2oLojgxzlHcTtKcJRYU/gQyyvtTg
0zNGI4LJLE+RM9gUu+AIuT4bENK1Z8u5ol+4yMWYuUyEgm8cfc/togNyUiNvA1qa
KxAU16KQBVhVD/a6ocm+/hKfIqx4QzBoP9fIXq8Dkl3+YRoptmjfT9jjVu1D9MRg
HDWBlcNKGW40wqHoQi+bT5VgQSzmU6gaAHkNURs7cxTg39sWNkTXhW9gfnbcwMTg
E3LkE5/3P65dKlrlYXwHvrL3gISimOn147p6hT9QmVtegI7Nv6RbHcesMfhwAIjg
jEPk0HKhDM/Cka+lX9Az1IsOhRLPkE4UcVjxIH+LOGCKvbwWYByYb10W48AeDgdU
sNdQjRFS4NgHrLrT82NqXFFIOkKut+oCRgtob9oi6mFZzxQNJHNrDU0jIIZr/fMM
xbrZZrqGhrMyzYmYFLiUDpPqmaJIZBfnunH50+eXnr0y2dbAZ46JP6iXAO0GkzOH
2KudKG0CX59Cm61sq72qbF8abalmOXvDzf4NiFcUAVXuj85I24TsaZvXorQOvWba
dvZq+PrG2MQSgehEp8LhdG3COtHePfCT1J6Apwvn/SBp3Q/02NfuFsVcM4/ojnLE
tnrlKNCsCKNBcviRUPsH9n7AC2CYl6Bd+EKbhIdmw0vSnrmkRSSlCpSTnYlhq3Sb
jnNt+NpEK4QhGchluW5WoPRZi/KMJkp/yn3nAR2K+tUbbvbYFNMTIPJlBSa4W2ri
j9hFvqukM+qUsoaDcOzzu0wjB1C1we4SyjerZIhIUnRbRep8UYaUmHSXblklDVWX
pnsE+8Ui2uStdEftvF7ulS8WTbaoRPFC+pB8mY5SONnsBUvdbqFPSOX4EVWvvwcE
087HHn2SZBlyBLFOrNjQsbKTIwOTrr3NaNOTimXZcYQr2shwXIgWI6CjNmF4bglb
TyrDhJpWpFUw9MFwMVCIHB0WXzBI9N+ak0MenTVFcPGnW7+wukccK49+8Fd4YdKL
NUhUB4A/C/ACkw1vUNk/5gwsbiDBXLIo9OapWAPAK687Tj1Iht9PRc1hnDGtAJaG
IJDuRfJ+Tz+XIAWZ/CVI9cco5EaIAbfOhG9g8M7XIT3OxPCPb54fzFjhtnjaO1GN
ZFOV2+ktqGAyAB7fBuFo3fd6bW84YbIjm3outamtuO9/j2aVHWa9Iqgez8CS+aZm
w/jKrj/Tw1CbgRzHy6N6t7oZSGtirIZEeKjTHEkmNJ2faLr7LwV+l5qLgix/CZ4a
EVsi3vaobAhmv81GrvdEzryelF+AA8nxi0kG4rBJzQeAd0zkJXzCZhrbCARV/2oJ
zmx6a0o5ix3wylWYgxqr8Y6L2mSNeCSYhgfP5MChKxKcjL/IOXZzhQ81Xb3cloct
HnRA4usEmv7QJyCHBRFhjl/ojSDk1CtChd+fK2zLaCqXbW9trNLDgQXMKbmzCrzm
IiGqsi7//CPlIwAFN5JGN+NSaOmLQdgImCzEUPCCb4b5SHDJsIGMzYU31KvN+LyG
9Z/dvcrvtbYVtOQsYp/m8gWwQzNIT92D5j3itjvkEff7aDREvGJLVcJ5rVWMU9Tj
/0cnK0uZGM8JmMAO0ljwJ5HU8eGqfY6DnfeUXeKgXcaBnESFqeg38PfwbHxCqA2h
vP+ODQDfJeu0huXfS0DpMMJZR41Al0aMbKBup7/rYJxBriU60fyp5nDV6aqOCHkt
+mu8mW07MQ3HR6ILeJ3wELWHglxY8WKULa9A+fvE4ONTNymoiC1qVnO4zxbKrCyS
yC5Uh3PyJISkyQLMhXAkvK7kztoSmXad8cdVWBZMhWYnjLafIiX+IvXAHhvzuKg1
AYN3+UUzIS9uLuUOinmNBPbACxqvnPveJnjmFURc0si7kK32IIcpPbZp+y3L0yBg
/Bt4S9Wh3tdK5BZ8LbLLl8cWZ8HoQwE9M0pqMSw5Wlex7x0yXE2OPyv25bdijWd2
HNiJKorKJ6CgW4lNg217Z8W9dSMRsBkoMerpykHPEB00167Ng9R+6BdNt03I4CZw
j0Q0hqp0bloPoPC1GYCPDsIndszGjmNMbJQK7OdnhPU4jLM7HGCO03lDaQEiOSzp
WnEYw0HoYPed6ya51ng5C49H7v5SI899n4xFKYt4w+D/EdgiLW2q68mI/MyZkeat
hivGWaB3mdI22qoFN57HcHhNSCv/16n4XY1VsBY+WjN8mExGUB2rWCb+SvXFOozK
NA7ST2U9czt1p2HxJVJDcLa1fRsntvvheZZBuZZIZXhzUZFv9DSLHf+U62OV+nnF
IEdgpws10UhVvjctdb8v+lSrXgL4E29+Bjs9vHM0aVsgNL1zla3SCj8eX4mao8q2
5rGv2DjuJUdnTjg7BHQicRuC8AcO7h5texaiTbAZDrTCkXJJVJVaX+ptQpygyl+9
YeCVcOSrd7z1xPPkb89umxZBqjTm7NfcwTNAA5fxULLdHowh18j7EUQB5yfwbMmt
kDAdOZm4Xl17F2cM7KR17pROVGysERiQeY7TzzQtQEz1lakczKfyiCLXnghgyGAq
D5knLIp/vdZoBXVTSQuVLDReW5pwrmrT0STCOifRbOtC8yj7BH2uIaOKNKHzqtrt
j63H6IE3cr3IdVBLsWgien9Rfy7kosBjg/0OfR1Hxf6Z43Vsm+KoH70ycZYnn6Ls
ASyHHCBhqbmf5J96Sp3u5bqldPj5u64jvAUxc7xYBjoTc/j28tqdZYfQAuN2NOtS
AXD1B1yECzSwEAN0FZHGHcCBE4ycVSxOiaRbu9bdBMOwyucBWM9UEMobh0R+20VC
LeGMDZPxyMmSTmMEAPr7LIsJMayMs26MPodGJ0bX500s59PJ2o6X7otGluyAGhYd
Z0uIDdAdEKEVlIKfMpInN1qIu7WlGBcLwtodkpOudvXqRF89QKXpiYc9lLu4Ms6g
Iqp6nMrX9AH8w50Yj4QVX/wMiFJ3wDjblQXKxTcUDtz29EurRf1OxYEzizAdQXUK
JTDOulhdk8J13rJJzsUVkZ/8e+C79V1YLdo4Nyx0W29u3VMCPbEcNrSbLjp7WMsG
JbUNN+VSf4Nvf/w0xMC3inZSKmvYBLw1bimWKOfPrT/WNRrLBIaX0DkhwZtbkBz/
zIrp8Yq1oHgQNbY0uD5WwWEd1lpRuFN81qiyxoozQ4pDs1zpd8kFCrcXXcffF2gX
hHHEhraENMEVk6jigFSbrelCL6b3M72z8DmI+ro5DmfngLlaNNAmycpLgiRQpYHZ
xho89wDNKrvmg3vmuht1mmOqokq2mzogKd3getBMKjyg4QhMsfAG+vMTSBG1R71V
396RVtlGL5r6cTrjSOVOHYj9WjOXjylzrjZV9Vd028yIWNCELyyQlC7Zzafi1msV
KWvflW4pTSosHB+b+9V0U8cXFX1ARCDDKmOHhUtQW92Qd/yDjMFhKjD+xSbPj43G
xyNCB/vnjLCOig8EjF8hhsmGCqiEykDjLXRu6yLH0zYwEoWkSyxd/5iyv65Vmzhl
dGej+CoYwwFJyuYi+wZKqpjWc8xja3S0RIEsziT335MtVq3nnK6jcX1ZAbiIiTOc
lgY+OLi2NdF0yeXhmY+eOL2+0CgSQmDDcujFeB+Afj6JEvF8UnFR2SuLW4G6QLIX
riI75oOCAnMyIdKi4IG2tx63j4BEuGwIH2U/P6XpRb50EZ24u/T5VwwZHDkV26Ej
Db8bspa1DF4w22Drg/Uu762Zq6qaPbCwm4jGHqaooPY3LNq1Z0Mdu0D7asFEobOb
8IpqGUupgMEyQUfx1HvknvgQ4C5jU5vHdi1khWlwqag05/HddkctSo3eqSIXcUtl
2/dr5eclsyrrHtqZTrzCm4QAuyE5djvA6Y0Uxu0pkw3bWQaSc1j8opvPrljWLyIH
76R37OeRnKnqPL09g0HY0lhYUbnUNCyHrQyWJHgjSenrBTYuJV86sCpejasCYqgR
1kFdx0rtDUL923+fKdYtl3bblBvYwpzN8CgiwXM/saBd1282gF3zqpgy2PfrVHVy
oaxpzRxduNN1KMSgorDCEv9tFMyBCj2wP+tmhb149g56sR2GqRTcq51+DdR2j0XE
eE5KQplvKleIjV+guUpcASRr9P+wESvpVce3/SNd1GWaNIcKJJosmbvsXx8OfF/6
W8sQv444c0lkyHylqSjtxK09VdRd7PCk6WfXksIFBSsKwA0Gdu27uayUnwG+UYzT
L3YzrCtHrHRZhvCjypb/l8BbXqoZGOuXTNcWTlmlSOLZwZyH3dUaP9YgIXzDpxai
dPORNBD6jhDs8zPTEIRhJFzt7z7nsg2oYVG+e/S2g6DUATP7QJ+lMxxP3PmWjJCP
7qNa4ea0L9lZ4I2bl0hvyzjf9/8GpSjZUj1msIAadxbB51ViZxA9hmq6/SvBht/L
jFfGagmj0u8/w+NiF+69jW/+T4iaPU1so9BLCMiKLG6AprMAYzdS9J0JOq4UfhEs
q80e+wQdZ+3AN93RYy+oA3QJ0OBucPOrveHEzwhpHIYu+remJcZ8gpSGdcTYTV+u
5q8nloALyrBXr1xmO3TBV5RJH4uC6t/WMj1Y69vno51kp6/B1qcWe/OvOC1WZhiS
yykSAOw0cBBvilx4r27lXoM68QwOnQUuBRzGGlMA5bzkD00vq/ahU35MN0VoV+Ea
aJgA3uBbV5QIVZk27bn7Bd5Vz0XPBvke+D0d1rx+NR1o28GZB03SPj75XsAsOln2
kLFSI8AKomlJJ2Nb8si7vy3o53eUs6WSXudUw01h4W2Svjom9QG/EKtPSMr8cioO
ol9npI5V4q59gN2tvaL1ubKmucSoqfgRDzveRiP4zvgqjXT5rOFgg9toHglaKj32
yrg53sESKfYQoB4gQ9Qtyx8JsWsQGhnNm+inzslIrFS6yBL6s/K2q/Cm/+CqDa9J
vjsErMu4BPR9Ezn/8v6+9xad3tYfliQRodz/NFHhbqdEwCKlf1kmk2eby2raOl2u
IJhUl7E0rjzl5/0r7SX3ir+L2wlTEjLg8Dqkgth90SEFej59l6ugB5a/lEG2U8JK
/DzrDtZ+GP1IfHl4OFT4OAIQb70Ybd1LebYL/A+Q/05H69xNsjbP5JVR0lu5Jq7Z
XUxWZu1h722MG7XWH3lqfANPauc5x8j7kZPPk/AI74+eRLOhfwgXma699qwK42Sc
PS6yO1yl6BPL7MLnUoaKL+HToUNSVSxEhRggHn9Nh/lYL3j7HM9d7B1w2Vq5AmMk
KZ67JT53bVMojEX8JISqPmB37iOkl2CkNcESLsLcomGSmSsdCBe0Vc/X3QQeb/4v
4HCfTEBOOQzrlmoD/AExzU+0xMYv1ZDo9wvbSEAQG3rEjLBpISfrraJ+27iTwJzR
ChnHBaBTIB5HFs/BcC+AGDuu8ZgD36sO2bpiIalz+QoGZeBfwPR3+Bc23pkCpTSW
RMIaIKWOJlgTkJU7r7BtXnenGZIDkOELOBee6BtoKAUUPdt+kC0I+OsNGQGhTLiu
kmr5mieawyQg11LvaLy15g94F31WR/q6woMG4zTSE4lcIXd5yfDxJ1v58RAOvpdq
O36pwfW2sLqwI9aAfVNrggBk8mYyxV8yOv3qywSp8Sx2hvQwLK6gA8wNsAk5gWDh
I4AVm/gW1hkQsiElZnVo5yC3Qu1r62toA0/sykwp0sNXsIJGF+C+CW6P6bd4NKaw
S8GPYKFHwvi1dpvkoPlEk89KiA0gbtyxYfofrfrchRkdSlDoeaUDQBfyreUP0eIQ
zQcEx8wycjqUUVoCm9z7Z5lWQ4zO4aSLlPUuR9ALSm7uNTC+0lxdHXBuouP7mcVD
LrbOiFhXAj8dgtCxc0nlzkPyHtccT4YNIdhlHbP7lNUUBzGJDdx8ZC21ZE+36aC4
POv3sgBtBURZMOS33k05bNZ7K8BKVaaetHJ7vDwZL6E1fvZMNMj/TPRhz3GFVNxy
I8Z7jnxfSC19EmEiLi/e0v/SKSOThCDwR9SQEMVUj4mmiShCk69+8v9T1qB99a1V
oqe8s7XUTKjrm4CmOjLCwb/AeDhhmlsuFWUC0Tg4bGxzdgL0qdSDM9mTTZ49EReK
0BHdn758ed9GEbACl5PuCtmn3Yqq+wReXETrpeC2LUjiI/5nKvv41immSsYVdj7z
72Bx20okXRSNZQM8pJDbBrBhrSkxiwn3ncsI+fFJBhzYb18DIDfGN6nIGdIVqJWE
SRJ8CbT9nUGwXXd6aLngfmAo42HICleqxZ4GDVDVj7gRZ0VqhvEl37mFzyzMtw+0
A6rrVax50RphiO90+nxfqVkXD0xVXkvW3+vnAOGjMdq14Pr4mRxXDXCCg38uWryO
mNTec0WT836nLTbU1OLYev2sOvCy9zN7r1fMfSSDBQF3WjxLQsRH1LK2ca20GTcz
irBBw4rr7TzLEzNCDIkFw8RXgZWsKlAjw9AOQk9NJhWxyzDT8TJR/Lly/SUXbjTc
3bT91txvy6Ca1uFzVO7PQeqfF86id+VfSeb1WxWbkL2x/b7mM25gZuXrvJvBlJiU
GNE62mAqxevgGFwZe11bxgtKWBM/gRy7K4dAaBUYHNupc/nr/fdOOTn38o4bmvsa
+4N8czwKj7lOaCrvLJIP7U5ZMIBTqTbSej1YNVAWD3va1W9pCtwkaFcS82MM6D/0
yqvlOZjZOnbl+YVN8J6156tFnQ7XfZT1MuhLXNaaDoTB2XgbqDYTRrFYFGkcMdCD
ooyYLUKdu2hfIWG2pwxhvYOS9rElJ9uyY7ruY3uBp0L7jyjoeAnnqNt7AEbvF136
Wg9yyrBosiSd7boP/NkRiy4ef8R0RrqrKqDDyKUcUWTy+qJk06zscHq3NDRat2gt
ZOFSGvAoDTgYk6Rc1wZKLzrG7JNcdRZRaEovfniBRnlvFzMTBiqYvE2yhDxFxTeA
wLtQzjMV5uVuCeyQ9wnYM3fWi74m/M/DM1UXpoxsKLhp+KEu7rBsB3acqgSV8ZjY
aRX2mnoMo92fptzV7AaRw3o5TfVcD29eTeZY0dv3L7YJi7WKeRdiWR8UOvXj/B33
fzGHcoyr77Ftf+1VLl04Ctide/HixbRzH8sOXfw6RHbRPDgexJdJuMmbuTr5eH6U
zgfrdNnwaw3HmH48wyTsKVutx2W7Obx/SxbVxPPiCj8dkyJ4KastUXWvv7mdZ6qn
87PTojdmJIWS4Rg0OwXYKJKNv0vBFAnnJT7/1xEMNVkAOY5imgzjuMPFkBvGavm+
/SoTyM+0DmjJ5XortU69DGvEI+5un5Wu/g6Se1WxqPaQcZtpIp5qDHO1xMJOqq06
t0jHOWUdhz3vzdOMLG9SX4lNM9oZmprL38g7mUzeDLinszOL6J82/OxuXYy9zR6p
BPlfLjmcAqXtVZe3T1x4yTIGKTt1kMGR1YoA2glR3m7dmD3CF7h1uaIoXdTxFTN9
YJ9C7OlgkgCNT+O1kSa9alBHSjhfQZmFN5lXJtIqbJC634qPIFWapD7eVHQBXNpt
2fBWBIWHfJtEC9Gxrh6XeYu3XVW4UPwUaN14WFKBwvKorv3P2c3IKZDIrCntyWmH
8noqSW9U4m7Nyw8p/zJyBrV8RwtpmcHmcWcISK8STsj4HyYYVGTQAFUZtt6nGZqD
HchjgTH7zGlYsnZzqZSQfELm17lgug9m4mwWa6oTkYMQvCRVWo3C4ZkNoBIlycMD
lE+c3RB010Y4TnyZDGnvNaoNmpQochIF14tYKy6huvg4JPqbRzNHhGsNXzO5ElP8
gXXrzsAPJfVaIpknA0ywM8i+EUBcWpdGWR3GmlaATe5+Kj8XcAIl1c2/sgUa42rx
mS+O0p+ZT8sYUMfVa1XD9sHrHL9XfLujP0r21ezsmxBAsUE+gVmD72LKggvR5L1W
3s7miD5MivXk9acTsbXcdOqNhOiiBy6XVLXv8gC2yE75YWfCVBl3gKl4kTFitzde
gvgHXkSPGshefV/nCajTJUoxBgteFzGWSxKRPQectMGaoCXvpO+rbYhvNE3wt1l/
AiHYIlsofXRcwtLnwhzGu1PkaAUfeXAL7WI/YvxBIh/GH4dptYdAQBS5x0aWrdOb
Fujy99tjCvotgDAVY7iS0MqCi3zc9Av+3GLeOp1nlSujPkaGGT2dgy6V3oHlc25J
z6K04h2CJtDRaVhPPP8onUX+68cLYmHybM/aDKDO3/V+ze5caYn5gsYqodkFw6+B
xJG+q0HIOnRjHkpsmXj4J79KKib0ucSnUjATrIr10Je1/DDoO9XfxSiLHsQUcIdL
CVrTK1kccrbo+c8W6RqgBlhGJ5mqtF9QRqcYcFMm2ytG05eLqwsRoclpAfgkEP6U
WjFYoJq0lvczE9l4hE0G++cNJomdkMxviUWrKnwDthZ+EUvbSus2CyTvYVXZq+nC
g5hnkxoxSm0rBp/MF3KkOwJvXg5DtgizbH4Gni0Njw4U3HpmiBHBNpISUYNvEHGC
95vHsgBdjXssuuS5KEoWAZa2xKMZc5v5ZgBumACcjAElVtg5ZmnnH7S6YZzZJmET
AFuWI2/8DmV+Swwv3Ndw2vMT0pFJoiK+nUdNHbseaGWxFs4slRyXsJrbD4zMc4QH
cgNV4u5CrZOwg5OlrKbHRfe3uTHrn0bnGMNXUOZPnhrROH7/5/upJcWFoqDrBQ66
CgoN6wTNmSitba484WUHsnu1ferxGmMr02Tyh/F+LN9MjQFK/Z/aiVcO5Rr42lnM
RtLoKtluVN51U0ZFIpBllSEYw8yG+ujAkcfKvxMphI0HqeSE7Z1PfrYODtnmfhst
9+tj8g+dPLcueJ6/l9nQB5mC5p1QopivS3WUvUSqcUJv/pJwmznDRteOqVYI482x
aOFC/oyPBBox0CvHpt1EIpdr37WcM5hrABQuxNfoNCH2+KVOq4T03DP2yPKCggMI
lbFjcIVTw4fHL9LdeNA0N3FD8aV6HokkXLM3R43BX2BSuz1SpIlMFFYy0IJ03VAr
FS6YrUOR+Wj4gcDViEClPCPpeojhg4BalVTnt4qr2aNLuQAj/qMnTYQX60bQNhQG
zb243reinkXX5Vg9bOf+aGUtLQQeM2yUw7wxQCc/BKolqNg62v42D2RV2Hc3FJsT
nlpKWzSb+RUl/IbaFCcLvIHvq6H0+1HsXx7ZqPhtAxdugOrQIIDlJZJPgr/fJB3v
YRA9ZQxPycwLYGnIOZHfP7pi5cnWW3XVSuxnp5iOpk3/nIQ6VtKac0+20NE45LWp
5yktCp02a7Tz7eFuLZf69aM96HdImmmTAGoJXe/KyaqXuF4i9AF63KOW0117gVn3
c5VB/Me/oWJEH1Tye4DLJZ7ej9sAnMAW1kDYSdqAzujIcCCzQ8YV6icukAhBe+9I
bHn0eRy2zckk2LrgWZldrKbqg2Tq89aekIV6FeEFKGOhvefYCKf6g5iyF/PRaIHJ
B0FKqN3gxxT7s2JMwqVig9ACUXDgWE2wO1nnwTCJGfIdqSfjPQTuyYbKT9mCgup1
Qc1V54IwO0HWj5LofVBRbfIXcAVUPN7TWDpfzOUAoT8KUkhxqwN5VE1Hm1RwPZ83
z26eK5HAWNASizlhYn4rnBMKXfeAnxsi4y8z1+T+Yed3CEbIdep2PxSZeUD2QRDX
69vGRLSDsw3ycBuxjr1qaJtlG6PkBeyh+1JzbSemPPWQgpInAATffGl3yrETFPwY
OCCxpzWgwI7HJXjyoo2O1zzaAMbAQnK1PvO+FVZgE+mhJjLzwnCmayxHjwSq+Xji
hKd98TV/Ux7xwmSHf3K7/5nj5W/H83NHiktrLY1qI7ZSet56cqMFmd7GtHA4G2IS
xQACzgtLvaI7kLUYQU8bS9SSfS/bLhk32pq9NsrioL5KniNR0moJlpuSsMX/DiQf
8ggCfq/tSN0E27UFa99xDftsPQfcDO4f3H68Js1HhFgRP7ltM9nSBcaZt0w0B/B/
DcgjgwesNX9NSUzVMn+UnJ4VADyOgnkYrYrzZbxfcnv112nMWKRxHUtsDJi1fYKB
ru5jEk53jwZfeKYRSe8gNe9AfbPXMpIanlCIlE2CNMSaUIMzRzKNv7RKpYQ14I/T
fbT8JhYZjVSA7yJN2rwC4sQwOkR9pB40510dEfwfZlNUtR98SfdyrYMyO79zzUgq
UhdLu3oKat9DwqXfISDRbeKk/bG77xlYw9Q2ZVzOPbFOz7NGFZCroh7FI77e9bsw
kfsPfaDbwacEYuvoehm7WI0zif9fyEPKCvvn42WemdqjHfjcSN2Vzf5rPKPCFyM3
L1n0htS01KRAb+YI336SeVXvn2UZOTS2bVyk0EeMKPQS3jmpb5046mpB1NpQXv9V
OVCzj6nS0s0WEX6LPS3NioL4MToB/KY6tu6S9Csoajd3NYBFJF6yMYZEV25mGNPN
1Wo+GdQyWADm18ULbyCEeuV3b4YkA6Nkz7yWv43vZzx7jH8OsB2uJbEEye+MUol+
p7fT+PvN27X4FpZeMFQsga7SCGlpL9oKTe5Yhn674yw+z1vvMvUO3wZ9MarfN+UX
SJg7zaYqXAvCPQg8ahTYmPY7gxbO7lIT/VZ1IiVBF1mMM8Ic+pLsz7VLSKwCwE1+
4FdKur/tt0iXkKJeFsn8cGCqovRmq+C4Hf0SY6AUof4Jv0lIEGZ6Je8IKul0TS7x
jDT3jEEWVkMMCuKngmMybl8e0lAftbnyL7d4EHIeU+RnrQCHC4QxPWyNnI3iWEnJ
+M+6ubmD21xViHrs3uzqyfuU0x33Bds/ALdiY16qcQV5oD7L0TPghKcrLman0m7u
m3R7g+/hE917to+/9Zd1j0zz1xMme2kx4dqDDhUqAB2PeqgkvsgZr49VVjyqPJUz
ZE3KiqeM2YNZxua7IjbYDqNjQuvLXYEb0KfYFCQBCWbfHUcVzGmPr4Ap8TpxDXlp
geS4mmGYEBQXBlIpFYzKM/fAw3AfkIcNLED+9RoqqEjDjLaBI2zIUsB8fVFbNynf
UReeb0SBXWEbOW8LS+yB4w5+ZaPIle90ldXFG4t6GYD6aWStz5a6p38ex7yDhLwL
ELISog6gOQMHdMzfGyMUKByRxmaYw+trgLOnWH1zJwKG5pqTxFm5TpCMrAl+bvPf
gdEZYK3MbeuDA2BTAFE3xGYeHWzXvufUzHNIZEHROZwW2XzNIp88puVs8Zn2DAW3
YQ6uKmTTufW1rDOMvyG9sapZzgvqG6H9YSgfNSMA3D1ht+nonlXfVr+4bNDrYw2/
1He7IVl1lb6NmLTAWPeWKPSWlbkyxbZB40UkYnPOai7cGn3/8tbNmo/AQXXJlEYQ
nekddRV/Tznj/L7XRyZvx2h5dKLnOwQQY13nBZAvS/gIu2uAf1wrG5EZocA5jfsz
gbBFygwjj7qTxVeSooAo89dkTIKjX+DJeksAiVhaTZFOzd12V8WjL7FO/KMjjdTJ
CCcCiaihbUrABNix/YhqGZiTX1CSR5E/fRG1HTCNAD6psR5Kr8ydN2ilA003NHCW
jSklzN5fU9JxG/XXvKM0OyUkyH90EcQIqF97VNeR0kquQPh1w7tpSUY3hQQSUoxJ
LKdD2GOSvpkKDUTO8K5SOb2CG0vWtSnact9m7X/plX6xkJB/Y5GlAISOzzJYFR0Q
2PWJJLTFDJyjCraUXNFsL7/I7PGcySbPLEIFJFDeGkf0jUCHKtsUZShrOV52pgC+
CeXj30XyvbZ6621aICccP5vcBK/Y+dlcq/V4GdEaqg0S7YJl1sM+q5W0WlMUf32v
svNoXcoZOyUcQNgaCCwS6eDBGyLVNWl1pf/YgDhLdLuuhJMVhJQFBeliCf55HBad
05CzCKyRWIkRKix36owsSF0Lr1Z2nF+o3UpHxbH9vhHodGMvFfW1Bjlzcs14MObQ
PvbhA+hjV+vA5XxlSdf7+NkpecsYUcTOcUCMhaNgoD4Ff2qe6gsoRUoYFlc2rNOe
2FEIVE+e4vyZO0L0OeJlYaAAi2tnqA1D9ahL5xazJZ8Ncq+XjRa3I3Oqh4127GKP
g0jVD/aXZYB9fgno4/S4YAVa842tTr1OIioVZMLmot+gqSVJxQ03UZ9IeJ103FQr
R/iP4EHLLUJsgmJC67IiiF1siljL9V0tKSqQWGSswUbG2J3N6BhC6FQAcf8Qr9KL
YhP9tD4I23e2K6X2zz3nfsvl9zFAlKdxf55TgJssYdf97CS44z/VBANhL7OA//ar
EXUa3EQtOp/BMFa5HDvR25On3WweGsMWRbf93qcdkKU8GqgTbDbRRcBINjqb78YJ
TpFJ+oUXPPasN8Xz4TwY9RVB7QCaS4pthIAE7f4q0SpZbM8AS/9FZZas6pKYufDh
LsLKHWedNMOvYMvf9uNSF+LmiUsmzTIjQhco1EaQa0+9DEUOhnmzCDmudbx81on8
9mMLWJjyv1X33+Zm6oP0/skSRgLGfCIGTYzZvnE9nNKSc7kZfSLTfzueMfqTwneu
fhbuAeK4/ubZJs7SPW8NT6OjAIsSVwH5t7GDEc05w2voKzsBKfNvbOt75WWnefuL
saLpgoF5NM8QOvckIeBwilYqtfZM2VLbXbW05e0fCfpf1E2z7c379tU8kUZbqqwa
eTujo1R/S8ENNPxXvi5IcErCG1kG1vo93g+apUAGWQXoC3sy/svuTi8x+ehmQV2B
cMseJxLGBBUapJ48CiBzop+GX7s7nIYPDsmlIPfJe5Bx8Fnchqp9NU525jJDp+p7
zC8+e0iNDJhlQ/jJhG5NhxhUONi7el87zZOi4Uk9h1bzChSklyQz4VnCOSOkQhbz
qgAV5yWWOsRzsDeyyyWE+xCwoGQunH/nTFDYpXSW/48v6PRZbD99yBlLjFxIyB+F
1T/G5kAN3LdO9nsEmmGwNfbFZUnDcSFtxWzHEo9e8uvklrubedil11rPWqjlLDhk
NUuXNgnm/p9yjZ2+a2VLcneD6+VCV+aRWFuZAntbEFFK1HNiCTtYk2onMBmi6/ot
NZCMhsvg/wIAglJvL08KzUZML9vSzdKQUn2EKErkiRWsNI5X7mCr+wXWRY5bDBEy
GhBxjNBIbkrSwoeBFcHDGm0ZBPO2xf+AfcKp/7qyqpyFrSgwGpGbe7yuJLCW3q00
bDq4ikx82ST/p1QnXUfsrWsNLz8u3LgQ98ikvnzKue3BqowVd6WPsVgZMf9yh5pi
ey1ovmhauZpQpsD3h5imOSFORlMxIugf/F741AIq1rStdPFyxEIRRZswwyK8frdA
jr9Y2UDtl3BGo3+WQjXZhzsRwi1+DeNong4t5PZ4J2p65bmmBobFa2jw0Xlcs/rY
R/H4HruYznIEYmCqcTPWrv2RJEuUMk+WHZRBwxa4RtmjYmBafpy9EuukNSvUbRuf
fovdxMf5yeGBhh2td/DtBqcCegRh/z89n+ujmCbGb4PbmT2Fm5aGX8ubsCmZ0ysR
EuWqQtC06a5wPvAWqPlekcWpIRVOe/QaapeB5Cp1xU1+pME8OtPyvQIyxTh217Q7
1FY2tEZjNrAsJC+YwVe3pBQtF5VRWNDE0BhMmcwpuC2ztrUoVaoaq0EmVrgu5ghY
k2zFKE7lKmN6SyRk5/A7KjKBRraUqCPBoJ7SSldm4RLEqI3mjFMj0nQlv9ANQ/uN
nIbf+jMpk0+yCkUfXRlhnX9xEQW0/bqgUp+3fQOYubZTsPFE33oMjCdIBrvzVub4
8UAw/3hUBoZO+N9RqbT7BXxalu8ZXM1mOfuKIduPZvn+w7yXxogzSS+Y80TGnJt1
woZfoazBHnPJyEQdy3DHmi04iSkUU6W3r8/dGYNAgtkUkINjeMJAS5aZLTjXia4q
`pragma protect end_protected
