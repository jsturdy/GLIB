// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LN7N0v6aan8UphjXgb0c/tLMmQWeE0SLpmG0A2Vsfqygl5Pg5Mrf7nzWT5znGwff
rKV7vgSXrc2Ln9mnCmL5f+wtfMnvxkTAlJOoCDnvXr0TTympUVi+pGSLcpSyn04S
X8XP0jkCcKjPvfHksyVXc8mBPRcYXqfearQp0pyAJ7c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 75536)
QXN7EQO3hKrQgyLWwTMfcXbMhxaNezP3lftkp7kKAa8CBVoTHDG/zoEuvnOeramG
9CmOaF0yyBh8cRpRRIynZ9CQgdB20ZtZseqjxyjA4a4tciGyJw72jpF3qGCh21NL
x3Yzn3ilqUxtoiJgFPCkjUfz2VqVh8NQBhf1pUSUlnixGpZ81JDsUTvUNkW1PZZm
/308x7PRxwe6K0Uii4TtIvX/R8kpBV8rc3QaGZutkFbwf6GCfv7grF01cDiGjAEZ
b9vPYfMc87lNrM6DCsdoEPIbBVxALtb4f2eTEZaJny5dZIak4O0EZ/xChFPXdb8H
9x8hkYpFCnUoOOaBfzTptyAS/lO1fVchrJE/jjEYNd5+UksH96KLmMEg/uIWk4Q4
nUsT+bWSNokB08+Hb/QUxucxT07SYkGyC2oLO2bMwSU92eztTKQB3Y30FhXYxf8i
8vOI/lcYmirOLd1WvaWawoSOOEeZh4nB3y/5GHxsQAdGxTLgOIWp+vEh7/JCfqbU
3iOXzGxguvMwyWOyRGGffhpPQgnc//5KGzwX0Yb0yNXFppLsDgDRhdN0Pffb7qmL
XLziFQCEzx5fp+Gxo8kHu+iF4pGxf0+ljIGNHqM9jdaw+FRtelCf3wQZTOSeH9WV
DajR/mDE7FM+9xNR5NKjDyYfHXCFKFmkRBTxLUZzdQ7hpWEMj68CD3anRGZPKtg/
v8EPliJYJtd19pSA6+4kibfZdICRH7W5OdlVJbH3jzdkpbi2an8LlRwPMu+1d3V2
pvHBZfvyXCFkqXRa0abI4L+lgi5W3uK8kdPdF5Tr0A8P3qVwBJ78ZAGG4aSvBPdn
WfqDToYFvLPN8EFm0MdG4ZM/C8fNmJvIPyRj0Weydv42BxK9wGH7ItwFaOF0VTKS
CIGi0ySpg9cnPN8i7dGBG3rH9vDBqFJzP28AQcqJgxcWSH6msPacTRdkdMS7begp
o3ecux8ghFrv/t4Yk3r8rxptHJrViNG3Q1WAe2hkasG3ZJ/2GB+dFE+5LhP5aRlF
rt6OMJfWg5Ea4vNQgbL+BYvZLxwzA28tVC5F+ZRgUQ3r0HuJMeOTPAX4NQgrTh5W
0r/0N1fWkCYw02HlpdiSD3lCXqSHj9/xZBx8mfCkXbftsI3ZNXkwT+BfXLINMyWe
ftsDaq9+LCR+6WVei6/6anMGTZowoh/WVM0mViQVKGynmmoB4Ki15awj/WnKxJeB
EJq+EWiC+MBcY71ehPSa2X/8gxHwH9PxUcx2fsfXaHhoFp+LXuFGKs8CQiD9Gt8W
0P6JNxPhOqddIYk6W308wbfl3hR6wFlityLuMqijUwfc34DGbRe+ylTuKlIGOGOc
uiEZdBZYO5LEjF8/PqwiEpcCIrBdc7XQIQevHkNGrK2Yjlh75QeQ+HNrQr42UR+p
EfzzyhimAgmqPR/bk0XOq7QgpvBgNk5p1YH+deffKAH1TKYor82BtYdm5Ihsh0fE
on7kCdiHxEsqsxQGT+QmhTkHoYOkYozhsJrxfncZKKxD2tnfpOLBHEolkt8DgBOV
rGQs1pp/RZozDB1jywj4EvHnhjY31mfM4Ne+TdYH4Q/LbAJl6nlfRmGx7rQynhwZ
ougklEFfVI7S+KPui94FJBEOzXb5eMpe3Re92S7mtJdYenbYWbvU46SLt2GMSItb
iPdntr5dF+zv4z5Qq4mqbYNtzqool2NXDJRz9lf4n2Bk3S/3wYO80cZv7w2OXlxc
GYrJpgw3kuqORymROZBYCv6H5Sy47znh6uKSsehgwJ16liV8IdBOMBAqzvjdE7Bn
/+qwoXCYcQJ6qN5+lL7CQ1lwSnePQTjzVGbEr6Eotxg7EWIJFPXHL1EOrBOHdUW5
jrcEl2E3knagM8VimfPfel1mmktPCIu8utdbkaEap6c+EAZYpS9H/jzKU0R4Yi2F
THVZ5PFp95PtRJ+tRRvGKBUxT9/TQZdnZsxSCzLs2fncjT7mp6Oym5ZjGEPXOR8s
QJRJMEtS4TEApIE27NGETC2YWthMwnBZgXY4z7OTuUJEn1rc177Vj3/cQ3+SSGof
i59atFfi2QCupb4GXtO2IvDI/I1xkDxVhmrxzOIwNpWONA2izd8smK378WM44Apz
m5r0dLZzbdmk+nkslpBjM3XavY52DPlDLpRIOhvoDFPArFoZve5Bn3InkQDnD0un
Ud0d580Zk9pFbRayaRUMWa1D7FgiEgR5rjivl8e0IsBLYkvb9DvxEl62YqngPxDM
WM9riQvO9FlD8vL7ZUJM5oq/49wOCnWo4RWDpoL0bnTGn4xoBsePw5UaM5V41YYI
DodsIrvP5nf+odI3C41kLgJlPLlOzuyS+iPdugTfv7QITq0e4R5+zjQZMAwlf9ci
eBX6L8L/6JG8rpux8gxh5P2fWH/QHG8BbkFoBDE/IMq4pnNY0e0yRVhqgUtA0fy/
Gqth3fwO6LyAEjo6/DIqmBZV/PxBx/cZlONBALZdW4eshhCmkmDIupS79/3XO0cw
br8AThoJP3JKeB98aa8wUXzsS7hUHQMO0fwfOJmjaNgFsAMxunlSnfQGs+c5GIS+
k1ltAwLqWG38hhodn5Jwdh/K8T1CCKOErQ4nMB17zE+R8J9vSvf+lv6AuV1AZinl
KFL6+3hImuIRsliH3mSgz/jDafusHvsfnQWlczh5iaOKNZ/jOv1TKtA8TRWXJvAW
AUatRZdxyyrDC33EtGVcVjnrNzFOId02WszMyfqOcj0g97jwgXHsdgco0uqoYnuU
4zBTocV8VGEeMCXvzFlr06cpAcjJEiT0nqiAwM6Mc5Jc47vVDuWwlYQWn1B96PSI
JpIDgLI8uc2uNXKnaX8fT5DhJmZAIGqTcdjubyrlME9P+baIfNChrZHV3CVF7xaf
Qv1dznBDlg88mCcCRpzA8d7g2SwwBA5eEgEgVqS+x6jO4qNpfTiPVreG8KjOHe2x
9qAclqhLzlFcuLgB/yVSG7Y26JNVpyF7xBdWZUm4BdbFT3RqpQXOH3BHic0MFkTy
Lg7vAy5YQQFNbpPt2Ciw28qfnDGhgq49E5i+E6yVrqa5YwRIn4ogsFHt1XNlAbQL
0QAxRXTNHTIXjUgX96C8r0NjqskUZilhy+sIidReswGoJ4rbznM0NM8IoMEC92tk
5hN3MHh4LySKlz5rbCbQ02ZmF6pSErpaCMUh0fxx1cN+E11ASW70UxscV/JcuTpa
UdwrxqaUFcVrlgJn/6x0Hns/7coj0qCKEl+tCF9nW6Y/VJnDRr7tFvV1k0L1NLfz
n8VOCkFhuIBy+PsnOI9g3AVrZXYp6P4//zi1NkeeyQPbOVQCb5Cf6CLprC4Eg+OS
FsiP8u7Yf4DEPx4CDNlmHUzvGef8gKJQMOXovySfLBaPs6UlUc/pwJEHguqhkhMi
iKWEQtn0l7WkTLPSBLusgihhORRCzvA3hAlbrKZPOWtf2f0ldD/Y8tdabe2z71LL
tnmZaD+VcbixPoac30hvTJkYvppsG6crEEo2OIxzz4Lb/kaC0ckEs0lRi0l5k1v3
qAz50j9MkAjcijlios1AmQ1FSdvPR9Vx8PeyEbPLfVtbcJmbGRvSjtZKookF6SA+
iLYF8Ldi8Shy1CyeO0+G5kZ4MlcUcw22OkqGtoo8v53Ol7yTaXi8cnyuf9o66Iou
HGI+560MpGg+9mwWC2ScwZYrcMmgqTV2uZmUqmh+j3SdG3M3Nu/K+oIwPUuoJens
PoP7x8LMpIj5lNz56tOiO0CtR91QJOG53zGOZRwv2dwfmj/A5YNroiRH0AZ60vjc
QtW/Yi5BFYS+OttyR7/hwYwfYFEhcb1dC+UJX+enfAUOjZwBITK5KOcWBtpOk3YO
woNwhAq1D7ISFWxHDA83YMS4gfsEfydigWBujz5Hmn/w+oSbWHS7XOteraIF/XMh
u806q3RwoE50MRKQDMT2J3Bvmo4MQadjNBOLVRKEnK3xlujXuY4Sa1VMGSqDk9qt
9obs3n1RcexxHe3EAlSGBnBfqVLd/kLs5rsH93fXP1IRK1jT4GomvXVrXjVJZCdA
wvI1hFG9m7LYy+DSlOOt28ab6AsC0RoeFKSv16NZcfENk/COhnBdcJ1TViczmlAa
P6Mju+fBeSBioJ+g5PMxJAlnXSTV5iVTQOvY/xFNIXRHX7nXVVJC/MNtgPW0bk3E
0GxEsoHNbrmr32jyiVDr/2WUmHyCtVxeN4ojQVgFRTs+MafKkg+EBRpEoGX9pxiN
0tDX9AMn1XsjumLPMVDxJrv5LzM1IsFmzKOYy5rWQbhD3g69Mj5Wic1d1UvjbZDH
SzuXOBD11nVM9A11OUQi0ZoySRpLAQUQVGXv9KzWMd8PArzNmFYAdQSzJ/1j3a+d
QGYqnQrbZXAYGV+KTJ+g8F4Q4aLpSvBf7V4gvTLciZ9dq/eQ4VxZw2Ugok+s2OUl
Uu73jXQ9Fm1j8MKxiBEubeGpyqKgI5CsAVY9lE+ruNwHjApsez+IRYabaFaWfwbJ
ke+fO1/3ZcKBXBO0j5fGRUWNR8GMxr4R22N2/dM6uxgnGLHbOnk0c7pq4zMabJCr
9lWvADXgjFHiu6EqJOBDARScGxi0BgdNScUwd/QuMnpSWikdfWvln6ZQIVxLOJO7
Snowv2b8bw+ZlvnJ/qZZUz3HZWB/EXsigPWbahY3C77i0vz7AnLpUYLjanCzEQHq
ve60LbClAgS+NW11JxLL8RSKWjAjR0Bhjr3igNQTBFFlsPU84xD+SbQ3dTNK5ZsB
IU3CaAMEOqmmbaJxcwpl7IXpMisiPKrF9uR0Gnv2One1nKUpCAX5hSTWa0obBbl5
mxWVDMSzDPpqU7slwkOspUc+sBSIf6uYCQgPMN/FaNQKPjCvbR7CwLaetL5xCbID
PcbtHaPrLoclzrK4qF40xy4FBVwalUuz4p0nDj5oKJf4IPA0htoeEIy7epc+d0uM
QW65ztOsKP6r4NhB8G9lVVlyInVEzCYw8ng+VGgJ9VJzdgqm6yA7sPQiCyqZflhP
enTJXladi8nNIPWfby1AsI241B8tkQl1Ie1QMPUMWaEqJO8HwIB4af1MFcQZ5LRi
4LYe0l05iFbPk+hu8+qxUaCA4wc2JwUs4p5dLw5SffWfdIIwbSl69gqGzi1uqRse
PdW6+GSrkXYiJLEjKsx3muRLWo7LbcWLmD9+doXtIobTjlAP6Ob/VCU79nwaJOXK
9z4afKMhj2qGYcf1LVUgKIW7KeEckHtV86kMza+KRBNavHQdyRJe937/L9Az0Yyb
LOBHlwzzV/mBlJYhYnFTmOu0atpdSdfoccd0LE7pOufhIHNoMLu5QiOP0CIzQY6X
zcqNDgBQVveM87kDl7sxgT9OaHXoGxhme24sA965iQuK9CgrxQiRCFInPZHtah00
C2daZUOEsrBSIDBp7kV/V5lQ5ZUpzj8fknxgW3mkrusXX+TG2wvmfPq7yAgjKNQe
Ch7nqEuDFGzxTHlJinuTkslIpZk9Zqqn9ZspcM/X5XgLmWpE9zB6dad4zOpmC2ko
XxRF+ocSmz74WxKP5dPIDbIH3mKmpqdkzYEUvbTCpIF+QnVSnOsiWONz9G3DB9+n
mkNV6ayWzNaUGRRTc3rorfL8d3SszDEafhTcsc9M1mp0sY9YKHPaOxQv9Tj/yojI
Q6v8fPzmD9rCA5kXU3y5Zgn3CvKiCc3QxtN1wR6hVS0XaH9CXCXURA/lJDK4jea2
hWybSHh7tq9krGKywknJvKtNTLsmI36ifNlHiW12Ne+zprJuYPLltt3JkKzym7v+
khA9j96gg5mDcZ/hRzVXIr7+C1WWl/WH/dtCpYBb5LCa+bmjhujKMNmjflZL9UD6
EuuXrl81iZ7o44xynR0vbxDc7oZ4Kztmt/HR2ciPBFQx/67BaaFRo78TjxDsI/Yn
0gwW5064SUXSsE9QcK55TbP8HTkcN2K0uoS6oROlLxEx6ktExz9KMgM8/mQDByjE
ebMTtEqrR0QZNzJqftP4mU9UT6JthKdBeI3OM249HbxHLofYpD27wHy1KBPEIIEy
BzTvbmXpExI6+Am6vDn63whKPjiEHogt/PjOTWHnWaNV9y6JSVhC/IQ73Q1NNxu0
lx6w7SJDiLoxIFYTCPXFEXU0CopTesP/f+ieGgGTQwjbcB1B1GTdxILt09hDHUAA
nRpaBvlt8UshwX6alQeVl3+hvEO6QP1D+9cqcmibHdBo/ZX/ankJS1eUMLCJoW8G
nUUCKxjadXGCXKZVRueKxyl0CDi9UOI4nuTrc0pTn5XfHn9kYvBj7p3sBLfdCtiF
31g5lCM1UElllVuKqbpe4WwR9MlIBiTz0faQfRqHEcntsxQwqooQIFLfUqQl253l
tWN9XKISpCloHIIxLL1JTpV7E/ergE+anltS172d9LP7Y6r8Vq2MuzVUinNAUGVz
ME9jJAno/YslWGYoijdxpW0Dv/TG1+hgP8E8a/DhndjHeNi2D0b+IW+SFUAaz8Av
n+j8GVeIhuH9dMxs7fP16b56aS1gDqMQk7gK1Mke65OtN5BxNixDU9RyAzIORDD7
gGQI4HuBU8YbsEntmbB/B5iVmQRwucg5CP8paSdYQuUE9jP0wHzuq68dKtRDqX4L
owLDCMFRiWY9D4wWFtktTftFiyw12gsOQw8v5HkaxJUT+Lnmd9mdwoIQBm/+ggP5
B1GP/8yMbReGwde2FpahHRV6L5cTiPuj8T2Q7SyhBl+KfX+FD4xy1mXoNCvqN1l9
g6RWb7so2DLr88CqmHS79tMwmfUu+xIHbjRROTZaP6VTxgEQQW/KgOKi2Yuiehpl
7349sqMZBCH+jR9vR90yrRR1dau6YJijfhV5k76IReBoY4iOZurvsBLj8ZCj6gOm
Z+dOi8N20bzDQNhU+oYSN3ZwadorhZq9wNmg797zerCvsg6Ruuvgt4AyOoAC49L4
YmMCr5SYL67K8mGtj6XWBqNonpZoYzHAYPa0ZXOApyTU+wc8d/y3mT+ZmP+n8ogv
+IxyFY+7n3s6vP3aFQ2OLzJGl8AUVv9+q+v+gI5R0p8hIrdb/Z/XK3bygT0+qFkY
deVvtyPB7XcW9DenbAjsiobFPtBLc33auC0QWrQJzjOpjGH0Esmu+nYbh6+lok1t
fPSkREKvQEf3Zyi46dScX9m7pOCwB4TsQ3XJefVq3jMCsqY/rz4maUVK7rx8JznD
oejFc3Xp5Trn2LjfcfXdQ9oa+e8x6JaU/9ObRMWhX8FeMensQfklSlwuSCeZFn4d
LcXVt8kaeXhJy9EuwntVWbcWbWGHTrIHcP1ZTbqy1GVoFUFIBc75JCz3lY9ay8p2
hqd8yfnJHwD4BeLlKEpBe01Jz82acrNtj3yNlGzRz6xqtqhcQ55kqis0U867RArO
ynoL9Tp+c0MRAuMRYtVvFPg3+hR5fyHHYLzPPIevf3rPSENHuGBK1hDE7AzH5pMv
1Z1/02fUdSITWKqiACmaUkGb0QQbyn3CyJxmFt/8qSuoRBGRlC6so+zlbzG97sfz
A5O4/l90k0VNMJ87680P8fTZHoKpEGWoE8zBKCOSJB3m7si/O16vMqiFhhiQUu8H
fziOZWLPCfrthxoBoIyJdnwr136GgIGT2YaKnD8/9KufWC4y0YvY25cFaekCy09P
EB2KnlfSuP1j7WoScTu2rCnd/ZB7gTwLmBx+kutswSau+pSu/QiC7aIq/ndb4lIc
k+/RGF8fXl6UPxNObw4pqY5MyuS/sJFUhOa3IBDHRX/LAL5MOEY2Mkv4UYaqMnRS
0j7Z8ctVr3gzBOufcYEvcfkp9fzNSm7y3srQQ9QeZK7vp393C2E8hnVSoHGzVMEZ
gJmWUYCc2aJgGQRvtTKzD8GmFe6ko/00A4QPz8LTWtO7GWbYGgAK+hDwvlcMPl3f
CP14t26eitjn34ZXQCGlT/zFM8Ag8Lt0oTZDQ9IoLDYGX6SfRFQ5fkYs2rwWTJll
0CqPDZS05BFZgrQL6PdvNzW898aVKQEZqXmNqhyiBnWO3PPWmRahA8ACZcR0gicE
fwBpdCRu+OAaBQdTpF53H4obMa44w97A7+DfrPzrlckvx9oLWIxg099fWZTZYJeR
D2u2GXfAWEe1DvYekgdaOkyyKLMVJM6hwD2ddm+aBk+67NcuU4wUlXHeHK/lCRQ6
qYzltxFakRZpPZR/9qrNQOuk+S5IhLxrwNDtesG4WqeArU4R438mVAUoIEW7MZfa
59dRbfimMO3lcGVgoXQyAl4/48ebUkotV96meH5L9hbHGSaU9txOFVl6EiED/AXF
8kbtVthKz6CIO7hfrCV8JYAAAat6h8kx8JGDFP2MT8v0QRGxn3Qxx2tvRTbuZklH
EQLgZ0ktnvDoCacbeyldKjZUaOUP7UfCWudpPFMX4PUA6OMMpyS30OvvNvvXuK2X
3YyU3OXPoDOM/vq/cvid8ow67QcYTk245FYbLsM//+Txs7PkYAQxyxM6IUwnZaXi
ytpgfJqTWyMIYuKqL9ec9NgH3j/xLRb7eRmT8u2ZY+K+kFyyc7/BFt+rT25Kbbnb
galWTMDyF5e1DXhrwMMAn6Ed0+eipzD2a+v4jlYVaBQUzlSwu8vbWd4hAsXeUOIW
B+tjGLASjQba6TD1mO3a8Q6y7TX1RFIsjidEOO3l09opOzw18cldAz3+EhWIGY4H
vgOKYRnEDrfDfpvd0opFn7vKaIH0SAThItc5aLDCQi3KDXxpB8oe2mc2sHvuBeLG
qnhFuz9WMCcgiK2eT9Z1sRo6SsM6e1wo+4A9cnIHYXOOUJBsSzuLi0pwp0LfdG/Q
7BA8bnY1Yk0JqanxT12pGLPNvByurOOrYkCxFkfAuGnEeAfI1cwMgTlzB4oqB3Lp
Ows3J3asfdT34gY+tzBIPtVFWzkV2whSsRrYd72fjr6iQ3LksZQgM17M6ncnCjJt
TLuNhVXtfZtQ3+1fe4/F/A9Rm/bWxSt5Gj7ykUoaO3eb9vpCCTZ3N18LNkgdSSMX
nPVO2hPBiYIDyPUBOOy/RUFdLPpEzH0qtaZRWNAxz+MdTiK6FObk/U3TXbpJEAF0
PwRedbT5J0KPL7ZfyevLyTwZygMKu+jdP9N+TtiARY3QT+5X+5oMaf/vsm5u6uJE
rj1Nkbw1OB8oRNxLecSW2CFXu4+prbX3z6gXcGG+JWUExb8eCebSVhgca4C0zpFX
CrNGiO42v0ioATliYXd0SSwikwHi7LIegbBDl7ZNugdSV2uvpkrI9xBv/ET0FeQC
yo6A1MDqxWhPhiGUecO3sPdIUJBHBwuePuD0L1aPdI+0Ck5TSEuDkhCw1HXJyG3v
KBS3wNlzjtC6mpI5NgNV/aJ/2LTsM1/v4/jnc+VVUwB66S6ubkcUc6K0KNrgn/oS
MacIl7a6QAqepYnJpKhbv5ybOF3SlxQOv8ARD0OPsrwrTeV5Iy4BJNyisIS97Z0U
2FMKs+FZrXQ0WHrklqbQP63rbv+g6/Eq+HDe9lmW5DrXqvesKgO8PY/IQIOChVpp
JszOSrcDVP3lE1Ib10p5X4XknVvxHxRYnS/au5v9mEeC8I4bUayDZjHVE69zMcf2
cFUfH8LRAXIJzRihmjyJkiJC+kUGzBieLQn6LCQAbeLSAz6V0N3ubqSKPJ3oxLWG
cFyrcewsOYdTz5R7zQxGd+rwQC1S1i2AsnHEXMYW4now25mB7v0vnLEk19H/nPer
YOEiYlLgzNR7s1gKwRDWghjL+q7rOAPXN4LvaCpfU0BZmxPYT/9CgEBkUIrSxE5K
lJn/OEUv8bdl0p/LziFPQHOkgHlbP1Tj99z7YLckqKYYt/5/UpclT1VLS1BK9GEd
ZT3S5HPRm3ZzU2iXkXNT/50d5IvpVXdMsbLjxXi5SBSph4w8Cgtifn+KztAn4omZ
S6bWaDNsblVLo/cY+voA+aC6dG3qTLhQVNc4lPJalD5umups/ttgiYqdF1T6Ncxd
IW2iBttiq8DcaOEaizsDl0p2uZpzyQj+m64FmBZHJ7N2ypsfN/dZgmtlUrxOYXy4
29mqijO35lETe/pC8A0wkwXecvpSR3w2cZn6OlGPqMyKWtlazhD9e2musqiw0u1l
5N4DtCuBrcz6L+aHXJCyXkx+a9FzyzBPKw+fRA+KtFGvwDPAY+W4BGxgfmBXuc4h
lF55ZgPrINHjEPnQdGY1gPsAAnNvwArDNITZYwKF4MjtilR30vW1njhE1BRXl9DV
6EF95qGIXXBVzpJ0Qk2PVjbXPhmMWZpGJlmbvYbmD6sLKX5vsW4RyNEohzlGTJcD
5e540lco2KkqRirj+iGz3uPmjWQPwQcNCvN7hwCI2SoSU8IYvkeWcWiQGTYTtf7P
uUFVytEWAmOU8HeSxML1xdxWJdhUVsSLmVD77bYEaCFyzr0VGJBKvkvyVYYaJuPe
2mKcR79/d3deFH3S9QxFAJaIFV4lXUfli70mubMIiC/geIZGQ+xHt/bd5qfMRXdx
sJQMlOe+PIggECDz9bMevKLSvZB3zemT3eHnK+lhsDG0T5LRDJPHFw+3zc7q+NuG
tZc4Fd2VQVwo6IFdDxYKgrcP7ydN2dpMHxoC/OX19KyjAVKtiW84Vkl2PKVzOBWX
bYPEJn8JtLmuXPINQPNIsvL8mHdEO0WtuPY9/gbuCjcL5j/ZF7WRyVW/bTWjRrUq
8XJkYZKNhXlh7fGcVyPhHfHPzR9W63w4nmOra6Wdcr8VF1jX8IUuE4oKd3ASJoUH
kcD+Ms++H9+p+m6P6FFUTOHMpjDbOpLXKSbwgM5ycV7I4Od+B0ihMtBvVJF5Mrm1
XYtWcYPU7h3CoaPf2Necd9eHjzfwrlvXWZQzKu/DvaMbeBJccucdZk+5Fx6UyDPG
VUuIzPkdhyqj0hke+9XRkbkirTCjAc9otW8iickCknDWgl6D2DkqC51Cof6vz/27
82KrswWvcR+u6ksqJlQb2332plaLPNNss2XYY5xsHNuBAhGZHznXqlRvUhzEkIT3
4YSCH7p0BR9bb/5H7TgR4Z0olWVLaYgNRzIpbL2UxMtcy495nBorGmaJtHDsLjg1
kO+xwVa5f1SHCeasOtlK92d68xmnbK6MR2Hb5FAfUnyAEas1A49XaJtl+Wc+i40c
gDv1RjKRbf+yacd/kBEnrXUzdgeE78Xw02HNpjPxUE9h9XgBm9HlkzK7bROqmQmW
WVXzyrSvOJYPQQeVBTqfTsfkqvkqZAD0gelg4aI1CJGidLzk3RZhFTiZZLFSDMXd
sBgH+wLtn8uATdQlo0ioKRKsIaEllINAEBpoiIII7pKT+f0CahrKrWXfMmVTdrVP
aPkypzyRv99rrj8eizRj+Q+aEJ9HChUE4LN6/DQfRc8NZ8ZC4q3aU9ohdvipGcSd
6kMuOGVUvFgAi8sZjHW/uLjaZZ3VNLxHU3gkNsPeh9WuI8nW+eyXG/EfrkRdjwSR
rcyiCbNDRefHfCAcGSdbbRaDyEIKjJrZaJqTAYZuh0rvXNFSqwdMEwwLAyNCHF+w
AGrJbwvynkCf99Y/rxM312F8sCSwO+ITkqRXVsBeuFeYotNEDMsxBg7z5Ubax800
fkvmzp1fLKQdymAs9Z4wtM0fg/d0eVhUYU4BZ5QtneWi1LN3DJvPpYaM3Rtwvxr/
mvYTqqotWtGlux7OpRYKa+9q5iUsUA6dVsK/ffWa7y8ZC1MtBA9tGpcMKJRJhoJU
TlJ9xUi9wsIy8ZsIu3RZNUhXAabhy+zquYQw+qLPobms0nuoZneNKjIUs1AlyYpK
QwFSp0/gNGtXsO9xuRmNrNTx1zuvctOhJB5osjtqC22dzVpkZ9XTKG8amzlXxU9O
AnCV9HRFdzgaYa1CVKOTLpGspgxEesRinsm23VJDZQUI5d80gF2hAVd2OLIciQQv
zNpnUZ9WYKHrGIRDeAMgcunaQxYIY5/WcyiA4SazioaViA3W1EZddTm9bnGxc9C7
z1MoynC5wUHoxmBjpMYWjTmMO3zb9z4m4OBjbtLCKXjaFs0OlyubSVMo9UIE7iDC
R8R5h6e3SxSDL8nMmsIrLW54L+QMpVPHSy40yZLHsM6N96U0aFzKOes2HM5zOk0/
KNCt0GVMKqE/GByORhn/lAs2zbZ9/6/LkpXOUz17JFbd84KvetzIE4ObfVtEWucU
vuSNFD6XN7DmPR/bGZxGDTPhMmDn03pjP7rpSIrsQF5IM+y22hnIF0c6V2FGQj8m
XoyhT0YMUc1+vYR4wflvd4SnMh8bwxJJCU4PQwMdG2Uo8tcZn6K3B35BXZmL063Z
pDgP0tItbmWHRae0lTcHkGQmfBYZfabOyaIx6PTazbnWodAVFAw3gCKmf3+6uZs8
0o1wtihUH7trdzcrpmYbPHZ9LLwHGtnlIknJ6mUI9qP4KdWPqclPjMJLPHPT5E99
6OhuRJ7t12mzKF/EqAFjAKr/5Bk/AY6SyABsXfexWlU4xBY/REYH9DzITSn5xxWR
CrfG3mf/aVgEIpyEroh2YUIvY2VUg9qm1feTu4d8P7IHXPND9u6QuOYpGB56qhZo
ZXPnLzFAAULqhtwHrMgnAwXuASGlVO1urMZcBjoTJ77mcYTqtGAxY0pQat8Ur4kg
2gcgDl/BbOFl9NMBNvxOKc0JZ+0onLp4lU/ZyENSGA5GFggt4y+kmrFAaeOGRMMK
Tne6+ImQvPjNVKLpWhRoRVHTeA37wBs7kNWFMpJeJM77nYt3f/wBCsaAD/V/g0rN
+6v3YL0gXwcmGF6ulh2xtAG5l/YHX8aV8lVtD44cd+FI19xATEeLGsY2+oY1Ivmq
gcf1u3s8Wxq1xHT0Es+7IEOlnh8NNlYalyyp4FKr6Elj3K/m42k/iTbxd7zPifcT
XKUIhA6ygBDU0EGGHVcwOr9KDnyeAg5FQglK7SIavN0Da523Mhply9JaVALLL8+V
dPSJneuP07w1XnGNwx/6UKccsixrYp5nOf5nCUw8iYqKWoL7AJGSfr+FdhF2sHHM
O+Zgzo1BTaihuL3/UKqbPe6j5Jv5lZdGMrX8rD2u/eIE/nVVF2QASJ9MnikkoY5p
xIDDx+RhOq9MUNnpsKRjt+fGfaNuIQTHp0QVfNRVZdy/0wf04o6E3Je4LCYxjE82
JvZrVnIQo81h0adAObdOeuhnl8oFwbLKHRk+EzjhXzgywgbN56rrsULG7U8jF7nh
XfVv9yT+LuUfEwhoBAXwvh4KnbLrOEYG/Jx2pZYOY2knegpvTjto82mnLRaEQZ03
cKI6ErfPXNSO1R2D+THLd9pJLmlkysvcLIYeQY7EQidcbEgVT1hz03LhwxP9PfRl
h6J09CJC1QZWQgMdMjZxueQibemQywQ2KE3NcBsSScqolzU4GpBSp5UhplLzzN9y
aijhYAlG7jelrMmbRXR87sCyWTaqE4GXny9KkfUIw05UWHoelJM+H7r9wtKjOM+p
OkLwlBokRWVQaAWTqOGWZ6MFv+uIDtXB5sF7kMa7ssBVfjPxm4l31/3czxF0w7s1
EaDldpnBJDSBDi4sVv7qfw+akJOJ7X29LMMkuYMuwTusZjAqGDVxeXhgUX0VG2jr
GcsYZ8dL5bhbCZsX02ahkvCw2R4aYM6FzGo6GTspK+ZMQkZ52nn20qTz96gJMxVt
cFf0YxFdpfD51g2waYA0HOAws/M3fVtIxQIPVtkzFkPs+J4BLFFK3g27zfJVVTS2
ugAXPQwL913GDIOSNgKvvnrkL7quOCwWTQO2lrZ6/sVfbSnhsP60estJlycYQNwx
11yKQLUOs/5ksYWZoY3rWYlcIi/D4ylaG4nNLHda8b8frfJAFQ4x8y/qArCbYhwq
BQje2r1/cyu8NJYWoequ3RyLu9Q6pp9E8Oj0SOJdOO5PEooSXM0jcqU3deRU6H95
oGhZgN9zW6Zpj5M0WNlqwdnMFX78lAf+oTi/q5a8Vq5mRlL6AYcGcsZ2mHooB8TM
dvqIVUF/L5Wieobc7rzjfj+MlciZtICYJbApbtfW7OiNoEK7tFtzLsXdCjVQmunY
BUhGEAA9DGxWasQ+VDfXOTQV/SnnaeUFO2/J29JN1LSMBHGhOvTNPAW/Bh8k7pFJ
5w3bqZEr4RJ7dZllZvy2o8b+Hs5SAOM0i55qkQl9gtXz/wMBgW37cnulR0NFpgpw
6Q616HkhfzzpmkiktC5migRH2y9oqzsqxYz7y4iX5k5AwHq6cWiULHR+ppiIA5p/
4UrE/5t7PULYdnA8NZoBx40dmE4JlpUBntXorrC5CVljqKJtbMbhXkP+oKHP0C8b
ejkwie3i80QNpnrT53fizgbqgn4qDJZrICab2KpdyWR0tD3V/Zj1MKoMua4LMRGi
iD5LqIKRv7dsS+L/pY6Bb9E7GR5gulnQM/3SiG8g2so1c31PTyUciLcCwg0o2qGb
6EFXZW5OOIPbFYF7lnRSWtT7Pr18lDuVGMO4Se9FIfJrmJgpAlzsBNFgyVt1S0yc
l6DzNRJ/tqsvCu6+kmSzShTCVHWS4dDXx7Chuj9lRO1tiZLoN60gjggULEezrHbD
rTkAvm3Yow2jsYi3oe/yorvTzPDE5Con23ql8pko6tMLF1f0FfeAZJT14hyvkcRt
aTxs7s1Cx0CN/yGeiGGzmi8fbOKhP6ztYnLRPHh4CmfcAWHAyzJqsP9rco1us7MB
ePUx+petIBiOZQXRkSJq2ceYmApdSWVKmThOXLXi1DCQ8q/nWgogXYyoGDAXlfci
Sv6aetr8rXTm6Idoi2jCQP4zACRTgBpINpRy9dBwKAhqEFw7oPBrnA5KgHaawWk+
QNx2Mmjb0vxa5hRjOWDLkPbubA2UcXeNLpzl8JBSiqJm2w6X9WrDF0ipIKlSRO8t
zxSWVH5Kwac2pNOIPLyss2F/n+Xe5/C4JN3yEIZLIabTNgDBvhp56vAOh7+bw7vL
NB4BJRryCCSEkQQG/j82nRzQxZM0KlIhptoqfM8H62s5UQOddf+3MtGSw+X4pSdu
cuLWjQnSbEZD7snN5gqRedj5y2qrq465LBgr1RVXZxJAkkrWK1C70wykJxmceO4z
buLRfriVAKAbXuI9/JsWB1YhTvLIu86hslBIZzkYcvgMrZup7e6Xkiza4ade8guM
cC+/mRCJfm+0UkphKavpzX6ZGgazT4Fkx+nuv4zzUoNH1kryK+8b4d0BB67bsegU
UwVEBoTQKG07o+EJSZXFVyw/Y6LwRL51tUYq4awVMs1SyQjIhABv8zhm3kQJ/fvs
SmQLV8Mx7i0vVQ47F8bE15D7dfBLykU44Bj9Jdk9k2Z1Loum9OPZbMTt2XQvET75
VbMLVwsQu6NEtbmW3LqRzaKl3r4L5AhlbVLHIARii4sUdohdPGt6qBkTpNJ6BWmw
3OkE3ShZVmx15nwHEeTZqre+Y/TMQQ8CpXJelHOoqXuh4Mbqoddah6LvljsbC2Tr
YwH9gM7Qacc7gcFZte5/Oh4L4r1oUXf9Z15iy5KHmyo8S0+e2PHTK24oEfU29vh0
V8Ew+6JvYQRfoaMqdFNsUBJ9mfZrVOZgH55visYKGkF7/Mr0KDgFkYbF9yeNO5uY
chInGUjHAX4IpByZWhFLXakLvfrUdD3Nvmwk27xrt3r2t2zai0vn+6RbByEoKXKK
j8CJqQek+OTJd4hfVPkrk8x7pTORVrOkghEowIH1kaoGPjnFQEKKgSnV4h2pRvRR
clQDwtqXZqIHgaR8rWkd/ELH6SkLp2FpuF6ySKhkNqlWGxqhG7rJ12Pn3K+HCb7n
u47zdPQPvHnQFY5vQ5bLbiY0AV39oQ9IRRSSaMvRfZxbDWc+Rdg//lMJDXgPegYM
IbN4ST+VqMizkUpLZzmZOZ0bRor37Ry60kdmN5E15/Djg1TKnMIblm0LtEya4T3x
MZFwvqGE49+ipcDWvrIlZNdbn9/PiG3RCFnw1Uflh0ROlJfBjGQwSG74Eds91Ddw
nyZBxirVox/dcfpqmQIqUBF9O4JJomRTY/p14dqu1A+dXHvHJVE09lzSyfk3h41a
nr4JWuUWBuPgYOmR9bl8CfiwKqPfWe/jwsbSRfpQHSQpkUd/J18apbM6ZsTYONYr
yNVUyzBOwZ9UW3T/6yZcge8qkT0twWD90DQTwxui+xdp61LEOLBWbSmGxhoGf8/H
/df0vrbuD+wgsX2uHkcOLIYmiJEYW4fB6ZUP96Fqady4vHL0B3CsYkjt9UqxJ9L2
IKxyCj6VRoY65lHMufEQngRyJvEW9h7MeCYQvdns/+NY5Qw4rIYNN/pOuJYAqPiw
Vi/ZPM7ix/BGZJ+JvwpHgn2oebTh9Uzv6EippOrsIWaR5Wn4fAMY7JAbelMKQqYA
OvQOBcaIGjxhC0Jk1LbdBM1r6yNB3w9KclLZBlALeQSmHuSnZ/dw/zitNHTlCwqE
kP3JCgES0NTyltolAyogI/4Pwvi9GiPuzUVKqGiBDeyWovCwoklmly8qBIqmSDYm
Spi7IF6rin1xnc53m/Qv6oTrDeSGvFt/NHIxuStnLi1RccEdBzaS6YE4uxqSiwK/
xoSpSBbeBUIt+2fEbHpGHHPj8jdGZoIwlmzKzn3puUY8SiKJbeLNMffqGXgv2drW
+o6Zw/BL+yXsbfzTlwuOI+VAs7sx668zCX+8MuAVy18ON8KP5glZzUvzb62MyKAJ
y0HIraUGC3O6mpU78RtjHYBqrS8Th/APM8XMfPFYogyee2z0b9358Ymd3g4ikaGs
MfjktW1StVspMp8Y+9h5WBAASdVfG4j1GSbQIaHdY9VM/2RzXVpqRsHjTlj5Uame
Q4/a6II5a3k9aNyXPsvnR1QmzecD9CATtESMHz2XrRyrkWLYcdaq8Fq0CgTugZ+Z
6aeljtcxKAbhZq7P+L7zpTGrDadyqSJhWLtS81NrVaxQmavVhjMU3dFMJsmNm0uO
nEMzUJNCG90efXaLiI1f5sMA+xr+Igj6fdl0u6KZlyN3fG3prz/1CCErQfRhGoss
tfT9vh5Xq7xKbpK1AcvoNa29voUlmzOVi5qGTymzerWPQLaEpP+tjBjdQKbtMFoN
6Jr7FgPrAOBb2RWAxfZPvBnihOuUlbklSVsmSsSk50t53zaIvwkRWAy0/YyC49vV
JuabIiyP5skSbzAtciOjN6OIZzxLVyZ/ypH7+9i6tMl6/H+L1hvZUqmECrEWqwi6
tOjuZ92ocDNezs0dT6I4WB7JqcRtib75NddnRY69mbwRMjkirLHOD/QUKeJXyQkD
kQrgVCSAyoROviemi5BsyZvi2NoXxT/Q/O6sVs91IaVLxLdCBgWlCrgHz2nHNOL0
Nj2pYjAw8XZl1f2L6D7t2QjKKXQDp5cunRsMI7mpAi4R/C1zlgh++LL4GlDrXgs0
+8FlnrVb7bas78DyAtsf334hdWVyzEALUdKMK9lp7Atk5kkK0xd3CU0SFp6Fppu0
taw7KNyTRl4HoJHAZ9esk2big++AkysJAXO+xqkDjvrvG/Jm2wrH4/u4Wdk1GdKB
vSw7dPGlrqZzIreDsOppMUPhK2hZpckLjkcBEh7k797THTtlQzuGqqX8ZLdeln3r
fj/JUc9W7265phVWpzS5M6fPcJUmCQASOhz1wQVI9oDuh4HgNuJpBdDKB7bOW1wZ
Lei3bNjr9fKEV5MZ64Sau1SF0pl3aYjUSuLmP2HMc9gvbruwc6TXqvtIkINXb/0W
i4fA4n2piTUXH8G1rmPYB0JiCaDyLpm5/4XOyuDeknROgZnSMwwicL8ePgJG1omP
ZvlO0k1JhXFdnGNa8P9GvebPG2XXqWmg7llcEH5IOekYPf47blsEq5mF47jgTezq
J3Q1KGJbNb7j/7amQmIChj27ajsApa+gGCY2xK+QuQ09jqz49Rw7PvuJsnM7jt4H
OKfoXq3VYM32nlOGQ7CxKaSzJVjys8mRaPMSM9DyXjXioHVepPjHP2OP3wiQQyqL
+JFc9RiWJcvgWwp1hFR5445hSIHJ+Zo2WRrVjMuY5usf0dLZoNq/7ILW9d6VPT4E
gUop3KOcy91Fouz9JpbvTvdnXA0siQrjvPUYU1kVst6wxl48Rs6WHn7Cpe0w/Qwl
2OoE8xl8BEsO+ZfmyJy3alkFKUIt407MNSrnWuj2w93hWgq28w8kXTmkrMHGwhGG
pNsod4cP8cpRfxrvgs4tZLCpAtPopsqX2kt72a68C/5gDBa7UpE7KBBDl+4ziq14
giJXLOwxT3ap9qSKXN3IktgCu7x0V3AwRiWLWKQz/PbQviOevlGTxKWbvOuakOhw
lANBU5oBkdQI2JrCw5S+zq89EBaFergTNW2j7atp0+QGn5968zFKZQ23+Vd19q7w
Iov/SFRH0hmMBtZSoCFVF1j3tzqzrHztuF+3uNLo9JYrFRIAnHlD7JAHERTwWqHH
kIshj6hp1sDEJ+F53jtTGW1mSCijxQkTvbjlPv+yI48HlCX+OI/V/naki6SBbjJq
klS6SCfbVecvYPZ8/S4ayQCp/3+OtCDquZZ0NT53o5FskdfgZv2UnTwyc3IcWB+t
4eAB+gmDbOSEa73fNEzyHxiXPSXDPUkM1Jwi8q0b+oQZpztDRuy7J4+34uq+Mbd7
YdURtifVgABzJsAmirzU2tdFJFWXLVySDJQh8JAAAXEAcE7pXxvAMQpQWaTynYmm
P5tYdCQs6KDzL3Ov7hI0rmZFZBqF2k+4NJsM8CMWBFb9patDReIal3C4ksU4VQzR
jgsii+s/S/6Ni4G1YDyqgRxXkIlO0Se0oZlNhBGFR/KFOABFVshGi/zsvSDbKJBE
v1khkYULtN64DHWSdVmiWzpo6Bv3qUJrzgjsIF9wqW7Zp1gvuUzD2yyNPQAaRvFy
Wo4dgnlaDABhEjA+TYqdPj+eBbo8HDFFJ+OrpSvF/tvZ3fNJbohS1yEvpE2ytvyj
lkDD372LavIpfog+A3kAAVOob6eJCdiY0L73iGTqZ9fuO9RB8kZzGMQb6uwNLNO3
KD1gNGyle1aUJMgH2OF8UMmP3NrdigKWexCGQn8Fnt01Z66p0rKUJEAM4IrNt/zm
UKpY/qQlJYbNkQa8fkuu4YGL8YvBDDlwqTSzzrjDl42FMDbnE2IkNm0smWBEmJ8s
mhTwPKkXtQtAhHT/RlabKLJCKXuZN3tNM5NRUlYlNvcSjaol6RWPbdCWExI9nP8Q
7Hho15QyALjjF4R1hzuH7OybVb+x8qEcmoOoYBwLt7k3i3Ug99UQlDC6HNiRt9/1
BumeBDt/tljhATYzU3uES8CbqLYs+tiDjld0XOZbQW07AUR+8H1bEHMK6wYPiZ3E
RUCRqKkzBb2dx4dcbfmfkNLIlvTgew6Y4lQQf9SfyMeJlM1z9S1TWq6KXbZD6KE1
hsCI1DBOw2iqFGlgqKM1N5nCS28QHZXZvGELDclPyocusyPuJgb+BeZLUHqS83Ui
TiUbb+ONpBp24MnScGjd9V1MAf3GR4L9/TEymLtvCt8vK7w13HQX7YSnaWpXUoUj
xiEB8WMa3A46gVn8k62EhaDN9c+4nTvhSN7GNrqy94amb+g85StHd4dgzyaOLBbY
JyfxVnf4UEh3bLv6q2uydmv+dCAkKxV1vRDQcBn2BPW+ZzJ3cbdcBaF+rSfm/gmK
BgTtSsAwj6JwPbOWtvI5SO4qMA6ofDwuLgvKO5dzkKHORoF2pfenSNh/bw3+X9jr
AeIyruWlAsR3k4tJj+aaOsVj9GqPW6H4Ut2yTutq5JAuobt5iCcifsI1/NQnGXj/
uAULMGzNnT7VkuP5wvk1XAiKcmXfd+mt6uee2Kegc+71U+kxfgjs1XctqMgQEExX
etu4KiY6oSOLpO6vAM/5zhCu7BNeKinP6Vf0rhDVcOZjamAoi112M6ot3vAbTiMY
/zwbQG3J/kXMM7tJfUh3O9AX7aV4idt+xHVZtOZ39GB3OszhXeK9NQSTk54SM9IQ
kxjyU0K3OIcZfZvVp1xDccpNAfdUsgS9bh2wKb3X2OcV9lYVENpG4wF+i38a9fo0
a1zZEE9FG71VI58e2dmVv/Kpj8O5Vkq3Hkg+mCWgLIIsGmp7KDqzPX7Y9q/aW6yZ
iq+eDUASsjBLJoRCf0zg+1zZRahtTlgVc0Xk6dWikrUT9uR2d09A3lxvWxeO0hma
Oj/4gVAxTAE/5bNA9L1rlSIS7a4nE0CdSATafGgKj7hjod/fw5xesNXNSevWiIoV
XQ5P2PCTgVj/7EgCqeR/lMy+Gj/pNOzsITIy+wvw0C977eJzVC5tr8+6GA5ISxYX
67Cf/bqixysYM/zzInpoA1gSj9h50SXGCOpnjdWOtriEtDYpL8d47QhkKUPWbPvM
1Ezfp9GVACYS9zyPhbiveiV3a/P0henjgQkwBkf2/7RaSMJ/ppbTYukpGMYyVmS6
jpV8mATFA4wxWqsk2YhXPjDfmCQOPrDaFysGVexnQATPQMLsXUVOvKIv9d6CvTQX
rITlfkdfyTXO8W4w5hylmmCj0RCr+RZN2os3cprFhUcvzZGFxexl+G1rqYfz14eF
22jM0hSIGNbIXzg08RtG6N6BxhEaL5rIPgD1UpuNCexcdBH4VgUZTf5JrMD12lwq
OnWdDQ4UDXua+xCpyROWxi/wLEZLFX8dsDd5LXwBzVaQpOqDyI7AoYigNnsztkQ5
Te3fFDpzbWi4uWAlOpa33YQLj4O4VD4/gSZY1FR8VRNXdG3wZjE4wkO1YvkjH6ku
BGyLak9xv2n/c7hJ0fJw2CS3u3bxri9f2AZq5cy1+LKTvnGkxsgk2cCuBmljvu4t
pJJ8cUZGlKy0MnP1JdbRQUJ9ximP/nbMIEz+ZRM6HPLqEw2YAYdNKOLBN/N05jE0
d9rLmnd7G5Ks6dkHgDRpLFNIOuW1vHSRfB4KcK/QaiQUghvpW1ZqIlT45MNToTgw
pm7sDNSC7tg1z+lOArO8nRB3ryoPvRFGWp272Dn7gd1WiKgYpGHzD3cHNhJFgmg7
wfQBZ16cTWmD82NGdWkMvDJ1ZbzFpuTNCgMJvurgNHTQnSgnMWqTFVhvO1xJTgFb
VsH+yla67hMCvphWfVIz3sC9ca2l4zE61/Hy0cIkqUjirFUFntS+zTVWFYPdx25R
2Di3eetkBSYZigs4KKn0fk3T3g81bxclLfgvth9wgLaStNb5+UZ57kHdi/9/6dCj
rha2CC1uwAMEHNNjG5aQjkMBP8FjmkxXognv3C3sBng6R92qnJYgNgostzoda3Nk
Qnu9HUnbwn4S6BAhjCuC7jvQwhUOrbt+YlNtjD+wmTuCgmg4ngpAIdWWUKLRUmuB
F81DSaugur8tLQcHXpaoO23WfLDZYg1GStIsyVvfceKUDa+41c405Z6cWqgDzNHX
TmDe+L0lunp3F3YcJs/BIHzihkYZY1uO0ImXQANb8Z5y7pc0UG8a5P7+0Z6LLYX2
6RgR+2t8HYzOAwM9XkV2zMhYY/Ils0aK9t05fArI2LkEyZi3/e90vvXvpjKBA34X
A9T9HtEwkC2EjkUp7BZeuGd5rYcQkVRxXWY58eZH/FqvhQHTUsmxix50J80sYqAv
pZW8m06DxXF1O721zgOzE4dDC6btcp5jJWNfqriwZAvd5/U61b0fS7Ndg9xZmhB4
eQfrVXsYMZIqdbjqibe52uy1jfuge3dcKDKFo+C7xMLt+6Zjl/ixaXFS/tZBvNMH
7o2nE7JQTKw1JofD5QzrH7Pp55L0Zf/E0A2WjV3qyheKVZNpae0zxl3/e5k/1uSE
WMmN7RrV9Uz5qeu4EuNuezm9J9/kH5+F6jZnE4ie3WNyHqcz43bjz3/MfiGfZjsc
Twmx9Qr9EXRDinOwExxRQL78n2+zV//PJPosGO+d1NO0ifJ0CyAf/jYacI+6svwy
TFdEXG9CIj0F6jVI1q4f1kVaG2jtF5OyDs+WRSRRkl05jnWYi3xXyE/scXufpdNm
/J8uFWNe3UAbt543WA6tT7LPjDFZVI4p8UXuf3ez0vfriRThWLMz3xQWhwG8gSVO
BnLwqsnMzFgxGfOX2ClCK9dYm3nYNkBaNYEiNurjuCoKocyA2iEteeA4aUuNkiEZ
PveNVyzuUwjQIRt1+SHF9ju8Y/2rOQnP/PcaTl+pp6+NUMA0aEkFRbFvO35v2G0c
rdmVsyCAj20qXXzHXzk598Jo4MciyoUNG2xj/PpTv9LghspyZZoNrybgakz86QX4
bKtnlKVbW3huTUQYUiAUHdO2KXh1omeG9QesV6/s6RLLhwHRrFNW+VF4JtxMwZD/
N+UOVk9pHL2CmuL+GlFsSYrlP7Hsoxuoa0XEvWTjnL3ucNWc/6OMY04PgD/luJCP
r4MTBaFNG2ARv7jIMdD0lD43ZutiZbYOGpwUIgY53Xhs+Etc/XQEOb8tcy+DPb8g
pxIjaEYu/tvKS2WfoGnyA8fQ3S4G7VQPOEAqbRqw2z+Vtph4CXOl9ip+3dLtzl/8
uh30C6ZPJsv69ko+AEfjE+fXm/dRNlgEakjk3LEZ8nbSadJc4shcPVlK7RGr6WCp
IHJ31PbeQLMe9ImCZFobnrAaSB7cYDuIFx1r+c7NE5+J+XT9ujdznSb8IhZO3xha
rl3Saab6G6c7bvLj8A0KQUE62CpFxfXexVb3QxWZ2tlS8jj9i2ZSmVxW+HNnTVkv
coIWEqZb0SQQT0ajhW72axxUqNywMOYHceecK5xNJMZAP0ItmoD0BCFEyIpqJQwf
6B1ptTdtjknuYN/U1o8B+U27JCiaihhI+cc7uDRWBSN8wNfS0L3CFcebW8FSq/07
LSy7SuPs+/nx6AKAIRrfe/95IS1EREKtKm6aoj3UIpufHtH7qRaD+ozkW0nV6AqB
g5A38ePbx9KUBZ+eugZXutY7gvPrsXLODulh9wnFu3d5LPzwcAGbuCz9NUszsh+/
vNidPdIMZlwnEKF25mTds8i0wstOHJcm7avXdV3zz8UodZmZYKAHK88HSF616kye
YqEACoxS/K8viMtu0aWwxtMa1NwEcMEUla3k1rkaw22DQe2T1Sbt9u+Y7mm9E3jq
1yszNv1NCAbe1P5i4z6usjhHFpJCVVZTSzJ9VO7+lYF10zvmrHBeF1dzPpGDKUL+
N2GNE2bo+MKUHeHVUMBXM+0S26Y46pu2i3CkRy7085T7OidZg4GQUVgD01PjILnI
0MiKVCGi3bHem6mhMkU+SZkZ9a9X7vAbCQyyqwB99vd8/U7mIkwVA46zSBBdjtur
qUDF9Yd3/hSLCOE/wgC1APjZFpcBojzmO1CLQEB5ToHRQNd3WqrrwDyACV1veFnH
GAu4ZEIvONZ6Bj8eZ/3Eo+IzRQOPdOAiTbe6PmUhSAo92e73tcRT2mXfsCt+lB9O
rZNOTszrNO6WGKOWnAxaJP7Wb55iC1jQq3I1h7X73XQiX3FLJRJcZO8J1QmGZNdd
3qb+DgZiLlVU1ST+8XtbMVREqCe9Gwxql0uFLZg+b+xYvBD1hwntuBYSvdsokE21
XHR8QHnVlVlYutQtct54IUJi7LmmfCPFKse2gxsQy/zUPlBu4UUqZ5zqAM9fNpbv
AIQXpU+TR5uVzqxJHVv6+KPCXscUP6Qop73OJdbO53TOpz8yJYrWjNoFefkQiv7K
btKE3X+0gnIxHxQ9yyShwTzJj4eNE/YJyxsojeUmtboKA7UcIdcvBT+WdzPL5BZD
QTqkflWl/sAL/FAHdnufLcYAnjEcPRajABZPMRfmf+6pMVvJx6W1SJjB0S1PWKHS
o7UxBHT4nz1LndEFLbHS9RPZpB7p6s96Az0qPxfEkY26711ImKHU9YGamOpJRsuc
rX/VFckTd4YkIXI1YBIbojOXfyU2bE5kdxPqCzFA/Hj6WpBXKZFrbgqoKG1Ra0EK
pAPIi7xTFLYEqS5eVCGnuZIuyecpoq/d/NbHiDH4TdvL8cpcPSW9lt/CmrYnx9RD
sjrnmpcIo/58zqKGH5SPd6zZ+gjZgXmHIYMfFnC2LQ4S8WCd6PPOFo2R7LuucaH8
JEUQJm6ht6UI3Fk3z2dkyQCTmYUB51ryCK1URkSAIJKioVmWg2JL2t6k+v4jWdu7
ggYGX4fX3XH3RiNZOWpl5w+iI8D7vyvhXbH88ZNmn8/guu8guVRWhq2BR4G/ZLTY
9aWhQTjCqHAnGmnKSDQtlecITDaH+fNhX+98nAVckmG8Sul1CvsJu6MF1VAirKZO
kJp3SpaU1m63W5ODeV4cY6eKTP6qezWR8ZsmyOyEIddUmkwM87GqudH48WA07XmU
TgeVd71RVPAbdZkinTAjpxhBx9ofmnSrw3SkECO/KgwBeNUhcF9apGrhbwEWL5Gz
2iCMAAMg9R997aIlk5p26pp5kStDBjf5vH+s3ZKOeYd9zYgrGU5sfjh/z2uvJeuw
eOmpXAL+XMnVUPsxiflKfhd/lCrncV1a1kRF9wdtkhuiDXIW4h+eq2b9dAq/4lme
qoW1/zre7yjb0MLA57P0yyB5ufDecC68fDq0Q6YvlG+TLu7+2sArRHMhfLS9R8Dw
g9uZmCO1vXk5GdQEATScSt4RbcZ9C+EnWHr8sc0ULywySYpqj4O6iiXVYpb/klS9
fEku01MSin7QorSvw2ybQ5Y4blQePCpvHBj2mUpeDpza3aYKLtBPF2EQXbpjqptZ
DAQcmvSyJKCGxCmlSi/wkgoRPgeMX0sP1ps2eRosQEBbnQsNiO4skxCbkVljkxsH
UErtHAwR5+u8uJYLxku2nz92nunxy5J6SM7135OLtXFTpGKA9ou7acdbbc2n/aR5
y/18p3y/Ax8icgCKPEk1vJMYG6WgzO+bItS7f/5FxlfHJaVE8vOjK0ZZs94t4XqL
6vyEbY+FmI+YJc4XW5UOE6S/w5R/xIHP1zAoioTvk/dvi+SfhZczC8XtBcQK7a5L
7EpEShaetBP+19/gy0okB9UwW5hmifJOcxvBvL/nmFrSb7UIWlLElogWelpfmvIe
bbIG9p2u+PEZKomqwFvKf5bnkbFKaN9NCC3yHNilHPQ7h1wfnyH3KOjbR85BUExn
Z+Pofp2yP3Z7qi9aQdk93JgQ/U3/bVCHlSRvNXWPZ3Rfqtnv/yHxh8Ui9Jwx17n/
OAAT2+0MJRwXJT5KD1vZ07E1SdBJ8yq4GMrwEQvpORbu0Qq/2QSZ7XM31Qscn/V3
jgl4zlrv3Vp7uYAlj84myyMFRGHrfMeNSEdqmAzu5jIdxpShJfvavHVXmiW6lFAI
M1isw8VNz0psZv5XQ2F3R2kWgpgUl7UcKXqKGKGBE+V72QQHHY5aIaWvvZaXZAie
C4AjhFnj29l+yacrITKF9hjaCGERci4Ko1wvco5vBxSsavOSDbqWhTXZmsjninMc
jrRoxlUowzeRaRc2CFlMoZk1R9mLnsnM/lm5DeaA1JMJc8OIAhOu7NfWVbyY/MEA
Cle3vNtChKfyDirA2UJ79ZhEqlzCdDOzmA2RFzBYZrzO1o025z3+MMr0TFdKyCq0
VkZOBngNKLfQnVyqu8A3RxHnSKuUXND+9mrsMKhklMnrHAPvjbdo/Va1hwoM6agX
+rSfqF5p+FzDTfM4WdwXeXER4HeTJAWMLf8ieR3wRFNWKrIEIHQue12TRucLBZrM
LKTrkqn6Y7b/KflDazChm/gxdTt5gC0GqPHUG5o5pInnVT7V3RB6cfrPrMznTlrx
9Y9BSADON2MU6o3/9Pp8p4OTEqrhq0e/2uPYRqteZ5+A/CEIpDSkofX47wMn8P1t
oyU1liHeP6CApcT2n8CBd5hZAdz1ubzfjOHYLMJYXgeFqURMHgNI7pXMlcS/c3l5
vO/Plql0u+/0vqrkYDtCNisZVRWCUo7wNry2+EYTssDK+bjYxOJ3WUou0J4GXG3i
RUyNn1RDTIQeGdaxCzJ1SGYFOBt55xmN3S/h7JNDtoNnMKc/wZ1/NeZLqatBSwaS
h2CJDB5ELTw+xYZSXPwzoNqpqvSpK7IH8hf4eQXLyJOLKAKB8SyNPn6arazcckN9
kY9Z4huoHVC5mBx8NVIrFF7QbNvGy1TjrD/juC0g03kJ/D1rNR6oHM6ghUlDv5tQ
mVMuCgYtryyakizCXu1/+zODphVhcnxHF4HSwT4xpVC5+7QYnQl48XSErOiNjJbS
cwf5TSlBeaEweu+Mzebn7g5IUeR2nGwo9DXnxux8OBj8JU2GYusdJWDID5nGbN7Y
Wu/lpHZXo77yA81cCXWdzZIfK6WgaXDP6Gqn1NxYhgS5FyGs/B2KIuqYI/8ETzRt
UvbFYdesZid8UokMOV7IQ0S2XTz4zeVJxe6/Wy14a1bTQGTKiSqyH54N4lP2yOs9
W6b3jt4Lkjvd99ixDt0ajskrfn7XNvwkDLuZaWjqYVIK19hJkQMyimkyIIcaUk/Q
CAP3bba+b40c8LVA4PVHnPH4ekd8fIv9VXlfrmDd2RMC/xr8bxFmYvKSo+UadxWf
78OXCGPSlO4PlKr/9QSi/2RUO1XQvRRNB6YfQiMjWXeRci3cC2IMP6M+q9azj9aB
ksyVQMJHB4HM6ydVM6nImihpTa2wUcXzSI88bTFWpOO+U3+Yk3U8qk99+ymkOPke
sQjSbStBemZ7f03VdBu+hNOwA5OfiHAqmMJbjgXlChUvVR2YxVAab9YmiHgDAE2X
V9H42Gt2BGxiFqKzS3tpZ0Go429jwWOp2dDWrauXkN4eXZ8WN5vxWRTAeg+5pe9x
rMNVWQ7aDqQgChYEDHehwTv7HKqBusZ9JBw7UaoyyxVSSyOR6cHKyW++4fijlI0b
5Yfi029YVoDCkZ45KcxF/wJA5D2C+KfWxl3MYrig05q1bM0QkrRqH8iL09K6X7jR
y5/JaICzfCLGdS45c3NGLqddnHqtm6DwwIJc1dIOG4HmU3lRjLL7CPfuD+EgHFa/
o0yYWuQ4xUYpTa9kM5e1DyHQA8fCk3Eq4A6ygqRu9ZjwX9aKx6Fpv6AlsalG4uLy
1duGPti+5ZArvqV8U6aKFKJ2UMmMzhgSbbQyJFy1JuDDqwzKz11vnWSa0YT2UrJL
Na2yncbWKP/TPVVatxZ/CJdGqTftIXN/uILSOj6FTfRtPehN74+szjFFVb6x3MTe
Kl1LUpFpNgOtJFx9Rc3r0/qCjPk1ER0B2Y+uT6ZIKVgpVEx/8CU9JbPUW9K+vGel
bE5DmCCPvsrg5tYlndqadqR79muZfvyEFIXE72xV5z8yayfCrff6lCzC/WOrg0EN
QHTvf3MC4ocmCYO0uU66PXuzNyd5mjc1ebT7ttFzWOL7JjYT8xOt5nF9+GJvfzmB
yPFbzB2uOg+wjRagAu3dYZ1Dy9ECma+jiKER9DBdLQaaCgk8sjsC+udfdcy18dpd
bK9Bov2snAHeOSCm8iACTzcg88/LFOHr/Nf52rB4egiJimAFUpYAwoEAlFTVjhw3
vi1bMCYhKkD2tgCxI34Hyh/PNXND6xI72EWRJPh6bzETIRy8visye/m1C9rCDPLN
c7ty8xbEMro+w04S2CHgHwtyiuR3r2dW3RfkWBsR6cEvUPp9GEwa7ysQTdFcuzwm
d+qHf37DCBCA4QGFvm5Tk+uTlJhBbl2q5JIrmk6BQ3q9jAmyqleyUnNgDKefCwXD
6TKZ9VlOQXeYCbtq7w7h5FoBlwIiteICMwWRoHN//n3eKV5GDClEsI7i3iqXvps8
tm/l0dBFa5U6IbYrlrudzeVBzocXO+9X2l0LqlCfPNeL+24Dk5fCgg4zP2YGoA46
9wTVfhnBkFSi0XOMtaTj//qbSdSde+ZW8FOyqxCYvijsjt/jMSN/afLbX2JR+PRM
eWsMHOROYgUx0D4Go8S26S5ldR8aK6Gw/lvL6P57XVYWRbAiDp47ydqN4bpclEUM
mH/5FBqzjEz6qXJSTSOlzC8YTYOJPATsbTqpqX7b084ItIo0yapX8Q+6JQqVTyW8
aKd0KFcNcpEEjI1Cto2npKVHBC51OYrH7O4ANUpfEevFSL20FXuQBk4O2+CjutAW
i7mbDXh0ZGemIcX/X03VJcZMdBdiknQ6NGPIBzJrPewtSKVv5AY68UdbInPIlyY6
4Wn+xR8UXBd6b6S0YIhzNPuhF3MST4J3tejxTqbg+o/M2iusq/JID5MU/gzZ0lgc
sSuWLIaIqu2gQVlQYZU6Id9zvrfuLN4kW/l3iMapcTMl4i1IBqnzT2801Arjl/7Z
kQGF2khiWrj9W+y2lJrtV8pFs0cqKi/e3kQhdrTPitYJx1mBwR6ahfEQXUfhAqhs
gFKgXzO60spbGWatVpXXXQJgw7f9mhShny5z9kIZud8SRhZxRBmotOfGssAlx9RY
JnZBs+7PzX3oFvgb9p65VyX4ca50l4dgtZz3ExEQsq2Q5axLeE9y8CR1OQRaOQe1
b5oU/uKpXGzBbaRIObufQ52RqmsWbqXfjN7x7NbL6hqROPb3vRDe93fA+RVKleRr
ou2FoIOQAKUy8tJBS9KhTrTfxVYCDhyc5w1tiV2oS9RCiPE3XIvmakwwxyS5Qviy
TcZFopllXDGkTaqFzDgNPR2HG3UDhOJFOlovkp6yHydzYZmkbw8HYi1XCZ3Ap9ct
lqZ8wnNoQlbGfP//SFqP0uZ+oc+4dF9eD3fpoymzWn+T/Umr2oTgy3JuG5x+MNOn
GWvrQhtuf8+UjvJOCYRF86VtuFxmxDX+czCM3DGsCqmAyLbTJZ/uiObzijNDSNvt
Q9hrhg6XiaN9r+Lp6rBwPkdXa4/sh41vfHxa+UZZXAWaCkf0y2a+j4eViMPs0FI4
6A1K9odyPHSSL41qSZG4paVzpHxvjoesWIvfrCoVV663j+MuvKHPJT+c8c5QMOyY
8v4ui20qTm1RbvgdPRNpT4wr7c5Xwqa7UtONEVRWFrSvfWjWteg9hKltmKrs8DvA
KmHbT2sSrBoA7bkXsVh7smJUQY8b7NJ+gYFNRQodOPBTk51Bqmkdn9lmDOq9J9tN
FPQsktw34+D1EYOblQfxKEk8nADC9NlxXdSvfNTFr+HsLQZIvA3pcXEZkcxTLcHJ
Sx9utdCLa2teuL0Vdzm6yA7copJboqk+8D2smCEBDQt+bx8PMkw7FQMqw2l60G7a
SoDo3Kmwv+97MZ4kLUKCQ/7r35se+fCAnbJNsQfXKfEMl8GhdaNNXxFPuaA+6O+u
ssi9hL5bKlDwHnpu66zwlYZWm8d/7xJ6U5OwBHEZ760gFUm+XTZ2sCR1p7YF7AqZ
ySrAY/t5U8wFZGlNYxLknyoVKm3TTfW3ShyyMRSAmRltFItvUF+6NSNUDMf2ilQH
n85IYsy30EfRwToNxgAaOI8hyJ9ywfMujG2WSl4YEW+nlynTPOM3kZZ0UmM/SIKU
D0BbGFitqTTdlnMuEhdK6kUVyjlQwzq3Xy1q1t6T6JDuCK4oJCOMnyu2AgNiEIXM
JvUZmZXNZrG0hAjMS1ses/mvPIvr1EBhYLZOvxPD/BA8sk67N90ADHTVIxBJGA/3
/uajkGfkFTWZmOWZxGKgYBQuZYBsptyY0v/d7p61EVq88U2K9j+XR41u57gPckyg
ZJxpCe1EbbgVvre9JYlbZZe2/XaNp7T2SpO+pdHo5ysNrX52mnuGXwBQoprMUL8G
/gdSN7w3v+CiB9IUy27DdbhKekBtvD2oivtck8vyNTH4gp3M5gdLoPmSuYAt7//5
Abojdg+0tQ8k2BJkJ+NomwBBPfEwxMrTb3vg/meqbWRGEne54VRfXGlun95MQoY2
3/5IFg2KZDcy8h6cZ393lNSVgqZoziCbcilOruCEcwpz1tL5lMSU+kn10dpWk1Yi
YQjjOo3wZqJ0z+qH+lW0et2EALSTJ7ZwLvZMH5xbPZOG0RbTJr6DNSsG5xmuN6lf
sQAFC+35ecEDbFWcib5rhSOaswNHRqpgO/1CAkkB26S1hnYaVnPSFBITL+KWF7Lq
I1na5zACnUrSw8dL4asI5XRIeQeUFWXY1y2EyIsjpZpq91mSWSdccYzg8XH2+LzU
icMm6pW5GYAe0+0mzQWBu4Lz3o6hIT/b6fV/S7opbVNqw5ZVMX1XBEXbMh58r6Ft
7maFoLnCE+qEbhSWwllsADAk/zNPdpU8jSe7ZeHAyWVePpAebL2OgvzFCR9bUDCE
X2bm0A6CINUc0+Zbac7FhdI5hX+fFbCo5JSGy+txwUEV9ALlfW2FwuGYKDooOogM
5M7cIwS3mJXExQWzR8ltedYmWTZZYRzpQrX4k5/5c22FRahQGsynxb2N9Aroi9cB
pVz+HztpjHyzylzyfkEQFztpJ2MCVOtfwUZSm7/koaWYg3J3uxySDMiKSRU5nAHg
TAPDXT4M/zV0mQpuTs3p7wJcWwl7jy9/PIvpUsqXCsLnxBbfeK1ysysj1Pl68eii
a4HeePba/a0Cbc8fs/CnsQwV739VD6l3zJmLMM17z8VLEYYzRAb2Wo5w+Vr7sYRE
J8bs9pnBrTvAOeZYS3Q1DabVY0A+6MnW5CwuFyAHO6GO0UyrHoQsQQ0Cr82mCqPI
33r1l8OjINK9rYfnDsQ6jFk8czofkGLSxtbAYfGycVy4RTDd8yNxp7bk1HGsBGqP
d9S1GUeB7yYiZ/FSIObfQrsSPFgYqRC9tMCNfuzY077rnk2M0bY6Xbau4mdWYjgy
IhjOQTJtgioxR1Dyz9RYkfdRviwyLyRXjwN7mmwMEWyJxXvkbbJreM39/pDQptWQ
It3kV605xwoF/xX5A1tVzWDIFw3Rq/aO7KPCytvO2I4k7zrbHX4MYjJX4pAXsU94
HiLJ+FFfsVZIn75kMBwwud3cC1ROuIArqf8cAyFawGIw4e5VFOaCKEpD/1S5GeNC
rygafqshzvQYus+M6CoIzzS8jXmXJiva+/TlVN1iFZTm7OSwyZVKjDI7wAGrQek8
iS4YFStBxj0QlI2pihcS97Pe2q7JiWv0EP49lwWAGNr4K6mXSf04DtGOyVMifFKe
Z076Tch5tRklRKoQfUcb9sCQhNggHCh0bp4052GjPz8j71uZ/Ugl74uQBxSA12dw
Qm0Zdi2tLLJ70LA72SruZuBn9lCURchhjtiRf0XnsEJvKEiF/cUF+STPDcKS3aVs
uxRxW6bwrHPC5djh8yBySB1mmfL4j3odlfhPKdj8f2CBucPPaQYdPpYDCRJSiCGj
yDcdXihqsX5WcNBfMGzp8AWzyS7BLbnyp9xT5BgTI8q7TdeWCVDIDGkvTI7sncIm
RnPCMQ+5zdQ64SGlPWmmZYFbvmL8YUKvYoZTsrjSoB5JazzbjrPxvgskgzxza2VP
RfyzNZ3FJ9Lby1OocBtGfosf/ODSDtPhuQZ0PP0RDU/tgtPMdoYa0Zz+vyIQ5VzX
2ZBYgEBs5S6gWgPeg5salZiVzvDNpwGGhjYhr8CWru/BF61qf9qe7cRldvD3n8IJ
Pe6O/YOPpB8QClUkjWG7+i6BAbZ2RjtQYIul3FS4/8VEbEPhA3ynJ7ghy/5wZECs
AWbHY2yL4gDCgmhudwAY87MiVlfTmjeZtnQO7+yYmHCHmIueYk1KuSzpz+2j8TUU
GsY3CV0s2Me9BoVTNN2MT5WomnDocPn4bMeLPMhwdBM2vCKs5UNxZMrtKUMXu2JP
5sgHxrBshTfUReGJHv9C12LJqiwwBV2+3tg8bFzEZZ4A60uL5DBu2OHNV9CIOULY
TdxejHuBitKUMBqgSP+nstn/i3Ocpz3DNE69a7Vc3/j7XVupe/PiTZfG6PqeJns/
GwouE39CUdOcK+7k7K/20AW06YDMY6I5TAQjdoMkX3lw8DntAUbK6VlqFx2yrU0Q
/pM4q/nwcGtt7X7KZQC7YfLtsE95F3FRZBKwmo++fg00qpOgGCs++mOhg9ZP10gX
svlCjSXPvDv4t/XzdHni0svsNIVk4fR4cpNb5fdvfjjwQGzzb1BMJFTGKPJuM7kQ
6EWTG0l+kBDlP0xmvX0GReGrN5Xb4xFFoNpN4bCDX4nWvg2G4XaJmQ9n04J/4z3p
NKQSEXJQBiQDsCkBwaiPmOFqvrrUTG1C+SJUbuy42vdOYR6UkkBXX+PpBVdwklA8
e9Q7Ynq5IqiY7uSm+n+I0hCeCZSspupK8GnBmuZUozbcCmAXTtFhx4lvUOPlCNtI
L0Wpit4nXK9uWR5YNPLT3VsCmrqdUiw0tEahlA7cG/GiiA6Kje90Lf5EqzlQc3Zh
sJR0cOhDz8xZLn0Y5GPd4f8HPg/vUGQjqkgr281mAiG5DjmKmeWhUBPrM2Ycp9wk
6CLgu8TA5IauZYXPOLp18XrDDZFaEjIXQosTCjvUJaIi1mNP9VxrDwRnYX5+BeZ3
XhVWJd99Q2i/f273zgaDZaMIurPkF49PD572X4TP3orD46r2rU3oO9FtVwxe251j
4qCExXa27aDzgaiqoF4kyYk4j1IgqhT7eSOiDKLwYI1rOvLTmKH7Zu8BHznWTlqJ
AgF9tJlA+eLr8U/F25+HWaa9i6zn7uM1oeX0vQfFmno7ez3lHsxsXBFdTuusgLtq
lqwO+J6O4e34xJ1qEQtWshsWil3Lz9aKzrztIp2BupFgMtjf96Kt6ord/+FQEalW
DBP6rJdxqlHKVMj4qUhcLIrbX7k6S9roa1nxnGgXoPbqBVXgb9TeAe13VHZDYBET
phA0kkAtd0nGnx6Nmu0REaNjNA/0Nc+IkS0gdf4HpJL0LVsUNInapVMTCRZpFSAA
BgyR8yayZV1y0k7y8GlmshYWgF/Ci4mmEjt9L01if6JzdvU0Q969WbuJapOF3Sbu
9ySYKsN9qqW9GX9hKsFowvVLNE00LrJFiL3E+qMfIdaORah26No+A88uveftx6Wl
PGyGdLXYXkCm+IJ/rfT6rWkB5jLfkaQZLrjpEkOZZFFsN3LhfwUxEGEoWg0CbLef
V/6Va8dr3Zgiu8Odqei4FmbU7quYL9a/z6xNSSW6FM/SohmRWUe1qz7BXHF2K9rA
9kslqLstqtq8xF3dLF6uUtJCveDEEdU1EsBS6bB7VM8PY7327QkfZ1c0ff5punNc
szsARulSCGC5i800QB8vvAYot7XEEXE6n6raoNWqOE+hOx6xXo5qSF4/Gub+0Xvg
Icjay6MuIFjQT23BhuXlzWjdfLV1Rc/NpOlEmfeBR5L2j8r53hQFJnJo+NLJMOC3
dztao/K18ptmLTGnlWChh5Vdwlz6ZK/5TQSEBJdhNMS6ufeU2qYl8gRW0haYNQVg
eopc26efBerNqkYOHXsYOlytiTm6sUnpctbwCYyKmSbpse+oVg9752wpXMMmp4f/
VIg5EwMiP9c1QrE+W7N+DIPIJdEv8Cxlaji0e4gIQS6Epj0gRyiFbHQIXeXLMH49
nnGgierrEbsuNKgcTsDVGH7Ly9P+sIdPl5kbGPeFB9m2jWqwEytj59YT4x0ll4+b
QL6899PnncRdWFonuagEp7IQYkjhIwrL2CCeSjnWVOEJQtXjAYu1tfOr2hlenr1n
8v+TBwyg8crkJJbocou3AzAH8IUKHcOkK7MW+OZzSdmGiF3KVO14T/yOOV7H31v8
+uxzR3wNigoQd0+zc3tlhbOu9h0/e+iYnkqop7xyaJ4H5/d36vZYHFqe7f71gIqv
wRsjw+prJDanG0AW49tmbVbJif0giRQV4bk85thcEa2TqI/tkKWhqko7kLHQCeFE
c7Zd9bhIvx2cjWcIoms2qjsDPVh9ylKxOUEdI1AvoKQLkAUecuXDB5aOSZjCkM2Y
qLRewK/0J7pawsxhnWVE2w5cviyo5XKatBPEovCWS+l3clMiIn/iO84g8VmMdtte
+Ufy3pdrJDtc1cL4bqa6YLX/RHlPtgiuw27ASlxjinGHdJYvX1tvI5+8QGQUk73b
JbqUa3fk91fPTemsJSppwDoyLNubuftfL0AiltuyBkwnpY2+bDQikdrd8awKdZEl
43AHCoHTVEpNvPgUFt4wCtevDX2MPUIwSJBgX/ihs84B4xX1B57ZdyrY6v4NSaCo
OwE3JQfPXQA7FExMYAabpLRX3wKwW3bkyWbicXq+wCCvl122CUzNI/QBXEQn+fv0
SzHbx4Cak8HXtzNHyHnhCLfmwtY3oXU8OABtOqVSCRnQd8pLX/MRv0trm6BXl+v7
8iCIt8/As42ZhUflxkMtMGewizmtDpLU9DUTGKWkNLAQ0ps/tTkX7YnEazMdaYVR
D1OcoIjz7ikcGARoZcBFlKfBMZGJkq+y52iZ39GUDLwjDxmWrss2CItML/X4qasW
FSUoSrCjNZpg/usICazeL+oOVGZsMh81vDtQLWKfDDvRfZXhsBZaltvIcwq0Y/C2
u03ZIUtXRUPfy+hC9cYqpTGQ8eSEpoNEi3VB2SWc9lERjb5Wh+a5ek4kzn/ohSEI
tJ0mzXfs7BcOqVf5K+FiZM7kUCLP/m6SnIkiysVSZkomTFCLPhaawW40hIFRogDT
sUjGT9yxNihlaXcgXOMVKWdpVeqRjusmXaXAhak3BKsWIET+UEyAPGHyeT0qopo+
hl7PlnLLkl0DA0XFmiLR4KU0kgBPXA5Nx4MBDELDKEupPSO0rb1qc47Vghi8oIsz
pdSNqJuidC8mDrwXqkV/XqcNFcTvkA/GpJE3LfoHNQpp68iXxv8xbZNhfDxjUZO6
IER9UentGO/LwfJ+w1WcLcLhShytcxrjJNktpXWK0jcFJk+EAp9Y0skMxYqqKOMy
Kiv5/uc04y2n7qeRHF0YeP8OQft8SMG7g7xMU09PZjN3EXwYyIxckfB1f7O2Eq7N
ZbygjOYrIzJNVNlY0X/5E2e7xi294JUgoqFbTxUx3hEPyDGiA9IOI2w9r6BBAfus
V8BhWbMgkoBABtQsjny97Y3D13ZRJhg1JfvRdSjs/HnyC/kZhHsSHCForEw+jikd
7MFY5zjjMPRvUmw4lq1bdpyh/rf89zR6K6r3uBzWB2qxBu8FMypE0b7cNy640TVA
XGqxeWSLwmNFWz7isktue+UXGl1QSJM6qvWdu+CVebrutAfqk5I0BmbUUydDivjI
YkPQHu4RXyJyqApvKDpSujubdKzvcpCTbn80T5Ksv64kB+bkrzvAroowqLFuYKyK
NxTmfyUcOJLRfikTrF93h5rOE5RIcr8jC0gLKGLlq9S384zdI/gsfzyJVegiLj8u
21f/WYkuR63tgWzMvyuL6lhc2ZkMvNB54lCAApLjCJBNuv/DldHNJsVlsMTv70Dt
t3gI74RHKmKFD4H8WL+zMZJ3L+tmjQNKsCgIyuMkG8K6phVhxhtbCGrXJnAKz9tk
C5GBTcgIm6LtbfHglpkJtjOLIGoAQR6WN+fS+8AROZnJWJ5zZaBkW1Zl0aDwvsE9
AhZE/LSJiL+t/UE7y1xkTrenuAVC4XPUL/AgATEeBxrpss9NoRi3+tuDPhAM54HP
OEov6btb46aX22kMkc5j30Hq+0KoofbX2HT59tSQ2hcUI1JZVrvhAEENPQoLpV7Q
1T1tdPn2TTSJiVke/OoYRO+mGWN4J4MaAT0wqSFXV+BiZFO5wofon4N9n+I+aApL
Ht92ug1MXIUmQKrFz5q20ouY8LzIb1wIIjij0drLvJwJhbIsMLzH7KHYE2GkXZud
A6v5+QvgAvhR3JO+i1qOqochTGgaCCMH5D0mAQup+VKYDn7975F9nA1gRoGGqe9Y
5y8QBrhRixkpZQ6BlnkHFKMkaCTJYEXc4NqSksf/WLNdNtgFgzggNqUmyOu2fB6C
V4jW7SHYKA9iS0dz4I1Yf52dumqC4pnpGqK6b0C4q7EJ1xpMXxcDWd91imUcGdWN
2/rjjpm5y18shooOnITX9BhieCbI14GMRuN+GgPGT6ldKzPGJTzUSOwnnyo4Co47
9u/EJoW8Q036rcSi/qDItgBsf4dqf2FZpFYwwwKwiynVtEdTdoTxuA3lIALd5Xzt
iQ5+ZXEsk9NEMFApPy2FZ1k/0WV0D0AlOCUqahG6OKk/AjUGbpWMApfVnJNJLJcK
I1KPjXdrCOjrA/uYoy4iD4Tk37Xfe/pLENftJqZzx6GkBOMfLgA6LPyEtAc59OnU
PQXHo3fNirZoghJ/Iougcq0eIeCJTV8mpOftcFwUHDjprGQvyWCTEuuSa7EmsLSF
fOkt4A0tNLczpx/reN7/j35SvkqW9n3YRJ/IAA5Hc8ZP6Do1Ig50wPh7y9JajSeX
5job7GGmymgyqtHOb8SmqVJXcr8dpcIJPQjTVgWFfN176P7w1iQ26NbXM0D8J190
NMNZDNYhd/DluydOR49lRTv4XafAdsZyYY/2dWrIVNN3aZRk735KqKmG8F4U8Z3G
YOgllbHQjU5XW9odfPzyQ/0jGqLALQdAfOole7GxweTCBbvWr5gQU5G7O7zVQK4U
P/KFmKlOOV15hpIsd9R/iSK41aw/UXTMShm+bizJo9tlteY+2vzkRCXJZtV11eWC
QS0iWeCRoRXfERxy0h3vo5lvpxLGlN4a1wFgpH43EtQqmvPfMCVsytcX6WcnIYMQ
mVVfY+Dx45LdnzCXuHnYVjEWfrS+2nq3pPfGflTMMql/QAU10+zgPpBFOty9fq6X
BiUqdhb5D8RdorQ9HNQYNIpvLD5w7UNmrAhvpl/rhDJFh/Y/oB+biwzdjIV/L2vo
MJi7obGifmew4nApW1IgerEaGHhIgRXuVWPEnO08GWvKPMn25Oj55yFEhe+LrtyV
i+t/cmajhnjuioAPCV+WB1iRtsyHO90nwEQowOENUr5B+jsugrNk3FAr9kxXaQiV
2oeAqqDpzxjMd1659dNIPZ4ZCPUB5nDB+ShdgK1/xnZsuj65326kHqq3MwzIyPoP
zax4J0p/zX171aNjrOnv6u2SXD1o5svppPklZHntBsjuRFytLYKHkVNv6yIPOFpi
eZDPbUw9PacOvV54Plp7+R+/VVMNz9XE1+SeMlFYz/dr5MPj44yESj4bi4zJONTy
HcykNugNl7zU39RfskbKKyTpKvdW7PvHZJz29kfKs4FDnVPsH6wWK/GDgYobmgKv
OPTHcIBJCIhKy4L0c9Ww28rqz5keznuhuWAlsSgYv8qgMKZwPs7olJcWA/EI7Tfe
oKXBZ6bstDW07GNxkJmqKbEKj5nSdqOnWiIPAJg9JSj/K+u3VRT9mdp6aF34JBKs
dVsBMvj2k2JHq+0M5wOUZJ0x7WxEws0fLQGYdASsP75us236ciK//R5ZD0W9w0/N
/e+h9rNCH4kSqicHw99Bfiik2bmsQ0Pns72vRtbjdwda6mjFtCTtNowK1PnkTr6L
TkR7gu43nOj+tVL3cVeqcFSb8Uxa6A+5ucpp2irwqPTysVN0Wyo5lCLCSVZOVGSS
GL9W5EQdw7lTTI4nf2vNDvOBKSfHUkmL2ONqqfmJQiRre+FYMx/Zw0PhRziXImG+
T8Nl8TbLK4B3FvJdMtGkIbTIDAoTlbN5MWGJ9S4uTUt3j88umGmf/TrKg45hWj4T
opC071ZlZ6Za10+eocnZZuY+5TJGkP84lqHg59Aiajc5OK0tERhfFG7D2xcjbkGA
w4YanzaviZPCf6SgJYM8lm48JPeNrdcp/b53lYPHeu/Cx2KEcLvBefe0U1OcQQLU
7HI1NXLMCSjnNRUHOY/jHknFBECaYm+knShcvGLnEwr+cVLbPmkqji+EAG6hfZ6D
KQxxZCUEOPQqS21c7+jSCcUJzy09gCl1G/A3py4X86Fd6VtIBT/nWiitb4YCtpIT
siCssJuEmVd18qHebNYooeQbqH2QJ9dB8sg12wHqWCgom22jZXnHcy68sWNCqVDp
0sQGaXpkA+I96wbD64UcpDU1rG9MIhhVknoDX7lAVgWB8C2VlWk61yXKvs6a64YR
nQIlr/lmbfj1Qbb3vN+1cEPHQBcbuL/owHmeMsS2b7cWC2WUNr3I1qG4vjQKH60Y
LdKyPYBBH28ywdV3fNKeg7Fzi4TVbNp7li2xgGK29U8dYACDQe+87m8pmls/wYMm
Ku5o/caQVgqN27E5f2ZHfCAJEV7QSj+iDicKI/xWzTQI6fGGjSOvZufg3Rwzh0OU
/PEJqCYZPA3qXj3qRsPwZKvpEVMZiXy+M1517R/rqedz39dBatHxF37AeaBXYFPY
soLjqhfvgTEHe9sYjNc47Ich4JezGs6T8byH7LTcGze+VRn7b8wxZ+miIYqXh/Xl
DweEKWZPN3CNYy7A9Yj7if3zR95KRw2GXbUI2T5dT/6iJ9iGBHMEAArDfQ8ttPj9
+2HWIx7x13LbFzlEYlNU/qYrEUrnqmb4+6JPtZI5tJLeJYPXZSvvv6IIQMl6x7cy
wNTI8Rv3yz+PoIn+gxwXlkh2bktfs5tBGTGa9QC9NNYuKb+dLAQgnpX1hWaoqz/V
Ty5nTlnAWmz/HB1vHb7HJXkDR9zS0w+5joG2HEyjH39vN+tY5vgzBfJjW1fDDqJd
dVQqIDbv0BmKcdCF5v+jCM8y/ZYCEfASSueq69Ur3ljnwvc88qskQGXs/eu3D3/9
gEYLzK//oBWd1SncM5Mzu3xxRl+Z1anAhrBf8PAOLDl7OvYl1w+outxauf2Ht8D0
1i7Wp0J0E449eTGK80mOn47MBHfeaKHJ5YKb4bpgjRsFJA63k3H3pAamQl3tokPW
XOyFABqZERCe/phyCa29fdIiackJ2Q59ePa4QRHsNB0pJzYspyhQdP0KrYaF3vIM
6kBhTy7U0FAQTJTjDx2GokHFHh7L7EpL70sIooCCLxMjnFz8ges0LrqavdIbx6xG
1azy9QVkPxazmeTBl1ARRtK/xRvL05zPAED6tjderwOWmfRng7taji2PtMd8bjjx
DaBiqP/3EoBYv/SxQAURxk3OEFzXmEwFWs7yTGIVoP5G0h5GE7FSJ8G9ySOrNtFq
yGpZer0XWMJ2uYNv/bBY81qYkOrfiEwWe/XxNHb2S3B0eIjt9sjATpTPTIvKzxig
bY/93LUGFdcefE5EUStwEu2jMzebY78NAmYJ9UJy72d5nP8PsWjMd0U89762j+0T
C465B4TRh5sVGE0c+URZfkHGLbMfZz9+g4N++I1ra4iVvOeBgE6YUL1ozpn5ZRFU
+iiBDf21pjphx75QhVjXv/T1y/26VYV0oDiSwn57FpFSqIrxyquwcSIbrD6bjtio
tWl9ibAP+TkafXgYmjMoPpH+5AtAJqtCu38EzxW7kJipkVcEXaBqqnLaAdM1Sk80
KLfx+aLMnDx4li3wQOm1d2EpdfaxDmFl09hVqE8e3/N30LzMSa4TC/jyTAlxnYtv
xEUWmvbvexv4q/QAEEpWGVDCsxnPepP/ZukhzKcsM32T+JzeFdoD3ktiFJelRiQ6
Yl0CxIwYY9dZqJ0F7l7VWtf7WVsmfH2sLJAi/YhKxNyhyz5908AuE+esbLpUKiYV
4+szZBhwldgeF8ZXvkwGhWnvEsgn2N6nDSUW5rq3eEgPOo7cN6WRceXAKwlUBut/
JU/5WBTR2c0EmzhpEGbnE5eYChYOO79kUldPvfx9G77+YCnpsfvTkocvTmuEoOJT
uLM0QqWgoAfM9sbpIVtRxOolN90YDsdevgbOq1KXXHYN3XNyx1CSB5r+h1RKr7Bz
baxf1iOWsp+tylE2oikmhc2RTf/J4V+MtLhWY0DrLkI4eHJBDkBjJ42f0ltZmuLA
y08sgHHU6HA9JzIHHQkO44/ME+qU2YvUhV3+fQVWBexreCr1O7NUz7G3qvXO9Jn/
x7Kg7V9LTxtHOS+9pdEXJiM9nGdi2z59qQkMYFrc+aUDD15p6hPejgbAv1HYF1i4
LGZUjnzAWh0K5c0wV+ivmxzFROo5OMO8f9502M/f83jYMtbb/mYVDf++lgP4kJ1I
DNL08Ralj9RrUX2FkZqwmMV5NNjDuTAeqj/b1dhSfL/G/1pUHRrCTaKWzvRgsqfV
GFuq5hJopEWCRACuwuxPPPBjVKC/a+fM6kkRcpbjJQyY4r9reBNURjzhQalyqNn2
BquSuDr6PPm7mBp6Khc46oDU+loP5IrHW2cTfLf+pg//rbOIQECkhQ+vy4dWnaSW
LPrR3q8A5zh5CCuli3zfCXchtY32K6o5ve60w9RHJ47lLiqaA2PNHr95rEu3TWs9
o1N9vKfBiTjUmv6HOGDLJUifI0q36kB9ggyDhdA7ws4es1IIwBxAgRlUtBWT9MgT
QdJG0LceIOl/tSWuKBqh+AlzkwTU5ATWycuioNRqMnBXWZbnOWo0SAyIXy739620
yFYZBDjjh/5Kdo8kMnmaCxmeFzJnxGwLoHZjppT9Z8X/xyIqUF8EfVL6QhZvOUQn
qfOQuUYaRpIpSFkqfovgtOHc/WmR6mVV/B1mwg8Oh7hNxR20Wr0TlybJzBcW8fDB
2R2brxCf0YFuYZQ9y5QaZQpn9Sf2pQSPtYk1/r1mxS2OkEgFpK/wMicTrLufVnbP
7CEOTxPApfXCmvEfJPsh/LJAv59jwFcPP899aEvt1nZN4Gac99XmjywoL/B1k/rW
33a2DK8+nLFsOWstSAPdlpkD7lfEErCye1w6BDdK+J6C2K1U3Vuy69dDWGLlOqu+
z7k5t9nZfo2reAXTLSM1VkPlIJrDwE63wNDSu5vUmspgHvPgtbfNsIlhTkV3Mwq5
xYhBM4y3LUDoMn2yc47nfyNA/nHbmCCKibtOgVvgyabI8d2pbO/qx/28HS3UnOws
M5AGacH3TD+YuU/PP1qwg87oCEPeuooO89VXlpL9QnIbhV/4TRB8EAixIn0KGeub
2d9TvQq1+ddgNUlpeicYhTaclja3vrDfv4gbrWzgTDK2sWYe5clr9wLiIFVWF6C0
M1ap94kFjTv4IDlNEswZBrZVJPIW1V0xNUHo1tW/4mCNi9PVp2vRH8vaKn+eFzki
pecUr1S68xRexT9tpVLz04g6v0GOUwpjDcUoZFW2G/NMnsNLbUiti1eqsWd47vx3
bsY9ZIQ+tJO7Al7YgTovxMFAInUBcEMXq3bSu2YmYK48Kp8pvGhCSP22mowK//h3
unDSj6cyeFWPAsmMkmgit1gzt7L6X1nGiQnAOsJZ1ZEdU+ieJZOi3JbOkXcXBiWX
t4GqG1DebJLvOQNGirNTCYGbBksu+5B7G/6iZLT6G97Cp+zpJ3T7nYpNMaEBTj8f
MuHOFznqF5aRWGGAgpfKvWeBKA9lh4H6ooOlpnw8UvKb6uf3w51XjGTqxwed0irj
ZXVuplxwt66UYXLEPSFnOWn7p/g5EI0oYH9gpp4qq3PfqtmLeLHo27RD/bVm91Pc
XFhKro6mqc3Uh5wZws7j7vSGvxVAQLWGJe9qlnCbHH0R2xjgvmjjUg3u/mBG0zo9
bvkiKl4dMpZrbP5LpuzCUDjOjD2atPJQ62hIzkSZobwdaJ6F11xgUJPgvi/nNpxu
z4gAkTsk6ii0O3peaXBpd9RMVrXm+mREe6uf2a/lm/eTWpUQC4NfmuIQ3SiBl1pa
pxAY0R10iZ5Y5iXxUk/6XhbKTPzJeoF6ksX6yAZvlOvCe4h0XTBbF6vz/5jbOntZ
gPXd91xzSW8Kv5m8y3xNRhG3MxOAQcNFUhEV9fvvVldUxIG7jK5izKBmti9LlQNM
4qQ1wSZIkp6NuuRK8duBgIjJvpHbhfhqwC+7Q88DtGXHT7SAO3mONxMLPBFEhSuQ
C7j8L71WkK/JpBbKIek0E8aWNK6pH3cdsGbvz0JAS1ybO3D4RWeoUMKCAcBtf9Ew
e7qd1ln1MSo/yTVPjScNzLQw0QbxYILU/0/T/AQhHS21pv7gL8V3FCX8ygIvqgqG
SRVu0pOem+GPEWXrwQXoVl/BdRGcWOe52W2YmQS/wYMWduAebA2TRa5jOtTIrxRt
9CB+vPUvSWLbXt7fvmPl9c8ylfxCou8caBzULLXsRIv36GjqPv7dPyGyUI6M0y3S
DlNIqSKR1Gpx4FWbHgsR7h73CNq7HJoUIFY+Lro3Y90w7j3xWc9s0F27l5wcuhP7
HFu5ql9qSkFkf5XJRenJZ9wgVIAniKBJXAXlWk6MP/DM2NovNblVuhrrzTGK3pVj
Hx1yHAZuK47N6YtLCwSufo/v0p+t3i/Fb3hkSQgllVtsd0p4tg9zZ6VwUi5wmOjw
/MSBP/cbrfI5srB1zj5ZJgxIs1QPvITJf4c9HNF1Ir/qFjKR/QkZHz4KLtOSi+oc
84pNlOug80TO2r2pfpC/4Ns3pnVHqjtOj7C2r6b8hBby/e3ibN3rcM2Di/0wRiTH
u4OvuSvBJebFUcdlu9nzToEsAwtvkNB6UpuhhCM7ro9gN6kHCTr92SqAYG16HnsX
h62jdfZGu2hpj6tzN2XmaLIf0Pd8jX9l704umN1fGxKegkkUeZ0oFzLlOD/B0ArZ
au2PRjSpa4T64p3sDSky7PSbsyKg2z5QFJ5qdkgcTVp2YSuq5iKPxYtmDuIvrglQ
Er+Un5aFJARaB1XfbpqGhjewzdpdXFAfPBm13QL2lO47ZvNq97jdQoPPLTLaYSfq
m/z044oUkZl63jPKCY0DptcCwySojbrqcLDmbMDLkj6JnyBmN+01Ls8oz4hVfcpO
+k9ee4uNxzXry7Uf7TgRWXiuybnmII7tqVxlpqzeaQaxYrqFX5zbUBKXvsxr7Zbe
5WV8FcAjfLQ3qByBM3N/W7MxLhSJ7gQ7H8tsFYYGovTseeO2uu69wUiq+VJa1Y2+
v3zFeSqSIvCANTlQFXGhb9DSouc3ewV470KG8y1YcKpm1uED/pDAqeFjLyd8xBYj
p+hnbM9+bd01GI+4lCdWArIUsYF4YRj+2Kk7JZG6glSFPxFe0e1PI4bnoEqraIyw
zGwYaF+jhgirjPCv3cufOY4ew59sBkYjVgRMvFQNnXoq9u2kyHKWTiZrH4J4X31L
lkHzzDBeRICMpdQY+SBeOVhFXcptW/+oi6j7YVcyh+2Zj5oGQKB5qHcIOeWMIC+V
mcMc8I/xEzj7D218jzKtHgFL+Mf+OEi+tldvpTsWtbLX8rdNkaoT9eh608euVTP8
b7JWfFccdc3PWZ6MIVcMLkna2x/oJbO4obZM48KZ+wAGmRgmqnoV2NCh+LUMJDfJ
4yDv/AaMyFtgwZ4uaAS5+AOIYNd8kAOWz7LCKia89HC+Q79OHGJUUCNAUvzHn2ym
mIdePL3reIRCdXylyiYg2j91wxJX9axPURW99cpvAXLGiy7COFUX5BRY/pjtb0R5
NdN+ZvVYwWsqIYUyrGgdpvrjjrfaTn3d9riZp1VasxwnTJcW0l+p7F0tfO9EeQn5
yhVDUvhOhvjduI+pKEXB8h62GGAPeUivfiAX6RLVoZuuLFnN/hdKE8rX3yGSr36t
8DkClNx7JwKzu/K7qTnIhfk4dY1NBS5Il6irNlNFRnibA7dQru4EmpFgZ1BvAkdy
rAlSNFZWkTwkWnIT/QKplSe7fGNk1YFPIVfkCNRZbExouDedOCtXI7sry+1SxCf9
hKcgZ5895PxhG9nNdwYVjTDJGH3w/UUxvJbhrFZ/kmVwHCl5x1btcwZ7aHJXSvSa
bKBfQolowkAjTUBCVk/Arg6BrvtORuNfQRuJPpi8RY4ecaFTykN65/26iOFO72FO
yAfF4aqv+je+9iWS2YS3rtx+Mz+xFTjK3UIDrgyiob9tW/gPuvEsFOmU5iK0uCJU
rsK7QQPFkxBnwjJ4iU8Ek27bT+8318DXy0JSLCvbwlAmSHeIFv4ohZvXMhYwlfjd
mSDYoD77fHBv11hNSSre2AH6VODN2AnGc9UsnbeYsgHsxk/bRaFqvEbP9rLKGVYW
5xm04qlt0xQY2tsLx3VakvBeDPY9UOkTQUStJWyMpslZEG2WlxO2xOVU0PYhZAnN
BXtwgtGKzqOH5zOqgfue5eQg8fcSAg6iQk2T+nXiBD5eefCT7UOGAO/uTheLLzx7
wmjfWljZO8l0Cg7UlHXrxuIU2QhXul/EMjk1zLf+zm2vz7UIUE2PKjBgJwkInf+Y
jbGykYX2LhnGPVR5xjZVq8+GCOsYKyGukvv7v4dHu9XoVgLJTEuWrwhFmM9o1uw2
yaxFhk+LX5wYf90YzpYkRt3pVnsfkpXyLvDSPiEE4Z3zKgfSMl9Bu4xGqxsa4J0B
BtFpbMbJkyhGWbrmUUowumEN7KaKaU2FgZ4H0R4eNA2Df63z8lCpYSEbQ5WGRs0I
Qve0WxWS4jG4mYYAVSgmm0bSyHnoTLhW6yFXvcT/C9V0q7IjAlmLdrqcOFSytyAV
B7GM9+eauBgJOnyKp3NnOLqRX+joqyxuvN8hEuRlW9QjogOnZU49g1SmdTBKdKBv
s9JueFF2FsLo5wEP62lSf+Wh1W8SGVFnWYOBkj2MLfTHAe2z0Zai7svS0DKKft5+
59ARk+B9WWL6XdT/BWh+0YUjyQDHSU9j7SMSaJKO5VsYnej+Zy6lnFC+1ezFtCMr
Q3MFtML6mKXiFG2PnqW22PTD/phMFwVwSmITsXr2/l2Fy5wGo9yB//+SxAu6XDMW
Xf+P+IpV6aQSu/dSKMQ/pqEWR8QmhmOTglFE48XjneLodWrzUxiNeb8PY4Eu98DV
59VgR4VKKBqG4SBpDbL/KMyygq53sjAQpKYC+7sj23YsOeZVV8ebYdjoHQ68KvBh
4+wWLHDCOjkEJ9eqd1jU3UBDb9RV16DB2koyFffpDvg+TcFF1yQ1cvqLt+Ev7eWo
Zxnk4Ghxl0nXP1emeZOytPHbWForYWJhDXyA5TauUhbZf3Ud/WwzU2P9R3Bg2rUH
xhkeAio3MFL2kPBZb2NuV4+F+VkCcQS460X6uB9L5ou5i8V/8vs0S1HGHm8T9H28
NuyP5B+8XxgLj+yBfTy8pODoX/WL+M73upSCF6RVgMoaHow7JxW1JaGrl0JemjJx
rxtVMR2i+Pt8q+6haPLBjT2vuD/kZHapOaRWpiX34DYMaov+9T7irH55bZVd5MVR
wcELekSzUmUHxeHzkzV4DMwzBnXUpikhtFjmueq+KTGySEBpiYqp5u7mZIPWZzA6
EgeHxAG/ORKQOEBSSATQV6E1fnlzdPm2L+vQYA6l4ygVlQxhoFexotB9quGH3vxj
Illyk3CTjjMv/OFBzSyuZaJtX0Ul6Ep5ZozIHqMEiKjizrlMkbFZCNpIF5Oi8B9a
3o8nCCrlXQw6k+iVikQuGtNLQMZe8Yd8uufLaldQlapKTfYfON5zZSKYZzNrAV7z
lZI48TTBhcEXVG3FS1uZKYbFE4Q/fBdh1T7RFoCzy6g0ZiqD2vcOyfIf2C1P28j9
q3dlJY6o94DbfH/y2j9Pvdx/iIIvN4laJ6pUXGSxXvSXRTY2d4uypULR3+geTOIG
0mmC3oSISXpTwxiXpzNJlXhDP0hBT6smVWSp3WxImxRN3DgvYdZwGfBQM3Z2gBrA
cZuUE89puEL73251dIpU0PLsCAUtn2u9RJWDxZUJ+mRNRLI1nzb3ryvKd9jcz/rI
TIBY144Ak0hzlvi5eQ3yJDWKVDDrNT5MAnENIfHn+H4zAVV9IvpyOXpe/jdwrxV+
DJF4iArXiIjmW3NOQOBgjp9Hw2lM6it3+m7GxC9aMAGK/TMYQaXKa0LXSRg++I8O
yR51ULl09ZtFM3PLNmdUGMlVZyKWSnvOI+D8rEcNV5v0kr06Txk0QBtZGNkJxvzs
wEstAxDtfjgIsC8NLsm35RsUAM4qZfwSTZw8JOS+wJXjZf+WfJkc9asV8zU85h4I
WCAK7KWh9AZtuwW2YBRNrq+d8hR5Zid4CPV8V3y1kTJ6vIQMPfKXJ7JpOF0CjyGH
RsHqdbvfOJUg6FCAJhKdDX+XkwKifB3r/OGyc2+hdpE0TT4hykWjFvbgyk9H3n2x
TFVmfUMrbTFj6h2K6TEwEcv1F9y2Ai93XjYit/zsndbQkfbkBlwrDKb8NWXzevBU
2ovXSsYKxMROgNQv3VuhF8rCsC/rx1FZRtdYIeFESZmXeZETqAPDHxoNtZvowjmu
Tmatp532URLZ0z6nGlETY8BIlht/Aon3JJlICEiSEgnn9DDfY6mNNxrUm7eFZbHC
2AelpH5Rgb36Y6jtXx4PhHKxCcN+Deu1St9dLFbdmN/ycWXicmeAH6+RDxlgeC0M
j2nawNOHhSkYEIMx41aaKv7K+YExMGqWMH3HWEKX3yS7bPX/Xa6pReLfK8n5kdOB
RBFgMdVkC5DCp8ZOk587cVWI8fBU5YqNx8SEbh6QBfomH4KHBI856lBKfE8bnguI
SXpVrEVZNEp3s6VoK9p4HYMHXu4JPA6OHKM0a2pS7AMPfEKeGd8gdhR9tF13VaQr
aPKuZD5WRdHceSvMcuBfEyCoSeDWITt0xWrKUCcGaCVn0mHqiz4WlgSFyPqiY9jh
EqlfAyDVC2SE/qCywle1YcihbbB6gpFKaRVzxwo5CzGPFycsMBP0VMcqc0dO4x9f
w7EPYcUKb5tPAF4hSYA7fNR1HsyNeEiemm9jtlJJtMe2plmgU+Gttg1sx3swLvw9
tWv9H6Hx9372D39wJRzptpqLR+lv3cNvI3HdXCLHOtlW9dwXaYhhY+uROMjMa3ry
KqPXUBppEupY5fS7AcNGpIlclahx4zypm89mylipH5deqkDJHcpzU8X2qlHKfFws
+JZXkmP6IJIvF5r6SqzhkKCQcQE6N8DBXNUfSDP+rDOe8a+MSQnSLYWzPZV/S7Ub
xKsjDggI/5PiOuKTVXrCOowy+s+Lnz7oV6h6glWAMqed9Qc11zWeXMVINqte7XfM
biVDBeJ71oqMpXDUL+Aar7w37zRkC/N4sjtjYpOEUE1FKLSYXNhWj/Hu2B3s5b0y
v21yiGfUT+XDZyUQbGzlcVd4M+psAczssI8vy140apBbuv/eGmsRNT76xKfHyEHE
IUFbGWEUYO/hx+oRldIq99XFy2O0vr3vgn709/gn+epIuh7FKAbJagzWLzHdY+yB
koOIYd7rHW3Js71MMY5jVyYEFhDdcfJTH7rb2TvA1wBWO9y1JVPj1F2Vwl8VnXIo
9ZWUgKrpPtYQpB2nC8YVMuLapd/kby9lpDBGx5SR3p+Iu+V4VZDF4MwqVk4ep/kA
A8rK7Zw9+rX5RVD1yle2Sct99N0+BXbb66ZyhgXgrlMHnDU2oGGpRf49/IAbOur9
FXRdoOp+5Xq5Xot/hoBVAQIn4W0PlefwH2rJ2FB4ddK4NygswRjsDtVNHJlZ+12x
NVTDf9zbFIUZ6m9MY7JmDlBm8U3hgPScjYzoLIBghDkZS5BMBDbWc+kA8BVqU9Jd
yhng/NWn4B3XLT6/gjOFGW5dKW838BEaeysfPJm782J1ptDx9SSKqLZnic4qCYo3
rLCBmAO4DvgparGQOBFIwy2sJb0UscEzA/kjOKApbnH9lYTebDBof3QX6FJ7ccVr
gyt94qFw3WLL+j2Pa9bP+hYUgGcXDVUzCTICzbQV7wQIEIUeRK6tLZu6MUhW1dzj
ubiTpbAIB3vxL1X39XlgYR3V1DEdgPeFic6qse+twxuJqW93NZFo7oRryGrkXJKV
1JROa1W5KaN983Nmu2sE2FAB2ZFuD9tc992Xthtt7csKCr5F0xj/k9ewGNeIKA3d
3NNS+8jkzytkkZ2ShLfKSaByljuOdlZrUMQ6RJ1cOBasdCrk3a1od5vi17peHt5l
iL2nbQYF07sVsZZdyFb1AUmo/z4a8ccA9uZPfRosaTmFXsAYh/Rc9YsJ6QY3Bnni
upb/U6VOJ3Hki96hJayOgPqZqvSsIYcPKbxc+74cILQB5dUhLmmsMzHztKp1aXPW
Nltkq34FBFVNACJKvpBzsw/JF88ZCudpW7AUCYbhptc4XIte7IUSAyNpAU/bTmH3
4BZ+B2KGzR2GhFYUSQQy/TW6ev6ibDIBtXW+OdEk+tFlrRip1vxA27TZkjNz2WE6
stQdpJ7U+FBaNTJKld4nqgA9zorgsbc230HabGVSsTqJNS84lCk3/8xgc7SPkZE6
PLl+gkp0T2nXtgkvZFNPhd3K8f1PLJMVq3lZsr3IWgGcmd++hPXDYMD9/9sGVsbP
d3bO+oQSf7nmOqoVp0DCV949WcwMS355Fcf9gm/q9Jt+Ovh2KMDrz9BiYmHPq908
fqmAMBVjqg7Zeu8qYIaL6X09t9PBTriCc2JxEFbZLI40grSr1sort+GB21Zz6dPn
ZuezPykz1o51NJcZc/SVVKjkXFmt9zqaLmgHCWAGox5bQydMID9SYYb/huKoICQc
KwBJDOy4liNvt+rOsACZC5XXEN4SLY4BQVtili6z+9K1+aoUlR3dZsZ/V/xxfaXR
dxVZHcYSJ1Y2q7VYpOrUbLRWL19Vm0qArFwErOIJ+9mZSlJfxHnM1bizsahE/Hg/
wGAcND8+Y7ZpTWop3KP4U/IJhSFWYD87vJ5Dv+63ZvbEK6JK0Lc8sgtrB3L/c7wB
0wjrbrhNZycZr/F83NgzDVMW6ekRqdUphemFPVXKZqtk33MeHzJ6AJ8Ei6aScASY
mAwzuGRhJAFYBXAuurhovoiKL8axIaBdmXNn3Fu9THIUPDqiMY95+CHeB37hE+3X
K/52k4tJswhhRL3bGjxQEWDLBh0F4UajMM/DQXw+y5pq6Ls/eDpj7zeZoxTruZrg
T1npXpBrkHJptR6vN0v495cw0U/dK+bs1wlIt031F1VR2eNHHQv8TyqjKe5pt94e
1Ri3k7Clh+l2FrWOmNwDNnV50MN0icYDQYuMQhXccWHe6Fc6Vaj8HZ22N7C18yKL
mjY9F15FvEislQ/elgeeNe9YTIh/SVraRbf+pTs1aGl3PPcRwk/TKjnH8FDCcmci
X5JvkSFLjmGYVrOgFibHeN0kcCoVuA53lHJQrUI69ktZsk5/4P1+VO56Z/jhltO9
YHXo5mDzKN1HC5J1Zr3sDLbIqzjECR/jj+0K1UmMLGNl7E8EWA1X+QA0gYunkRxg
CQC+2X/RuIaxSzeOw5o9+1nv83OoqvTEGyMyWctMU0ak3UA6Bnwr2rZwTIPvXgIG
bPzC5ZplApfJLR4TS/G0ZVrW+dMWxLAfLSw6LPjbDxtgT8RAZPuxu44Q6JTV59rD
nMWsv8XSgXi0ti2gpTRsfUKPARVLN9nz+ewIZwmlvUdYH3tIKXDd8pe9ald9Ud4x
Vwu8DCyy3j9D3Zss2B0LSQ8ir2YyUBphGa9+AK8USXqS24BdtubQWTLmo++Wug1E
MA0x6sT5RBzYtIyN5IFadJM3bMRhLfBjIxSLPxCZVIeBF0kEUloJX8X50Om70MXl
NCzyzG/JYBZuOdClnwNHnoa8FFcf1nSrOo7n99hJnXQsokR7burnkDlIT1TQwvLz
g9CcqLiywwFWBrop50p6sL9rm5WlnU0crvnOoXDLXXjE8H4zhDyURkswOL0UMCyi
cYBO0bx++/pWAKeV+JzGeNkoKcKXb7+s7LslI7T3m5A5a+E7/CBkxVbC1/laKaHj
9valCAo/X3Ttv73WUDMEIfX9RnwrPCnKPTzeNXxwHihqjsS/wl9rFoKBs/AW5WHI
dVNK2ZLORJydPtV/mdyVNacoaGEAG8UdwhOiGUxfWlBrqsnKqORs1O2d4rf0FRic
54FYhPtONOD/j6K+RiJVru7ZR57Y1qAFR3bikpdxmyniFm5DR9tGlVit3+YJ/2nO
24URuQnOwYT7wUJ8WQ62JHQeA+BHEKtrPPu9r5tmS0hw2pklHjsi1kxQnLLe30nU
/7QdOePqjKsAIeKtMvAUoXStasm97lqwOhy0LV26teksd4DSq6n5P18zMHPGUgN3
4jSVYTUUza6AGJA4RGqafH5czeH35q4+ViwlsIhQICIG40L0e4wU6KzmDIBtXtzU
jaH0DeE2NrPOP++IwFDmagB++IrFj1ffPzmiCBYewMS2B3w66iTAQcUsdR+G4JWV
miWfUJuR3gn/mTZdQrDUHONmQ1F5Smjh88l+Bd0ZLzoz9b8dsyYVAogAvCDuux8P
9zch0d5hVJRED/Fg9H8RxgnoZsCvvUf8WM/AHRcOWasOVaJu3oEyW43kqp7yLjZ9
UUksAevePOHN+ANzYkprAqBIMnRFtLrxwx+5n0TxRhGO5jyDc/r8EN/+3y1l1ab/
flTj2qD1ALjSaOZA0tDgsW+QzpE7ZgI0fSOYGREllZe9K1LLJc00JeAehhgPXT/m
idTInvaMkFuZSHK3OK8SnHGD9qHB7QTQN+HoSZcVb3vR0RmlCdbaodDbu9mF2IHA
dpdOHv0LZlzjdxhv16VnNCrbGKXnbbhWHPrSNkj52yaI/vl6Q2+PPP49LBllfhdS
MlDBezWZOG7j01ielXiphg6l7ypwmv2n4NnTuNkVLsdEiq8MYu6P32FX3DAhrkk2
CdTyXRKjwLRsye8XDp4+uC5nHKDI1pyHM+rYpopD3a953CJ6PvcWbaho09daoVDy
zUn6TvkmM8CAVmtxJZkqHmjNg4NyUz+SskcKWQSvMyzpOEHlS6E49Y/PmmlPYaVs
ep/FIso2FCFqv64OzBTZYcZgjEPnQQiYBAF4UoqAwbNBq3StNdx9M2hSoZZJ7RA8
SuqjYlPyT31AJ7is8kCVFPdqz4NRHTlr6LzQQCK/9zIoNDxgdpMNureY7bOYsN7q
kTYdVnkLvVp1gJqZemOOXfM2KOvAWjYNX7jkN/68zxpLPElv9B4+Y0hY7qf834Ya
dvfC/cGDXVbqZh69Fd+jZ8+wNIoKspiZzXER0paxZv7G3Cak9NJx0guZKK/IIMEL
uYCjH6ZB/y7sDqgHF8CtymUx4nUYsftSBonMPeqMc+WLvrZ50aizdjfzgIFuZnLc
4ZN14uFvTPtp+jmnZ+SWTEwMXb4J10plsBrjxZ8TVdulcV5ehrrTQEru99JybucW
zEQWHT2pSlf14c/8dwM5UrAd6D9OIaKrGSc/9y4PRszPo8B8GAUbiLb8R0Wj7nSx
GL9raDATNoQGV0Lt423eZejj2wZZz4hwoh8P+QakDi1f8qiN+Cym2AUkgirhiVRB
Aqa8yZo59fD4WekWKFMKc6y0r0zWjb382cUT4or1sTt+lYoNaRG5TB8vt0DWm6ec
2JtkEKbOowm69oZRqVg7k+b9O9b1xOpnVwze5VkwXngrk9vKudsO/ELy+zPnhELm
wLbZK5f3ofhWN8fIOAfXBYiRWb+8jFuYBFGpwkmFBfMlQvwkwqGRmUjIizZvOVHH
5/HPBuLaW6NGs0AgvN93/yZhrckpMY8I3cXWnjSU2+zberi1zezI7kJSNWxCQD+z
+A4qBDuu/NIa6dJeDtliYpOAUKTfYCQ86BtRqlcRSwYL1TfoKxeyOYTFXU8gZXa2
d09dU81VtHuymtbR450+CuTivuJWRDEu9boscGh+0Tq6pdmIEgx9GQz+ev4nVPqU
/ThmfL/A0097P7woL/GRW+egnGOemG0Cnk+WXiwWOcSwP+mkkCDgvjhNVvnFsVXv
SRtSCsE9zpDcreOCA5ScDGzkSjfHSMG1eHfoWtcm3nppRHpWe4sXr9N3RFJG/ImE
ZTUC64RvrI3Gts3DVI5o5S6JzObm/9ubHnXnVjULzgZGY9YPPuIyrmHuTMtTW02I
gidm3OSmrcaiMP5INk271WNZmAghw39OvHdDhU1uKfSujMWoRMjNRlTMvXc63a1a
tyYRKRQkk/kXapngSqxbrVWtODYGCaEme0uGaI/GWL96mDDvt7u/oss1e5gjEFpb
E/tZX4D6C1cQ4rGMI2TqXroeZiF3jgH0o/+UG/w7PixeaC1lj7BkqNDQTxuFb7o8
B1oWiUB15NFTEdmlCyagnD6AOlBlC4jYK0hi/J2CdZ5PUH/Y+H/uqTx2Fsw1kLdK
afuHcnpdoygaFLKktFQPa4CQuhDrWuFduPM16DVbIa/Adn4mcOnU6JN3pO2zcXis
qsmg+gzbg73aAp+FD8bxD+lGBPs7kGgBRzI4EBeVJWCUA61IvuabrUzWpzVgDKAJ
LqbitZ1QAJ52LO2zOA8G/E+/elCxeVM3yHfQy+FGDFyTlEjiV7lOS5YmNiL4RzBN
2pXa+ZxlXvMJ1MoKAFB8tS8/gTKwxwCWLYzFbaHsxEfoaeJtQ6J+QnUdrxXBSVdj
z87I5dF0Xe00SOEtQ46gJqOSVi0Bcr6ez+nqEjhjBk4YMKz6rHTlTpBCW0k6GKUC
P6vbYB3LzPBPUcPfV+WVDIgX6Ka8drFm9dJCwih89gZxm0ureW3RskaJBKbGtIZZ
ARC3U01yvU7MD43GEWu2dePDMuxozvOq8FIMD5Wfjok1UqMrCePXGi2t6/cVCuu6
BSeyRhmDONgUmYJTOAUQvkK/QFSw3Ptt7vH/RgEqcviy3J2HUjbjZWdY9LrIXoKQ
+TOPI7zRDxkM+dEf6xJXjss8aA30J1ahkjypDNHEwcX95Xn2ByK5/8DghAV2Ump+
Hzadf/GB2I6LL0E2ZQDF7rCwj3AE4WhaxFzBdKNSWbqfyRi8UC4s55zFos+HNuFu
LLwh3/Tj7gd4hoL0ECfdiZctVMvWUc77UMYGqHf//fn3UGz/8bZ8DlENRBR/4yQX
H1/iqUBojFpP3gDXWJgD+F1apsl6dnr7o7bZv89LjwPls7qXT0NrxskddAGM8tSX
y5OplWEqJ+8BGQhN8Q33bIukT1VLHi+eqSewblB2jmTAHoQCAOzzyAud/uoHdOGC
N0z2/sOt8lhF/DvY3JcpAVMKY2reHCpKgEKqvh6HLn10wfHPGs3j9hhjRGQ5+pSV
ke65JLJ0bxHewLbsUa1wf2N1oLXeGx/o9kRDISirLjSBs0vw+TRjkhGY3Cz4+2W6
QLlBw6f22FWgLKr2UnX3X6jmjQnXnJHowWU+Zkgc+xk/vsJSqiI+3s386O+7ZAx6
Q8/WKlZw211y4MV9xD08fEjqrqeQm1rhk9DiNfcU3uTaxbhYFpaKPwgiJf5pRDnM
yZPPkVK0VxWJ9nHTSZEv3ec+V2dLzpk7fa0LrMVgT4vTxKZW+crtKR3fpfKlsxdx
yS95tGn/PxVwo9VLYOiQzvX7m2MbGRkRHA81tAAuta69IkZ+DAJyB15Ub8czy5EA
51gKVyaxKQj8JFPxSqQawuusobbE50XSOZa3ZRSoSKZf0V8ncjbuhgEegCvQ5FcQ
DQMjSKw/3IQ0J5Zn8H594FXX/iz6BycdQe2De1IlxXLMo5USbzaW4cJ+XnqJPXk7
RViwYE19TJULBXd0RSAJryvR70DdBuexxau5tsAh19lyBEBbersEmpOt/X95V8eK
pa7/wDD0ayI/8MO8+RLMEkX3legBkZZv/CdRwAUlgG9434J22LkPnxqrwnazpZ2u
hazqEcIgFbe+kT2GTGJc/s3O9MPNX4j744yacycm6SqSHNb0BH2hUkUSdhFLShjW
tDfGKo9fdgE224zngJeDBGISRyJMtgIH64GOXQJ3g04SBqcvfPnbTjX2tEsEZasE
H8Exq/DRElQUVs4RLfABmiw89HkmcUyjD3rElBd38qwX+duvEURZ9X5MJCafxsVO
rsJgo0m5sOJV856kG4z9mVz8WeHcpwG4PKUtzCRNXtjsUher7Qy6aX/uXYhQ/PeI
va16yOBSjELRd7fWU138hW/SGWWp0Pym1PxJb5qQx88g0jRVCkxkHN+PqK4DJULK
8jwXQTliqgQGGjqKNRaR3hfn+oSD3tX+IQEci9ey86WxKc8Lj9873779bzmOYwRf
rfpCCe3KjY1UekTV5JegN3nkaB9X8mjfUYoS+cPxPIcdF4a07R6tmtUBNeL62KUD
sqkgZLGhNLEhdrC/M0fTWD2/tpyCgXkwTC4BJd+sS/UUHdC3/aRa0/t8jCJjQz2S
uoxuNXESTe8VpHPXl50P1IDqnrxEA34V5vSbkdG06I6MoeFDOl7xITvgBDDD8Ati
DGu6i83PkpIIjhRR2FaocoeTa3Z0LYf11O1JzZ3JCmj8v1mdG2OoIA/wYhe7h2cD
BJLwq4YUT0lfyoK5uUiOxbKMXZmLQYPhzA2Sskfe9Dm7ZYpOQeLhHFooe5ezjBJY
f0taBlXc06ePSPjWLXtuwCNFQSGJCp0n1oQueLpYFu2du9xk1z6wwf6h8Cph/+YP
z82ZCYPmM5XmIT2QnAZVnArC0TTHYRYKjkmHl5AeW8YlMmaKtiCVwEztM7Tbb2ed
4vMYQhHb86Z3/E9SxedxGHl5WnT00zZ0kFvIhVlMY3mbVYESuXbe2DwgDAc85MkE
fJ5UMS70wvgDymJo6ukZML0csuzutxKRorneruleBuoNcDAFU71c+nYWvBLLed0c
XaGg1iUKAddjdmmoL0Axn3JbrOkNxMXOaADNSi/kPF7T5sWQebk4Kz6Ir2iDqP5T
0BzTOB3UGICcS1R8UQwmF/I2muKom9+wqaJgnhioPCEFtjWIylI+lSYDvSkK3Oka
7hDiFOIPdvqOjZ3Bxj0vzVVa6ta7XEZVhOjZfTWhgX4SzFWvOtXzhe/YJXbP0NnY
Eze80mz63FavUuVBp9YZsT5BM33wFTlNzxjpvnqye2YlIa5eC+4VXH3uk7SFBLFd
UwliX23Eo9qesoYoo6NXL5pR4uFZ+4D3WM3kFpa4H+yoIqlCfhlv7RBj7vpdoLtq
By6BA4C9y3Qs64XMl2IAKVIL8JEXs+32ymxAD3O4MKTPW0BIQqjX6WhwOACGp+wP
qUq5GA3UEUDTqx/mJagFcFdLlCbJhAzJ6oYWkYybPYGZHv/+4Ugz5/y03nA5eIHR
GBxmmhtU+6c7yLZenWJlEnA4rYAJ27yjn+FNV/F4OBhg9eVfZijL0Ikkhp5a8ZoA
dF2if5rpiJ0lJkgsvfmeicjrEVw/KdOuZyHPKdO/UaDbgA9AlCbSY1UmG8kgd1Oe
ytPfaiN8VzdOzyooVNSjDUei6xZpRQ1/zdg1L8AeV2XsO39bIVV2cf1vP3vbEz3b
FwRtzyY7+58PyrYLkWk/6KUSln0+AAURIQibpXn4EyG45ZPMsMP0hnViikPpzi2m
vM8OEkwnBq4+CElVoxFRGy3ZNRypH4Dfvu7AmxSheAdyBOuzmevheWBO7rleIGjD
3xQ6eS4qcQmZkA5KbZzYuWjD8kZJKtRwbbVzxmpifQULSzHijX+Ei808KGPA2dYW
2QrLLVqAjr5YNuIxGpSJGsi0wlhPzQPQdtWoQq+QLLJkdbnEJbfG7Lk63TzrO0/l
mSFF4gGgzcepRyH2tRQW4tuS4Kydmqe1oS9IAvm6f6nLFNHBdX4PZxPeMWT7EObd
AkL43Be8sgtO8KxRKne/U6c93yGaQHs4hUsC7NR7itQnSaFSYiKf8uGTsw5r1ahe
bGJ3nft/oE4GSMGhlOHmQTdZmA5JJ69SgyNY8WD5lzM73vENhYueOd+u+fIY7udM
l1QZDPtcpsdoxpAMtRRCMvsxJqLznSyhD3EHQff7wy8xOChXiQWQZUYpMNafrpVg
Q71fQ8HfGPFu/LNA2Wi6df/PzarWWNUEp34zQmCp6g2teVNqIYhM75Wvl2r5dhgP
ykm3dR5Qaurj4fhqZXf6NI6oXRnaz3xJ0ZQqng+VjUpamS1t/+wrgWyXGnDUMHiA
QcVZsBsq72gCPfhvNrn8DGGPfTIfxItQatZR2wbwTxnelw0eO8mTExY+HROk5GyY
12JQS837PuLKMdE0ZYvofuxn8jkXY/2sj/Z5Kq8eUF+a4T3aFoxsryBAIAjyuvme
1vojvIcU5rzv1EYIUeom2fxZO8FzELSqPXnQCqWqoGsp9NHsoQ6ZfWBlmb9qJbiR
ZM3oAPcdMnEIox1WP4op9XEcdNXPiEFngPdKftz1e4w2vRqoMB0uiZN3vSvD6cGx
jnnFiYH190sYry5dcCYWLdehTSQqgw4mcRTk63EOQXVAhqt+PwLbqcwEG40n7DNI
wPrmZOKiEELd/fg1GdLKaJOyyNWDxw7aL/k8i3hOJo9NAZ00DQn/yBlO9jQqVRAu
QnuJSlApYQ+cZkaKzOoaAeGlcMHoGzHEbGQUi56wGlt0RsYQtzsKNMvFDcOwiGHM
geT7Ajzmrapmc+ecIvRBHI/YI7K7kPsIla0+msvFmJqHJLNO2uJhuINkxTlXxUiQ
vW4mn7J6BtnXIHdpkOe8v+rm+PXqLaQrNR0QTGAQO8QDscsC0Kvwkfa3NwVoS50E
cQVq0nfZIy44kHZKSLXdLStHPefxACQXwohL2tmfN+K17c1+sHMeRjeFvSpJJeys
GZOghhc+Gt6dHuzx2lDfFiKOe0F0mUFHfWCmi5AED4HCfCxyZvzHQ5QxwgzJrOV1
/eFMwPwo95qbkjE28tBXhqoHSJ7rEvrE/+5I3zDSfTmfHtKjshksr3n8XHA0SkNg
E/Zc1uEc6XMLE2h97gbBf/rrhwB/CMFGBA3JwsaejS1YRdtM45U8eP51I0x0UkS0
wBO1pS3EnuPA9zrmjSDtuy3yHxVSgANMjj5kLHA3MAstPIBI41sTYJKt8C4H0G4r
ZHTP+RHrcCCNCuhmPTsM5EGNqGv8DYx0MpSRV+I3JWGY5c1B3pgLOf3s+TJwHcrX
J8plDn6srY4hjJeXuKp4RYJjtvFc/hMTfz7sb0hl+jPCgx8484XtguzYB/F6JRxZ
fCXiakthUHDpJQjNQAhW7shz3XqbevCfv98JlpPDNGZxMu4Vfzj7OBFQ88uZuzx+
Bdi3HEkoffZDaOBNkcMJKZocdwspycEXdTRqk/C+xkqxbw9vshk1eTlXE/j/92Gt
HnOJY2cxLvnRUiAvrCza5j1w3En1RApiU3QjpyP71EiwOiQDHKmHy1u8lKZZa9dr
yQkZREm2k1Dj2fk5PZFUuubjMU/QvFB1O3TWIUV6M2OGouiFyPtKH27kaIjPeBb6
FVwz2w+fMJEsf8aynYGIWKeS58o44xEIAPrfcXs7GkZwVbByz4JR2yGL/TJVyHVw
TGkxy7JRNX2CnvkI8HMiyBrYA2o8ALRzy/yqVoUC+8Zd4x2yyu2eDNp2yZhvqV4K
WqL8QjmOwL6p8hl9bNOvfV7/wL81IFqH61mZt0dmkmPYVaQlquXng/Kg4JAN55RM
iYhQAPUaUZNMy3pxY6vbEYOMuigquzdqNfz3qU7PFr0I6JiW5BuE4zadZpz7VPmF
bu0NEVUoBlpm6b0b2ob/hLxos9/RPtLCVvDS+pdGAO5xGxzSmTAGHRW/5NPOXQqM
vAR3UUvndiV6y0ziODdh9iySheyfDK11uwKBpPaI3OKERtbcYN6qGc0Sm9OV2UBq
GmtgooWdvGRB/xGDMfSBKXkQ0O3mACe0Yyw0np/xUxvV41Jkp84zQ3atCfksUvRj
QMTBjw4A+DeDaLEes6PrExaxj0cySKFafQ6GTDlIRxsaJT37C4wM4Evfn6huzrnZ
j7ZVdKcOHuBhF4kAIV0tWByGpHUsJDAWJsmS6/p5ZVlygiSuVNizlda8b1mzXqk0
4DT0iHzPdldVX28cqQRz/bos65igUtE4ZnFux7J6P6MSUtTZ8Hpz0xkF6AN8fbV8
AKkQ4JOPuln7FMUDzKamiVGfSR5mAITFAOS5xr5tmaXkxuURCCUw1j9icrMoLswN
mDiJ0i3NRXMSfElxcB3RzmljCBasM5V/hSB2o2VhjINTc33iaKV6WVWzL1OA2s9F
YjWJ5z/tgrrpAqXH8lC8XBpsoO5X/rRmDWzgL9al/SqrvIz40U7C33Ncbvp1PyDq
VON6vNFwEMJ6M52sd0CPrMSln6GrjaHrI4YtKjd11oUVOqctQnpGtPFZhCm5SOpi
Z4gWKfxLsKxviOHPv6xrrPUAnECpKhGE+J1eouobBRJtw9ZNzIlyM30jtDcSlv64
IKh+I/9lf1rJPttLsen1NRK80rwv6wGHnISmoTt/psfKqlJ5qik62EzJfTyLsZ7J
3SbAqoF9cR5HKsB0s0YJ74yHXD4jZ/O2DkxPeXFs3RR/GT+L7LEyZvNkE9WdT/I8
rxevvo9/bh2HvGTG5WC2+rbdsC7i5pBr4Z8y0zjHumeDWHjTt1bZpG+bi9IaWK62
BCkKvYLh9Il3uLptORDSbgbmB1o0BnZ1VmyOoew+lU0XAzmwVAIeA1zLdT4WgyLh
g+MvLIQ/gnvass8z51wDHgv1giWRNpTs1VdPdKivNLW5KYy5cY7fELne/xv0bzKA
/RlD2IWB58EnWF1bJRrC/aj9RYqNaf42yEpVd9rP9qNi6Svs8vPmT6KVkJRhL1OU
AkW+9Iht+1+YJjrPZusyRaaaV3c0fcZIdH9ueZo0l2wFQamMQttM9wI9d1cA5p18
R0Xa6B5D8Jz7dNkh6KzCE7ivNsAO7KfO9sxycVdsy7UlLfxEOuHMpCRA9fUmfy0B
LpZZz/F8ojpQiYEplyWvL/5eHQJRCdwXFAcDfvgOlWrAcYSaub9wflPpgsYWrshG
COSb7HTsbB4jF2GSAfsGprHfaI+/DSSSGTbFlHuzHepd+e5gWnuiBxA1bGML86Q9
Oy85KILO9A5kZQ+QpagwhsuMkpCMdeQrnqSrMRMp35n8CRmPiNcuMFBe2M1Fotlp
2tYLJTXDjVUxLnklt3izpN/vfGBpbJJHHv5GabAz5liamY6y10zFXu/KXM7x2WLj
sJMzco1+OSaeIYC5PzqdNad/sSLjAXExoA7l2RBoPn+GolDKnsHCqx2a0IDCVlYI
oikrzRUv9IN5jnH/TDJtR5JOlXI1itvFMc4UNJK2Whb9t+XtJMm2kwWDVJO58piV
san4hTlqlJJi38wowJM+POaaqgseAJpNihRto64zfybMIAf3WUZb8RE1UrU8Z5NK
0g8i23LChQmCqATI8Li8rsrOrn4IIgVbn3UIwdRfQYOmqthXduiVurJ8n27X/ZD3
FIx62x+mq/iNS3UJbR6X0oI49Jm9NteYBpHKiA60fsJr6T+xT2q3J++ureaRpUmS
X5XP2+P1hr4QKUWSQICG7aTkbenbKZMVNIOOdEfZBHyk96l2C+FPxX85DYXyXvjN
YVgPnkjmlD3gbIeDIDaNHQaoJPq2NAQ1d/RN2nn/hxbsuRsdazz1OeZmSnoY71DP
KQVkjcloiTtvTwcsmGNAL8NkLZua8k70u/TaG6JR8vcneKlRqjEBsp9dOgLEqdSO
1fwetM/lJd5rKlUkpKOi4IcW3uVaBvtP+gKdcN0rkbBR7BOKwEb3gOOEHbtSGoSX
6NQNS/ky2RZWtx9R9Us1tgzOYnHJMtSQrcjx5JKgOQNFMP0ad0z4yqtNyAsI7sNw
B3aUoIbKCOj+lzayMqe4XB2kndfcWxc0v3rr2qJo2TJe7f3EFEFw1XbFnZImvfS0
eUFkfHvCWz6li9Y9PZy9YN44OvKXDp3Q+YQGaST2fM+XQmvy1v4dUe8blFJ21flP
N4+3d+YLqNB+M0OFS9KppBpJzQvR4JVS8wQblfoBQdC2jclnPffH70gqGgeMIbRk
PWm5W6kBYnkvXMqXXDYwozozwafpTDM2XFGoMPrNc0CSjBOGM8G8DGoSu6J9StuP
xHhuaxwjUWwM3QpzBN+f8t/5jntbfSphvyhi0bcNOs9LCy16fLqZ/tehxlfQVzvI
DkCK1o1t3EH7k5NptpaIhxA4Hbz2EdnEFInh32McA9h5uEKtm1vsIh7BqmK5eOa5
O+frCCsW+/+p84y3WCsp71dAhLvE75g1v6U4J/BRqOx98NiFSHfSNwOPwSL8iNbH
4uXi54Z/3g4nMWsePQ8FitHxGxPK+v2TwUWPrth6GXSpYEA6exR0RrQkKYmepiKa
9jdGJz27DL1TmMlodybKkmenNR2ugzbg6nj6f1Qu2nEh9jNCVcTUsaaZ1ldlBe5K
GNvdMG7qk/wGGzRGF58eHXaVPjnIxoATRiktYa7hq+Vk49iQghujm6LnfWgOlWmo
gYBcnARDG3+JAABz472rNJIZ2XzwMdIvKw2kZSxpbyV8GtXTgRhmq7WRS1oRX1zy
tdyh52+VsmEAXxGGVjr8ej4+ehZa0VosSSKO2gctmDSK+9E/RNkYS6Cs4WnG2NGO
rkyZRZFqSOKWeAkTWNuzM9CX9GgPL8HZiA076JRUFHdiQggAKgmiGgvp1xvGGXV4
ldvf9mH47QSO7btF5Ayi1tVqHCn6Ocm9fj0LKPz9Ixh7vNphzSp4dDbUnx0U75c3
sOwRdrr/SB61g0tcqBi/f2DrmS0ibNPn6zVYg9DgYgOxhBMj+O6knTzGRH/yi0Ft
UH77ZUiU38v9DB+kYuF62D/KpaQAT3G20GbNb8zc33xNiMnEYdc/WtNWY8f0x1ap
5DcyvEiWHITk6Hzjk/Zc+WyX2CCsBNp3qN8IjMKts75RhH7E9EqyxpMULyslmMxl
vYTPev6KETkt1ypMOAJdEUcdd8+iinlTRuPa6rOt9S5dUV4FMs9Qm9MgH+yoilHu
94Jwp4SR6pTlDpDwD9ilIABQTqLS2ds25mXmJwdcDDJpLKRb1qvbouxo8EV6Z2lH
mOkPUR8P1k4bsVwA5WqMqQrcCO5EIsaBo/rXHxwpOHMURNV31F3xJHImvuENtL8Z
dBwT5xAXHm7aAmGJiyrFiAi1eKG+QpBcXoxCAO/3wXlwySlX4QUWFS9xhyB0YbMF
af1NhvYmt8+JqDc3icC69R/Q2M5jqoZ2Em9vD4TimKEHjvhfe5VNcSnqhKBnrgcC
VQSxD/Jv8Is/Z9yC5fx3e0GpyKt9Hh744thcB2eHboaFIIjKPcQONQVAt9ZjmAJm
uuTBHm2hykkvQKa+2hltFMU3iRwHqdtTQ1gE1GQrvWCay1aWZEKI/dpcz/FbQdUr
6nTCLgab/YXdcn9f+dlYUqmgZicT6vV9MekfdgOWu79sL8UxOrKOwMDcPU1ju7zC
48W7p8Zj9WoTXqWdMt8ZAk4Xgq4K8UPu9J0I0Q5zxeDO9iecWMEbGHQPgeMy80Bd
2YAsD/SRXZRJ9QN1TcnHAKILxBtsaAXs1+IKWhw849kK4LuOh3RqV8Y8WFdc/pSE
6kuarQwhlu7rJRri9MEo+/7nuGsEoI3AgUBr4W9jaRWVjGcgHWq900m8mW8yuWhI
3ZzeaFjwjTMsfjMzOd3qs+M4Q1nYeS3HoEF0Aqn7CRExOZILQfxcgbDgSOwxPcM5
RyNKmwZvvKkJ+t1qGhMOddxTzqAYAvHYOdmhaOolS1v5RjX3TWqHpXWDgBREjdyL
iCGNUM16zttv498SbmfKe37HsEZSUSZtI+hmkQWiLa2QwUsi7jenwx9Kgxxakrl8
hFu/ydBb1yaF4GaHVkwJuAThIK0sLu/2wvjAwqN4mf6if8pMwOCu1ODgnj0udmTN
MnbT+FK2okEDfk8V5JNAdLw9yAIjz7orfuOWUFDWRgH3vErheltoGkVWD41gssmI
PxwuqC2oiI2mikE318ZB3QWfovch1wVD94uWJsoJIAcbM9HvdvGCFVLVjcMFy0Q2
fXSNu+EahmKMQmGunXylgoNjkPmWe1MJnG2ZYrsCl1bqyILPtz9vIA7e7ZDLim/W
m+b9Lt++148nDB0TsRKjcKEwXNvgZ0lHF6eks7MXtcHgg0fEnLTD6A/RdjlC7171
S8GH4PIrpbXpSKwAF27phwYUL8Cm+qAl2G7gJxsd/vDLlxTzXJwr57faE4ZFocNY
azJRYun1qFxH6mjBpGmqwPn/shcvhZymVNIrS0n8UyXmG7BBf8ht07R4KPczaH92
G3jYGs4h8eQ8vSc2qiNkXbdiOFWc2GQCyPIlXk14zMveoPdJR/UCo7fKlqgO7FeV
Wstq/Jdt3snzXqZuYpe6kXt4VQblepdjSiesHOi8lshJjOZkf+dJ+APXyFTQMBq8
9AZMllgmkQHNRm8mtHTumIDURpTncDsJ2S+CuNqeRE8mgL8evN11HtRsR6zUbMVk
pZDTWiFnLyT/WObuksM0Ex9v/c7CqGxOjSAM0Y9ldYtU2cS2Xo1E4lsYEEtn3aBE
v3JJIf6EaeE5h45BTuMW5O+fiTcKILRJHR+GqbCgqsiDdU4rFqmD3Pb2hK3u4NTg
Hx2Karkt3Nv170xX7h1VD+Snlfv5qvqMwLYl4v9wtbYMHuZoBY7LcStFUKjMLVjx
qItlkkHNco2OmU6UuwqXG+4ft8iubHAOHmRPneX91h2ZMxd/ZCYUUsRAU0PRxIBg
78gyqhWXJDASrNPQOdHog6dYbboLhMoklp2r7GIFWgixCL+AJ1WL4p3aA8w5mC9D
n1hFo6z2BE//wQqFpzLSAjuL8Qqhbr71fyylC4DJ2foydKyJEvQkNlcdN9XEd2Es
elNELG4lccU4VPJ0F1FdxAtXguxkwkhQQzQCp4D2axXlHJXkxd1D1RpppyYoSzYx
U522Gs/lMbf0o2qK1qBLjlyCSAXdrRdZojMJguaw6QZ07Zn0QjlmJOeQdiH7J4v2
kxnNHSxJTVWeO0fv2B4yM5Y7M46b1vuHpfKDcbFl8gyDHekYJSv0tJbJMVHIcWbT
CniLt9eElh45D7daijSMNJa6hVzdsvBekFu7M3G26iHtZhIVomqTeGbGpPaoEiM0
iSsGbduNoj3AaWMz6mTdfBct0JDyEUMbx8Ug9LOzGleapagfJ3+cuBPyAk1jsNQL
iFYHNpUGCI0ZW8CHgvz/tYDNgnXDPJoHwwSa+kbxPjqWopttN5jvLgXunqu2c0PA
dHet5zNDq0lkfqEwXpqD2a4ybD44XQOMFug4ap0pLNe91ZjbW+eydkJeuBMJ4pvi
Rm4Wylzjagn3X+cLAGFZJe72uMIvKI2ynlcAsHDm9B5s64sf7Aqz7fI5QSWdELO+
joo+lSB/GmcLmUGLZgDyPjBRq/8FwkJZ/5ts6GX3D4Ydm8U28K4COmYRjZVw8JtQ
nuTH6hfYEm6kSNjrC/ldR+OrcSleWmqWtHTWWnNWv29mjrWRW3xxiBcZ/gaZQMJL
KS3z24fubUifMU5PrgWHPYMXAYnlu7ozWyrNXOg4LFAwYbOBMIuaNEVjLAnS9j9G
kLZVhosmpL1oGWiKnA21APguKw4CeHFRDryR5NLB6x/vdvjMojQg7eGL7u5pW+75
t2AcyzUNNUNsGo9MMFnwYjqDcEvbUslVPNW9YC4fIZ3+aBUib58WSDCb7SYnUsHW
MpkO34V2dgw2sK2WJE9BcmFe63NGpwSfVitiCk6yl8j5Ve12kBPa8UY3a12puwst
VcsVLIePawsz+/eekdxIGWBsqWeJ93X7BZxEGWwfOPDCAByXKMr3XzDl/hE6pJPk
AEhkfZ7lDHAm8N+aMWvkjezVwZdsa6Gn0G7GZlIqSsqVqfxHpjPib+jZfqOx9f/V
83RCA6swnq1iyHt1hYnKFQrO8tnj8RhW1O04KP7T7fROq7atpSr4/Ri0GZq7zvvi
TDB11VP2v7afu6oIA9GjPB8KXsv4pckywF7M+mftr2I8tOIanwSntXrk1+IRqMQF
ki8fGyUNeIesx5bTVPFCiIsO2RRHRo7dlzdaveP7P3gGLeJ7PHe1nU7gKoD4jKxH
+eDSn3lKhxRiwmypZmAQnYpTCgmq8/0S6WUGIljVyUv07BvfpZjRRa+hwZPLaeeH
ULd//mM84V9oDKrM3+CbhP38pX0qgh5aNsjSPgKJVXbfvVF6KHFydDoBIts+3BOa
5NzBVhCeAOvf5nd+q7SrkA16duZVF+mPHEIDuX5WBsLWfVXxVS3LTkNXgZJawyFe
bW6P747LQsApQTq6mRZsJeJNSvkRvloKS2gLpUt3N5OpMGEmYd9ZFO4rYhAwXr61
02KuEOChC0cB7t0miDZ13BR66YrnfdDqIs/Z0d8QlcVmGgrEC0ci+UaxHdX6HwgN
6D5IYuZE9IOYJukL9Bsz33rL+LLwl3KHcq8XbduSmp69AhXINFuG0APGRxkOkH8Y
4eUt0ClTlMEXfCP6ZueMBS1Okt3m9R4TgFyx5UwWxAXrSDHd5thqDRXABIxmRkw8
Ynsw9+gps5QHdFPPhd9P55xrB7V8m6hfxwvBOWg/MJTnbgPD7eBzsfqZbu3esm5p
WjsDreiks7OlFMX6iTxZT/Z/DhneAvsNYZ1kGEzDfoVSYv0hCfTtjS1kmmrhJUwP
cqjeA4HjHYHVlkW5sQE7D3HCgR364SH+A4oUmVvBrh1ao22IIsjmPT9ye7v1sWtg
QsugHD3mB9okJ4svxaAUya2ORK4wSp8hb1w5rfl46hI2dP1ueIK8EgmE87HwuwJ3
7QrM+mTfnwnmZr89UlvunTpMED2VdTRU/1WyrHAX648xIwnBpGjPXcvmRRW1Mwmf
DZVLoANa/xd8ASOXCHH08/9Go+oSM4VR4+TSc2T/BdgVfoY42F0z+CAugGyZa4vP
2pS2XQ1zXOLvytfKLJCesq7Yt78lgBp1DK1wtJnUdjU2HU8HQ1TqyMq+j9H9or43
b3FtmBBQDYeeIJpXpv2Uc1+qShqKnnX55lzJbBpBTraOAwyPzE0RCa2Y3FcOjO5q
nm6MVCW+7YfG/lz2Pkk5YNVwj1j1NR+QsVA7DSARq3vnd6FsCyw2uR5u+Z6IENdW
8AlCoiAV/pheZH69tMLcJiknkJnwrMCLhktMVJNTqR9yJdmisRsPwVLyGXaBcLJ1
Et3Y4r0M3EqfSQVSZWpZSoFOppo6qOGzKtuldRuRtDTCfAdlUyWBk0gC5FoP+zxx
CoSttKsyGSgA/ErXruvYI5xtr+7jnRDHXrzTLSWYZ6tBE7CaAxXVCMm7A5kKI6na
QsOhyVpXtIFCgqDzPX9E0zuYirq9tWLaaklOeLccOuRi+PWUuJUYKpZeCbaOZGuH
uEjqkDIBJHbcVRuvmumXMu5vI7MyOwZ/01SnRWQC/vOesLT9arpR1I/r6XQp3YJB
emCyupen+tRwTiYXEdCCzlyHAiK4OaoEebVpA/gQ06J+Rj9g5E0XfJIQqz/l9STW
zl7Vh4ubm0pApflQG4EtH21kclR8uxtBZpxNQXDg660rbAyY9JznAqjN+TspxnnF
RtVfRDUMwJNmQvXobM2Jm0JeoyDTykr7VUAvuq7cuQmfVNGhuiveSitWtxViJBks
XLrbUZBr5DrZoZLAgKBj3BfG4/eSY23BP+JxwLM267KrB/kFGis+tERPP24bkq/V
s+2ZX8vmVdykn1oT2sUJVl1lO2PO6Nbrfl2c5g7CH22sLqkNCFv6MVyjJa2eY0ug
gpdrJvw53GavGoqaQCSmo4Otks0hJ8Rcxc+gjMZqUc2aLvCXObcqL3m1hDGR6Cn6
9WAHfvjCKYAF3WTF17vpEk48QPuc3utfzRYmr4eAbBm+UtB0bCxbfYvmS3XYIaRw
/ZBfetit0Y2MUSWwwE9sg5hpp46kk8Wt/oVpw2ZeVCbeFt7tQckUmkbTINIMGAHE
Arv2LYFwIgqvjFBanLZ4T23QOgyVUqAshBCt3ozKa2crdyoITriXmHYu8s1NTgm5
qQ8uDM3OWkqokkwt1+nqm+O4/d76HKsK1H0jOqCiBohRkZazlM5Ke86csMYm1Gt6
qrrCNSuBSNNblqpw2fvRpD9bVjzBHXV0AcFup5kwneM/R7H5utvkkELzs+7Azwds
//3PRezfuPIShlEn3YSsprHQNfbqN03AE+VzJwq+44XQt4qtF96Qu3L1kCRumhWI
i3a9gmq+PNLTgsbFb2xDqDXNLehF0COnUcdb3tm0Z+1WRrvwwqGk5y3btXrLw/Pk
vNoFPotdzN37JdR1iqyLsJzfzgeQFFLmYZO9OvzVM7umg47J/jv59MWazV5xp2jM
tovrOBstL4AF5CIcRVEa4ZBC9zFm25ieeR+loKeYbvuczIXUGfPtxnVeHyItE4zj
PpTeiX5MQ6jKNJDNwyKgPQzHOZphclUS17V4Gc6vVnQoDlhBdTJ9xK9V8GWFlsEx
PcTBwWg5pSxO8YmP7IxVzQJVMryKmtJ5qlwoB8t9afIM0tgWbNZdlLfNvXaiYvss
sl+8XuBEb5nlHZ0wTdf/LkJS24vdF7UvBYvaizB2OiTQPMldTJe3s9GIE0qPTR83
y5dzD0JWtTntYT1okR9Ozxzole8Lh1q6IsFeYONrsYoAS82T6R4HDf/ts92iBl8K
V2yILt1rnCEVLX/dUMAozvo9+KyevDzLQG3T7/gDlU/3OUPXKcUxiZIy0hS9x4ty
GxKr6oYuFq9ZFmNG4QivuRYWLWBc+eIuSiF8GxzNm24Efi9ETpFfpc6j+e3kH1uT
Lpn/RmQY03T7S+EjfO+P/t06cZNkWXg69Q/GbMstTv+cM06WAUasLTur7RjLJHCX
ZoPiJSmFld6Szs18eSw2j1gulHcJOr7fxBd2sPwmLXsD5y9j1OeMDZIq9e4twoAI
624artdwlDTdmpuvIMbihKf9RdX4MqJvM2ERIkfHFvUMmLpsMfsDzxL8EVTmfyDL
NBRoXII85M3ofFG4rOj/iQQEhDc9a4MAeptnPsm6WAvq/gkHK/rIHHUV/a/edwVC
HP/lMFxraOZJBfNmTWKQc/uTPTZaWTq3eZxaQU08hf3ZZV9JYsDyTkQPVHX1d1z0
kOewigl6eqf7gP+na/kE72VFpUTlGEee/0+uWppuo4Zxxlv1E4RCNBiW8mS95wkt
7ZPTX1Szp5tBTBnjl2KK0BgW+vgkrPLFLuU5SbFwXCR6T8S7stP81momQIqjLTKX
zlpd8KWV5b8O5y9wO3NpAP5FvQ+zB3iSVAo01mPuJ7QIY4NiuAhatxHRDi4/4PUY
yomg2hSQ7DRPojtqJfksG75jdtdHhN+KMS6olVL36x6kDkQKTIbbP6I67I0DwPNJ
FzQhIOCEI5XlOYWwc69eKkgBM2ZRBY2Anp6rndiTllM1JqaOBQKPIwbE/ZJL8XGK
0dt38EukG2iGdxM2U7GVhl7EWyvAV1e6MpNSB+5IQgZU5fGnZAeJebfmPwT9PmcS
rS0qxc3iaBG2LNl7h8LbKiN/9/+9CqXs8U/wWjiS5GA+M9k8MD09d+bpJbGlbNO5
RA36oJI7Mw4O27F3PiwGCCgLoFi2z75DoGCaXz/+vNPPzwHmLD92EnGMTfneBNOA
7QQUN1xLfjTeH0laL6UVdFAzDAmQAu9AYUCAlgQB8CPB5oWDjeAOEWyVpwGx8YwE
+hxqWuFux5XmE7aeDRRsUTAupPRDSVzO+LryrdGQVVnF5V8zS8XQ9DTPmvI85uQD
cvssEd1HNnJQ4E1S8MqmpwLZtig30WYqBvwcg7xy3JL13a1EirA1fuRoAoC71Kog
3+MWrTz+T63JCkqM6x1mg/yKuhrIsbzQA5QH8OWU8eXhhBeJjHoH96usejXOAgJI
I15Fb4ZO+VgWOuqN1urlxW/ystgxB5dgTFgTfLoHTRjOP9tdZaVzo8r58rZqsdWu
0uBUTSUPGqbgfY886qQf8A4FTBVtR4x8DPQp4k6ysQMWn4p4zrr6slOf6eVsuNrL
CYzTewGcFoOZcrG6H2QDZuSaeX7Diwz0ev9tw6hQ6ypfWQJAuq2kKj7UksBR+mtu
rb1hke8cIm5/3cLz0Kjjvg6VCAcMmkN7r7xcAC7RYZzcqlylIwXNlAgQGjK+5B0S
3/FGXFzQ/hyyGm+JY6RXzx9bmrcXePI0Ejki+9euCYXKlaBAgqIUaJSmRG74+FtM
zRYXDkVyP4zmRMkqd4uIGDAV6g4ffAHYB/84MJIhWaSRwWA89i1PqX0wHdOphz5V
EdcHL+hlxYEUD1fZ0P34eaaSkLqz8c1e6nBn8BsS39yKT+8gq9xJRD8WHG4emuzU
heB+g97iAStUIdjtl9RQHNRSzqIApa39hcVFnTMqC3b/hnU3G11bP+NERQRAvqLl
DGmcy8xuJRVgQ7OPDdO8QJZ55iYV9brmxiJYqfynVcY5kAlWVjysWZmAiR+K9iJH
r3+EPOe43M5PzePlngXPKBORYULvBo7Yfei22bURLN7W++ExDJWbanC1fSqHB7Ex
D7ahkUwJ03S3BVnIBPxefHudM95Ri69IGrxTKv3n1VnP9erqK8KhbyqzmC9FWAGf
tMNgCKw8Wdpkoj+tpbmmhZy5WU1d2QQ41PsFxJ/yW/j2mDogMjxVWiDu8Xsx2p/n
bfyjOeuUNy0EfqeWdA3BU6E4wowHT/f+s4MLphbzZfKML2wAJZ9R2tzgbNlO3c5g
i6gDMgpJALdaKLq997zSWx1dtuMAu6Uy0qRv66uJcVvmvXS6VwevubYfFsVy+r/v
OFtBjE8Rt//RZTNL/gvaFTu5ncCH5Ux5dl7XaOJr+y1EYOZJ+L1yyovAY/aJ92CX
qjL73BSL7tJ+wZ4DtDMxqPCPetguNSXdge+H728M1AdTWnmZcwOFHTB9KJnc+Yoz
iIpH03qz7mP4MwuoOB9c756wmEn0lwT8wQfEIm/cx9RLUZjjqIeTYaJy3FuG/Z6t
qTPXw2J3rs1T6PQdX2sadpIJ55jwMb+aoeJfAeu7cWC8Uw0UlM59EgR/RGbC1/GS
l2h2PRCM4A6zBVHM9z16A1V1IPRoGSGCUAABc9/WHeeZ0SFxetn8cVJr6yDRaGYK
SI4fFU9YunUkRVnBWwq2iagzFKb6s/7pP679VUmDiZJ22p9rmPc0TbRBVWvNxhBZ
CV1Oskz9s3F+qgcYSGxiJVeHbtUjj6uDK/JC3YqrRXi5M/adSE1zijTujG9+zHyb
E6bZVYBn6JJNPl7LP1CXE64DJQJ3o3w3X/KB+IoXK4SDEd23ph7jRyo2ybp6kih1
nnDswZR3fFnX75HpdbDfRqy+5+M9es1XJHfgVuTuBrXgWy6E6y9KhPAt2D3Qj36R
qHMX82Vm8iHpIB7WHZ8F3YIOu0n45UutCw+Hn7KmH/U55+rY7dKVii4q6L1JCngn
vM1Ub+PgOFAIoQqgFp25Ovl2499CwAQXS0qLRcEM5eZZY54rR1tkmScp7//OGFyv
ex/maTkLsu9v367oxjxkbYe1jVo9+3FRxNkYilnwpk7zEi5utfnVADlNE2GYRjPb
CorxCN0prtmH+dYgyifcxw+b+7dMcF5lT6ZpCVKt1rTSmGFS68Ua2jVpmf7LTK7B
QEHsbyGWmU7pGXuIgICILcsUad7olrES/YuylCJMFtEOXbLvVhwcycqXP/9yeMVJ
5HUZ1kj/dqn2aLPvhiDSkFAHg1UeznSKAYKEb4jUYUp62CPMHDhmzCX6RCEKE4bT
H7vwG3hCMbQLYHGoRY2DuUk8GPsMkkE3QWYnJjrKrCVXGCF3EzBkAa9AzaTLklJO
KrkolOw5gz7ZoKradPc8shIy9mRp2sRcC6P6Ep09aJygMel24A7FfR9tIfrruvNC
n3GLjuM0mNYG5f8JmS3OY7Hb51NB489SqkaIrDIqqdNF/MdHKw8ZcqYlIXoO74Ox
/lPV56o8npQRfpnu0/tAvrwqGPMP+tt4Jgjm9UAdOoQcmoEJMpKs8niC6QFIqzXF
XCL4XfEEt8tqgdL5j9WwMuymmJCL05SRVcGnG86+LfIiJqjpTU6wVU/cITQ91cyE
vnAFl+aBB+RO4z9hJsnWq4dOU0tEbIkj9xohOACXDhbvwSZxOVx8I100hfYdNBQm
SopOKGj4n33mFaWLXOGpJ0iTn9nXLnCkhnTcVpbK51nseNdtgVhjKfu345lFPPJ6
FBk+8Q4YhgUU7rqJLCGq1Fhd2XLl9Y8zCyYwJgRDXIPy+Bdo1ZQg9rdkdfa2QQw2
FrR5r9SNAPjQhzkO1x+ZvJHf0lU6rNj2hi4/5Wju8a/bJsrqwp8WB683s94qz0i0
zp4ZiV3qJvFFn5zBMRyOz+BgWbx1xJPucnRhJq2545lDtYqYeblkCOwe4+udIufb
fLZ3ZNrtLB/dS2LIDPmDGH+iej+kMwtCl/uyAOwjhCu39TM70dBu1Q5kOgR9fzJI
+z4AD/HKopHfpLU9BGc3Wb6M6UjZlnUy93ioRd6EGNKi7WvnGVi++g+0EzAQCpzk
B+P6E2gnrFPK7aNTXW1i54/orRt5YCCRw9udnlPEDLnWvMzwt3JKiIMhY6mGTQ7W
ztDxIRC5dc9srAGCsWFvgGr+h43tR3RsfTIWpPNCNciSTR3b5jSF8qPXfiegUvs8
ubTmFOKTsolSPuiArhaENd7aTU2o4MrKcm7tvHAw3iZECzr7pCmG0d09Xv68WK73
E+JhPOhwa2F7bB4akWYD1xdBVPennllGnndRjTfDKlioKWaQf2U/CArlQcc29Kp9
08FqDZem11mqPkyjOUrfCfLANxArhgV1oQX3h7/ON5NOCa5b5SNCGkG6srsx3ZVB
0djQLkXzbynyBqHtPfOztQe/SqPYCr0GThKszzl+NGdiRmHKNE7q0dmb98+b10aq
60IeWGrP5kb4hwOZzc6RQTqBYiyp9fZgxjAJKl3Tzm2gmJKfQchdTKe+D3vFNeB/
myYRsOVMnAr6A+ma8dVuIG1sCmqYpGocDGds9qqaKGr3XvkoDgZRzq8W8hHQo/ei
2dTXxZoNWkVxMqnHYVbAwhsGih2vJYZQ/EwdP1Qz35rqEzhf5i4PfEaZ8KPkTn0L
sOlVMZ752gIc9LQMGNCYELAP7pM4Sz4YbMdxnToySDBDuSoCplrX8y4m5YkuKgYR
5YTDxyxFrX/svCicF5osKqNGhvZ9RCCS+L5guIdW9B87QrhC/X7mYtOQatRAkBfz
Bk3a3wPfkSDBoMFpcFX1w7FDzpjF/aAGsSTs181WP6mzcJkMYgsRrDZPvf0k03Nl
k/1osSvSvmVaBPpcAJpTXh1e3/F+cc9q7ZyC/vgkibMyQ3NOTJQhR8KSs45m2UaU
j/il+eIEY5yfP0fJ1PIS+P7bxlxuHp98SdB9JWwqVXXJTag8b3nUqFtTSaQXLGYi
WrYow8g7n9YUrwL9VUj7Wgc/BC08lw5dRv3hsGAvFZH3ZWhFbCrLb0PMLrNlCY0k
WP929LJQn2iu/EjhhRkK8KsJUxTK5BrYI/Ln6b+8KvWK8s0WAqXshXwYVhG9TUcA
5/IBvl18bb3AlcfMecles4+KRQi4qR86d86WbsZyBYUD5k9eYGUrKkwTuih+2ajg
1t6IArBvn0bgvZraiBvt97mKW5G2Z0h8Au1mpPPsKggQJbKKGgK7SfzjdL3aRfQT
novH4lOgS2C7OXr0hJ7FFAFhPpt7YgqtqBdGlmnQs7MxG1hwsPlV8PCfW1lt9oOy
/Goz2DSufH0i+/xDQkN4quad8Zw2Fr39RQhyzpY13yuZBLmEqewoswfGbg2NOi7Z
UCqyTJaI3rYSKUEgd5kh+U9PVvMcUUW7iDKZyGiPI6ApQYW0TydXVSkdIq6w2wmQ
GOq9qoCqPFN6T5GXa3u8p7iRimp9CfVC3Hid0Mnn8wmmhLJG0tyZ2Qln1tWuzFJl
OJIKEFEaPZ3RhzhaA3WCY1qYGADRgOybUtlTAyhT2pJ/Uwh3F21bJciP7+aLp2H+
ps2cTlIfU6oq79V5KUv4AeEdjwwNHMClwiUO7LeQpbIKYOWhSbzsR412BLEkldoi
WyiMNK1YNpu1WHZ5SCfzXhIbLi60U5ZHyv2DKb/f9qmyi0le8LKJbIvAxLnlnEDA
iqRy/jrJForXCbNjx8otwjvoVvtFbmUdbQg4oCaTFoqDgZ8nMln/ewZV9H1Kj01Z
Il2MnjzaOFzlhj0YNCaOkm09ntXWiyHTEUI7DUDwG32CDXJUo68YxZ42zOOPhDuq
jTAVcnWs6johzqGQtsixe9nsT0xsMnrRbSp47qSNs9kT3V+hgAHJXryYCLxTzdH2
ZEiApTGb1AJVV60kjsrO6LCwA2H3r9/RiBbRLwauDXwGlKgn12gFsZuihyXviEb4
m5XlkJnzylnG9/BeKnpAdfwNAcgaf/qsLugeR8vWXoT3wIwRq10opjjQTKKgqWaq
LBl00jG8e2Anp+JWZS6+KpfABYkcAJ2lktIbAIJHeRxuBNClo+GNibFbbtVcl95Z
11bitTqkXgYwL8RPqpATJWkCZFlti3TbDvro1W0o11MsMdETJ+iq50NSrsd42Sah
7gobhRCuZ/aHoirGWq4tzUEK9EAo3zp79pv4yL3AP5pdFCiM0KgzmxSPKaw3R3nU
YKENCWortFCKNARjTQUzKfhkHl4GCZklm9pX3mVD6jI/y/oNEOfajGdhUG7xX/5r
BYpU3OKHuJSUcEUZel5k3FT/gWebPIwWxQMWG0pxMK9lCOiDQ3mPO1wALd6h/zCK
WB3AigKUlb0zo6cCTWvU1ovTOVVsZqmXVxcKwy6z47nNiuwHCKcYnnUcAcvLBjus
DZFxDLRXB3Vdh8k5UwgjQODNduDHO+O4/odXO70aUXgrHZKLIlZ94PJGfSV23K/n
x/tMcsdukjhp3+NvFbarpYje4jXgL/RdK7e0mNmES179dGghnEUmLyRuzqpSpIqf
2synwhs82RSmctWNOWuZu/qp5HdrHEaFyk2ecifA+7ViM7HF46MufyB0YbqolOej
xr9LYJBpKrgQhGDsUkuP1oEwDspxlnIqdyJ3yfpFB5cM/LS72VV+xRPRbu/Hll14
xfZwEXkJfeW+Bav1fdOYpVjH4rD34lKwFkPs7LKfKCFxkXX5TylvAKfjuzo39+9R
OTYA7JDclXm8SNwWVywLD5jpuFXZa6Rm2PGLolmXjw2rgY1OnshwCO3SQwBiqEFU
Ycr0+jm29BGJZyXVQtAqBOQ9IAElMCoaui27oe2ypDb849DNBI/nOZLyuVjpW7gu
cLn6lAFdv8Mw5oHG0i33jApFI9z0Y/ntTtIe+XbUpHsaE4qI1rlqe2MRivP9MNtO
hF71Lq2bxBE0q/WtkbTSN0GKo64XTrULUyXuubpc9b3w+nMjG9lQ0d3ckt7HB5wJ
LMq92/tZP1OzNelQpo8so9xFa/QXnqerygnc45FVTbhswn/SI7F5zKuRSlpO3awh
p37RU2LL+IQ2iHOeMEWNohQebGbrlYTVE2vJb8P0zIoXTyKdfV8U9d4VlPiaCHcj
3zIMwHd3YOYBa2VqQMHZCuufAQYIGeYMOu/F4DijK2qXec/vWLfLkDqFAAXhXtRs
XRFDPQgShoRQClyCmyc2c/r1SRxlCAUsXHDW6tGTsU6TvYrGrRpIYTB7f0RMydEk
QRmfx1J+oH79qxwlsoIPW3o82yubaU3usXEyS4VW0HRcREudYCIftK1KHKsdOu+q
1VjTBjbPJjx9JiixgvdxpvT2KyE6BjW7Xx83D43bl+pTv+mTk/Gh9RI1zHjz5DnY
Xc+MqQQzu32OfRVz1Vv4gX7syalgD/GbNWNdXGLUg1+aSxsofBj6BlnJkuVRUdWV
CRlH9J7GGLom2Zr65KejRDfPj/Xh19J0nWDTbOAvmFwufG7zyCd7bo0WOvAAUjOA
/GdHoT7XkBF9ILkP8800e7y+woaXxWAmSG5KQJZx0llVnQ8FXPPPKW8s5YHL7Zdg
GIjM72X0rj91ioREPUj5C+E/n55JdhCVTpfnfp7t/vFITAOI34SsVlT8DSY3F+JK
c/K2Z/l25XDbSF77wdYZeiTwGLKMwZKqcFntLrSipZYvp5jPSmt5vq+YQ4mOUD07
QgC3WGDYf4ffrnflPumdxj4R48qotB+jrZ0hE45NJD7wez9kV61BUaRKqtz/je+G
q1yLWsoXnsI7WSUNQ7bayoXWTzi8Nn3C9q/w5KSiKzzkw7xDxbIuhArwDOa3QgAo
187OJiDvhikwCP2JEX3Oocvm9OLMHSlw9OjWW7ghFXCynnhlXzt6s/BF5JtyenuD
7cpCoYXw49so95bNKgcvlfC+5Dy6Cgj1j44jIWauBkZUF05RKA56OngcxHhdXD4m
HSjn/lmhmtN20hOji9/A+mxBgbuW+AfzpHflP6VGgrRP3TY99dWGrhvs+qMYkrCW
jBl9BEp2i9uCPu362QZPIEWtCoH5Bmt6k9/VrWBMaG42pZuRfqJFhQ56rgqP2nrf
dNaoMGhZm2/dn9iG/lbonUC1OyiS+fhhZbsA5Zlr+nFi1eG9lGsILvxlf3xaGDh5
V2HDqsBMyPa49lm/RIdmwUaqIwTrqnBxUQc5FFPxz5eo+ZqZurN52TeMuXlooK6w
lQM3f7F5LunMJMkdRIR9hEy9j1ZoFhikjbkZZ1ccnOMwp8/Y6kaqR4yBWUlIrCDR
MTa6dIw0uNmXuoe+VQ3cbCxfBfqqYSj4iBRLyrCVZkdsUEcECiMeNj4S3AHzZipU
iibjrh/TL22gdDKWjWxAeEXm8gwvgRCOghAey4FLkQjuJenkUMYyz8XkUXB4Xrbb
q+h/j/qF3Nk3PrB5WkWf/E2eg4G86bTNSC4sspNPGV82RcF516ASbhFRxV7Z1l9G
D3gl3Bo9hSai/zwyPmmmIfrlxQvvm1laW4B5yIvBn1oKuqHj+zPzlxTnOFdzHeR0
Z4ds1CEXeNTvDHKiX11kknWzy38tXMV8lSMZFQzPT0FCc+5LJXaUu1XRwcpN9cg3
49yZivepoMqcUljDxp6DLCO+OGo+5nyPqaeGdsr9wKAAneaCK7X7Qd4MnzfTaKnr
3cVbWdDZxKhuRQQQAWtz6LFMydQHIQFxBhrogBzlZ5F12YJ11K3I6umaqOBbhQtu
RvXzS/6yz62Ui5YbGPHCIh3e1ryqIqi6RPj4RWQcpvUje0aLZggf+CsxPcz1wZx3
3G6B+LOvH8fswHgD4C8Q+ufIiqwDRHW3Hx9/i407YobH34nG+hOQLbRmbxAnQ2LL
k3743xf2BXHHEBRtgqVqlxNhhSTsFzTSaZJ2KHVoLjhxnWAul3fT9tkdq7+SqRon
sKK6Ac+ARu5EbZndvTZ5te/mwx0yixCqnhvc2evizsOwG1X4mId6WUTZlDSCBa+Y
8MOcRC1I2lBL3320uaB6IYOMfW0zgWfjA+s2z1tLj8YGUzAHc7A4+Q6rVOX8HRTn
2HjU8716v48umed/g9gaVjseucv2rbAdHbd2hcNk05xDVNGUHqgkjcJZnVG6uLld
jwrHg4WN0n+8oN1o50xCVJi3cyecg5aha12SwN7X8kts2DRoTib6OxyqbQ1ZE+Rp
pXrxREYa8JOakJewXxlbNkccgwrlefonnUe34P9tlReHhkv2xxkrUAgNfbteehnh
NVKZy6jKqRoiZPUUslLwfAfkA/4Y5q+svsc98mwzgfl6JWOAAJlV9u8/QgPmKnr4
TqPsnJAssstnnxcMd8QQxn06qy+bvXVMW1WcvIPVukRTzt2tuHIdiX34u+BgNJUf
pgqT3LkKpe83AWtQfOotCEhnmkzNNvr0f611krCCJancPiiCweK+pa9eYXHkcp0Q
up4l40k0LP1Z/D+fc/EwnPhC8u+RyNjy8vByxeUWJFj1qUWj2gleEFKOf+xmTil2
quE+QqRXXjbYiEnWUIy1klBrXUqUab4oCDVl9CoqsC1diiTK/P02Zz4s+MDdVu7o
TfhO67uZvgchRpKotpeM3VYJnY18HxbgCuTxDZ6JMRk7YiMYcoquC+by/LH69gj4
Cq1l+cMkJm9OUYJOsZZVaDq1i3CNrLvwfRaIBYWqvGgSsbuZ/hu6TehxP9I97uwH
7bukVzxZaQdr6CkENfw8Ec5X+d0Ck1jWbjOK6R1KyYAfd8FaFboE1QT3If1dTSVP
q4brewRG+7E1GgqllpEFJYLI7bl0hBTk9+SVrRMLwpvdTzvQ266oM1z9D+/CLoWJ
4RcjiTmp4Mg+XRctnrUinscAHXT9qJldFf/PPltQSxAOiMJswe+44n6vtnvlnetw
30dtrUENJFiMlAA1/QmS2/+q7OPZFXcbD7DPZcW5v9+PBOR1iPgkJBHq8gYshm2o
SH+xsu34ZcLOz7dsjw/rnFGIt0fTpY7OS/E8ngFnUQalVfISz87+K5liitLqHQmk
CdZl5WbIvUU7Xp7nbZZUOjZWRhO9DCItWVZfognbZqjKWPcX0lDV9eTOXxhDbPiC
ZLh8aU0uDQzGGge7jNYhp3wzwJ1D50XANcnyWkvkrqOUcKcSszmS0jmnvfA4JhOl
NabWkijl7kAGIvS+JGq+fFNw1sBhU2VNOL78AJyyuE9wNT6FDeV40wcV80CA0c8g
Ey2Ote9jifKYB+i12JcpvboQ9HMqNIatRlbMu1P4TZasP0gUZJ9w7R/kCYwq363Q
FWCcHoarh0vnro0XNM5nSxG6YY75ydmCz5Hjy65+1fEzmYULXFeR1BCo+hqOPEyP
NC8qJ0qT1XbiqdIUXF6xS6f8t+rpDm4t3YlHdGY5mvJzxQo8xCB1/dswmhfFxTGJ
UlOid6I8zrg5Jz4x7iqlZYIST4SRxNisBmFqeesUYt4JRd2INL+EVZrE27R+l+d+
qyhULKQU+XUnTIcJG1kNGaAkRykK0ItzjwuRtbBbaxLmlqSzqA28MpSF1s2f+Veh
yxRzvcZdoG1ftuC4x4JO1591WoGMWLMvQsIVcBRKkRAS6UU/LkGun2ahhDnVt2Mh
TzBXjqLo4Bcd6v5woM8efGk3hXlMhhBxSdMyJBVKUpqbguM1awAp1jv+qY0+uZb0
Z7ev2ur77oCFJhs/9YiaHAnAnQYxhlbJF/TYdq5pq0pATdmHsIw2KgmCmqSQtvx1
NH8gTPBL56JnrBMNWehaUpWlX/ES1w+hFn5LNjh2520swuV2377PVuDNkqpsKuSQ
Iv78Dkrm/Vc7T4lcajMO2+HipHjgbDSBNYLj9YbS6YnIaxr+98FMuEJCW1p/EeHX
VaYML3LkPdo8F6e4Knc+kfy+WlpJVybpTAgamr/vE8+9YWObHwOZYGaPLKJiaEER
QHV2Id0mMWDM2Nr64SP+8W76d1itkB9QkEgNiu5tqTOb/wyU2CS2f71SHj1jtGCO
g8ZHR57mJCudL15evqynaT8huXObWF/vFYag3KCqO63cVRECDnUS5iS4ZWuc26+g
58g+K2JN0FohHX5qpglW3DN4Zx65ee0pmT6bW4lKMhBSetKaLvQxOOTKXOWPQax/
AyeJgbHPc6JQXtlWNdDkrVPTWruaNwpARTczXxgKeKI9puIvH+XHlWZc2+Z5EbCu
ANXlGCdwybayb+neum+StwXEgVpvdGul3FUZwOpCKEDjJrfWhPcl+FqjMNcJudnS
9SM0FjYpiSsKzA58vvbA8TOiRCGLFyIKQwmi1FjWI5MzqqjigeD1EPGI/1SU6KlL
PQxFEG7IaFek8cEXEy+f7KqzI1slmxX8qgxdf5M9LbSakfHvLGXoUiWnheSWwktj
PQdN8G+V12qULhM4a18mKftkMGE4q01KnBbdHZChga4nW678J/k9LUhUVAyOUuyd
ZuXznu+hNwTphk0gDtpSVrgm2ydmRQEcqEZ1rZU37UC8Mi9/44l+tHZaHKHM0MIW
QW5SLAadporCJG8GvcTXOUh3IiKE5XgZi/IEGdL8yoVsD6/B5Nry3qkzK1+owfEq
K2uKVYq6ubHndFityNfUq2h8cD+DUvMNZ0D8zUwL1aJYp5MjprKmQZNgOxZ3hs4Z
e9P2KsGHGcyCLc/Stw+0fRZQ60Sk8Ptlk723jkResANKQ67S7sL73nJzMP0PvYjj
8G0CyXVims9nh26pDofXk8bDyFBzo1tOU4pswPnWPR0utAaYx3QVxGYF2mhvi+Vx
PmRdA5008TW+3N/5Y77NrTNV26VsGn7/a6D7tFgqH9aICJZvLfFGE3jkJLeq3n69
pfLirZfY7cLujlXuyKNPVYAKLI8R0pL2Ri9FbftEwlwZw4MEQBZvd1DdhRNYZ/TV
oPyikfGcQjW6aHFzf3XsEDbE4AWk2tkFONXAnIfNhbXJSrq34B9l+z6FVesLfauD
oZfno3v2ARu+ggmzGpfZOCoOQEd2AAY3N6h9l2qusYyZyce30UCBsVDrtVHquMU3
IuNc904l5sqmxg0F0n9SyN6GliGzT8m6e46EY+oYQDU1Gj3SkP/RkUXKoFAb5JtH
zXZe56fXNnTgIPu5iL27ufxj8PAwHLucsUwGAp1q4/pFAJQMPKva5R4jadeiym2w
YpyZG8VTHywwPPX8usoVL+kNFa5K3o5LJaF6QDQUkT3zM8C54U+LG+qrJtpcuJVc
pbU1SVm5sH5sPee3a1R9vLWv7HCzh7lD2p86IX6/Zr4m97iQsqmyBoXxtrRAqHuk
6acIvNk7TRuO37Z9Ur3i1S1fWxYuKwfHM25K0OLRyestcz0bt4pA4UU+UQJK3wMd
+5YJj6oExJ21P4019PM3ZCObou+ixGCl20ANYwbKvMkH76ocdSXR4H5sMx9I5KJT
8+VDu22IBBo8vjXgEk/xgEv0GVa1JJ2+uPJPTeCF0LevOa+NYg87iwCADKlIHlDV
uzSfSEswHl0uQoWMzAwcz3tUbumhb1y0WjcAmK9kX3ksnQ+FLtDhdMZJE2euI3zZ
WuZHEgnKJhK6QI/6rCOK42/ZbmIluFLImjV8LQnkTv1bsDZQtyRR8du44i7Tb8W8
NTw8DXkpDiCtxHCUWuF9Nl7mpQqVFbOfvEwhhWJ2n+KckSYPFasC/eR4NbX3pQjy
f5VyUrBBtHCGQ2K+UTmD5SKc6bjRqTn/MzbfWLyDmTU9lzRdYxL/bvLUPYViyBFU
C73xV8iDt+oWQuXZzA4Vg6qr4C22NglolDLHZ/7hte2Z+BR4ybu8N8WL+8pzFSlT
GYzZ9a7VHAUBpkF7JrSvtAGGe8zCBOXwVKdZJjrTFPSXwfzoyopqMT9hb205f/vw
ei/3Hw1o0lEgNPN4FHsRoyoAyH2zrtDqEjY7Z3aHo4b9WO4+bL8UkW2qcdMwKceQ
XNFgrXVNfl3gJz71tb9jPmPg1MdG6VFkyDr5G61S5n0NLSd1U7FAvXzSr9azZKlr
ozy/Ker/O5TWi1rQE1+uVTQFNJ8QxvMnxcx5nvPtMt3SSTF/9Sp/0fL0XZmnovDI
kvu43YVxHFqitRa7HYblu7AtDh7rhEl6pJSPpbGBeV6uzm14K0c0q22MTvyMTx71
C2dPIP4VLyu3O6/m6Csdalnh7QeffxopfCLzAJF/ABpWvE0XdKNKVBt+JdAJ40qB
wUZpuk+hWa0PUQYHk+ZJVGotws4uUY9sehb8XmsUhvYFS5sDOnks59AFlKMvheEO
h7IiokHHxclKH6xAPqkuBJQASLEbql4MXCyZYi0ENdrvMwkst9WrXoZvQVE6+EYB
jueXx20aPNLOPgUJ8mv04Ypgs1k70IQRun1BLbOsXw/IOL0Zgwhi7a3iQLFWY4aJ
qcLmbZW7iBvHoGcUCSPtCxhDoNAgR1Mx/rIKMcv56gm02WUqrBirNicztxSIfVJh
jFP9lV5EzKgC55PFgQJjujUqGw57bL2t6jl+iwy4snj9EkJtuOMvJJy0GYxXwWqD
jQtxjD91NSJPYQfdYLdt5UPttgB+YR6JZx6IqYrTuSWvag+tGCd9/Hqc0K8X6cyf
ABEIakrP61HJiNf7lmKe/EH8zVaOnIrOc+VXfgwgDXp8TpB002+06vfq9GpMNPum
zBTe7RfeGYPw2/YZmiekTk94UA1pxTbxOtmnBtsrPW/tP18fFqrzKNlGth/pniLP
+ZJGrgVHqupuq/7Jp8UWrk5S26dnOHfG8LO4f7XaH1EDOGHWD+ZZP5E32bPTfFnR
G84SKppk1HKlq2hQV+rtgQH7gsL7F3YvdKQe1Dfk66YjGJojsRZdIio0ua9NW3AW
4QsH8NWSHClLKEBGF323rnmj/fccoWS5a/TWEV+A69TCVBs8cYSUQdjpEKJYKEX8
LC7PFsI3LfAEkohKP3Potw3m75qY+Mm4Uy5BySa543DdWAZYTdWVtkc92rhNiFTx
e5esNliUxbidwT7a6iY/1MIUEY0mEq/FbGRaC/rcwVxPiqNlOfAP2T6et4wpgRhP
ngj0HHGW0Gmn6z21pdqz0rWKxq1xhozabiPrR4suH3b0IsnRUr8mK/osXYYAONWV
uID6YC83g2/f3KAVRSxQ+lC0NUBWYYzCPIrdCBZ9xssJ9qmEQ0sJL7TbZ7ZsHndA
J0eTiUJc/GjD4mSlHcBZZjN6ISe3R1iIo7UFthcv2Ij9kazTMiKtfVyytjBFO68m
9y4lkhDWclxcYuQKS/RR+djaBD31oimxOZWbjHhHCuuNQoazr73GaK1dkrqOJb4s
Lzb+jlRRPVrMGrAifKei8vCSqCQ+aeX6q5XbTCiIA9//SZs2fH2WqeN/TgY6gAiq
FRVx1knOX+ppmMLhXwqRqm2bmN+Tds2AhSnApuK0HC5UgJDvmqLrU3261z56vjjX
5BIm+MTnQ/BCpuqhbMGo24Nsd5EuIuqOigT4oQ0SogJ3yZQE3gwRCl1Sh7pOQkTl
Q2+mWQz3toP+yNt9F4aPPO01RJ12SK8rDCnCUTg8vdHj03gqINHQY0fCc9J4MZvH
D8MkynP6s9kv/gWf7I9cIGs4QpVQFqlBmlpPIodLz6KreZgsTwDi8k48yNxgYhNd
8qXGLD4fExeeUmnyiTz28NXliq/WVu+o4fLtveyPaWgqWadJgxqUFabllS2hmnU6
9D4+iuu2hEeWXjewDWVOcc73KOv2tkzYWMFVx8U7EDUU6UI4Id+clRe78Ad36c38
xef1CgYdl4S3gDB+S8m+H9trwE4GUiDbn7Wwvr1zrrKyuztGyjL0V5a19I1qbcy+
v+4H/DgumKQfHXZ0wu/Tw33NNSOxlqlmaNG9R91fnHXgBOitZgJos2KWSCQqkYP+
t3OC/DHwHH2Q7JAMYHu0W0hpqhlH+zfuhYodBGFa64zXIA+Y3ZiYVyJyFFx/hq7l
GFGrnMgSHvKttTOXBK+bevLtx7cqCMmVeUC3ykVxoS2JUiA/feL96NweJkbhVObK
CFVTfeI3EZdJav8L2hnI40ZCxSr/PV0BuE2XElgasTxQJZp+yGInI30Uqk4K4YhZ
uhnBjP/nlxUFhXwDjN1mP4LqNULE54N+Ryh24rZdX23zZJ5hwjeDWFFQ1rAjYzo/
gn3VrdQmVg2obLmjex04y8gYRy7Y1k5/54wuzLOPAELCDPph3p/Ud98MGXGT1ocZ
Ui4+9alFYAHlIfDr9y1CN8Vix06wDjP7DDecXQVsfXjTL60BF8B9AxD+7UzTH86o
UqJrRXKLtbONaEjM2EqAFY15DAf5uTTGurkBOBrs03Hx68GODUJeImtG0/hobcIf
FvCGGWm8mg5uv2QVXVXtWVAUpL/409rMSvpSjm57x9akuzk3fb7aPi5CEz+9ai6u
pX5unDElC4Eecuwq1kjAk2cKevtYV5AwZ7ZBn3OuLJYymZlTsVRZTZY+LgIFGJzT
3AZKXEAobHT28/139DaR32eCGq9YK5DEZLTjdikndgmLUpP056xkI28Yff+5dZTk
ODLLGtTdd5CdXPy3xZ2VkN8EHRFzi4IlOUhTWtHnvEuEEx7McPxqCBu8nF0kpolo
Nmm84iGncNRLpxTtigQpgLfAe61glQpvLLLM75HArcW8tq2VHHvPlsMVTrQouW0g
Uu1NBsjTCW8j0ke/Zl0G/QDC21Qbdj8KwGAPDq6kZG3J9zzh/Oq9qsLc3M2rZLtP
lkAuyW+rfqeCqOEU5+ZQS79pnfoR2j1Vf8P6oHVGYClUYftC4zlQ6qEc1AUMVoJy
xUR/v3k4N0pT9G5ECAZDLDqcsY1TsBBlkMIX0Tlyw//UU9dNREcawnC+AVj5f2q8
hH4qMl//JHwx8e/fGLmA3WGX+8Ub5EptmAnTCgHUoKS1HJHVLSw2DEdSl2fqW8eg
CYVXYmD9atcP0PHyVl5/6/M4XSgHGSrp0vjcXncfsPNLz/AGsHpXnMCpBDlTSg/I
qSXgWi7kcbfurTqLWVXL7C3wYZ5hE4STGxM4eLZGXyITAzTcrILRQtSJKcYYleKS
jHnF+JOQjjNAWXNCRUnQcbUzmq5I2tNSW5WH0ePYUFUj4O0jjBWvodoiPV11eB+P
2hV0orWa8aWKdSjePC+zqErcJhpvffOYNJaN/Lxj2SSnuoomcUGOoxq13BKeMo1p
BiRfGrDawIWNHwGhf13xFm2DA2sEKxCXb9cT2SqzB1EGd+bNZyNIa1vy42q1Tliv
jHnJOdujXSOTTw9URSFuO2f6C260P8f9sL73QflSzDSs3KO/E93wYeYd9bbzqIv8
ibCS/FY9BPNvqEhjlB9LFWqVejMg4p08NsKGQ8AJwf8xvWhprX79NKKYq0nO7ynD
KdKkxK7ic4L7YpcE+bYscnaoMVwkvOHf/yJlCPz1vDVZ1olywn8L7ktghgGqlXSu
7ERe1803tXK9S1pINk3xtzauVYIHqmNvr55rTg8/wnwl3fFxv2+rQbSLzsvz4CYf
F3IRR7t8ujQn32lknYTpseulAgDmCx36OFGFNPQnIDX8tRWP2msdQHRQZ0gEBP9R
no/KZ35bbndqAEc6rYNbT3UDy4KLotDLW1FFfwSRbMejY9DQut8avNowlz0pBYo0
ySoAGuTEvdt0mYol9nyCu/5ddkRttikXNiOYE8u3I5D3N1V/hri8Zkxv+BsrSI3+
kduxganqm4nlS/dqPAPx9I8eguV4C4lv8zxbgn0n9OghHbveaUeVxVmZXSxNdTLs
TnpsG0gNeUIrTSGAA/u0LwW/muDT6gcjSO6sg2po6YWX9ZQMV/UiF+lx8sL72WN0
pD9pTzkdiFJDlSL3tbxfgfJT4fdCqcEb3wXnaQvCrZEy5hXVu5U6k8eENsw5NEYE
DZ1SX6JuEokRapp+yoNnqhlSjap5UA0XcbYh1ePRIO7CdDd3+I5tw/QfeZb45Ysz
Xfh9XD+4vPU1BwDAGV416wLpWAicbOSmxPovKrrawzbI/pWd4azm4U47nM+rfO2N
4YDWyHqMw3YxW+UnjrB3EgN5tENzkVRmqjxB8LxXo655sR4WoGOOMvXWi9rjBNKv
NrZCRDnuX4oLJ2ie9LqJiMhcmPa09d1vklwPm7Gw6hUk9VY/a1zFh9q1IDHO/ty4
kO4TZ33MpaZ21eia5Q4VvbrMBEf8tYphJ9g0TM+HfHxTMgfx0pxuknU7Xd55H+Lf
nsG0ZAqJ/kaW4wvgTLuyG8j9s/2a9FIGT7cbbk3Ihmg/qW1drzyie/KkwXDt0BjS
O/V7gIR/QLmc3SvO7poW5Tkg5gvN+DoyPeoJFyCDBm9/wWyvDN7Z0q0lC4xy6x2H
jMt7GVT1AtvmS4tPkAW5PkRZ9qEwFnCZ0+syVGExlcbJGS7QfOq2MFihhKzIL7PP
r+fX3aUrVN84Gh5xtxtW7xqDkkkUxzUis6QASHBSszGEf+ngrOz5G4CAVNeekHHP
cNcb4h2EZzTXqX4bwU4V4KAKBJG2GJWtjxxIanQX6TLDsHHFb8452z83owjQyeEE
s55WD6UXBUlXBlq3I06YkrKpIb1f5PA0TP/PA8VfFfJDHHlUZnzFKabboSwK4Nqs
Evjp3cRot7nRUEF82d+0l4+EqkT/tax/Iuql98lkuHVRjp1BsBBEg6qrho74EZow
a4PcBIZTr9AL1QigEzzCndlQPZjh3xUrOPjlueduRcsM3Nk/uwqiomj+Llu5lIOM
4y3r8sQk0vbOkbYtwccKN5VEmcjfpE8W4++zxjaXokD5FDdbXuARQcJlIqkf2TNy
3UKs63DP6TxPZVSgN1nmyLc/DY0cv3oZIjjukQ0SCd+F/Ac8BLNXDX6fQSobql4n
EKKVeH/IcTegNxOTjr4OXb02SdHNQS56rVapmGq8ostBYQwMuF2Zi6byDDkE0OZb
BN5tztb941bohgKs9MDA+p2sVr8EaoFptrO1xbrJKY0oOxwOjuM1SxAgkFsQF4MV
w0UdncbP3dYmf5Ad7Z1qVvWzSh13OwJqo0SdMsRWOXB6fgvsRmfMta7gxEbpbe2c
ZifK5bRNjh52t2AhZy0vN+PJL2MCDJ5iczUIKhDqzFEodmYIT8wuW9kIgbFrzdT2
KBLIM199lnMBIgcbD9tOjZ59foKtanFQ6cQ8IYOb34KxRLqjVtUL7gpFsNGWFlVj
PT++mCthrwDWmjux7L7y0fRrt8nuVVjACE0LqyP2YkZj5u8br4u/9uIMtrAthcix
FZ7j4T5Lxy5HSQurdMWJ77kYp0ubPvW2kX7BIopXSbCdCxWw+zXmnQu9K2Tr8Psw
vGCSXuwHWmoVVT10teZJmE3mHePpjo23bOmDmkmzEqU7cwKiKhu3WdA80Y+rNwOs
3yidbLOa3fukVJBj0VPNMkz/5+2ZwYJ4wPDQ5YwYcMHdgM6VI/qV+tiE/xMs5Q5E
A049/T3MCcgV34tgBSIDaGwixQybY9R5es+CN1vQ46yFZz/QFJYHGHXrqWAqYXvC
Z3vgrWFRSRX4KYT6LuvyeExxYz8Qn8fMBVFPKZiTovzrScb36bupw/4BA8UEYxZX
skg4vEFGexNd/M1kFF5gcgnalxSJcUR6e1ewfqypIvju17NefMZKM8NrPVaE8gKY
OqYLBkL7BKqOmslh/IAiDop2LsUqQHeQpbVFrIUYZJA7YZf//68g9Vrfic3FOuvY
ziRSl8byqFJqIdubKBakJCGzEnvU9dtuQ5PWD6TinYGn+GyQyN41IikvfJGzc5IC
pIHnR9e17iXQ8e0radtOzfJUUOxPY4cSJ7yvajiXziwzfR/WFrNplW0Zpikf3S/L
GwoOOZtvFuuhH1/DXQdeUhtxZkE3NufT26j9a8Yl4riIbvB2XytmgUmmyutyLMvZ
YYZZ1spZcAeSqAUXqSYTsvdisFUEdUulI2vMTPaxuS+uW7TBGvGPWs+W4uHdTEkD
uUyRi0+NoZzO9nbw4abaRoUop3cx55aFdaCztsGM9xejDq+ZYpfeUrHYMtiB7zoF
izzuM/NTVWibDrrKAJ1/aKay1/WI0WjJh0v4wyv3C5aYjwLhgdS/HEhMwqWl04kg
N+A6fhMo+JqXl1H/nVJ0nhUGXfSsN4E0mJSRQcfJ+mSqGZCxi27cztMCpJfpXM3Y
O8V52KvBU6DwsqmzHM+FmqxDfmqTnx2MadEvFoKt/ezNjeTY8b9uXVdtklshwZof
mX+Pp+Z9FO5e9udBtBz5ogZ1elUwg8cy9ejSN3NWBVWXdHaE42SV3lfN8ivVen8Y
sD6GQqTPEWnrvIi4jxNy3Us+oeS4d4abxncQNIk0a2y2NIKWbnhfaaLP55ItnsWo
zsY/RJr25s6y+j0KbIsCHK4DiA1/9rOKRJ0S+VjdHtSd2ZMKzOZLnXn0dSmLfmZ0
IXHAK7rBi5LFlu2ARsXeSRU7Zz1OSLCBO7/TkEMe2+WVU+CfYp1aJC6OKCBedHwO
s8F7VtzHnUVcDrrkzV05hJJXvX4NZNgdXBrLj/JfybIUarncLSzuKEdvSuL3pG9g
wjkvs6XqDQ1BsX3R/znGgEynYnii+aRALzvURls3f107D+Lvst6/FbdGUsWeVQvY
M4stMVvrnqYP25BClDyqrBq0JFnS7qGdmIKx+lJWYwr97Bxs/t999aRQlWDAnE0R
bf7ZBQbwn+A1l3KZXJIV9hU61xyPQ6AwsLDuIYGHVV7JMBfQPVGOwAr4ZmCzsW1O
Ws8aSgxq7I7iNTP1smzqf6NBtYHmL9wdQThdAk9Y1yb/H6BaTDRgYQ/BNzt5/eeJ
T4gdqxiR6liQLjHJLNrkOvxwXJTqO8NChAWnCzJp+IlEILyqHZbQth8dNGTa4HtU
l9OwuqEX11aXTl2iD78R5DtZ0EV3DEKwIDkZloCcooszh80eNT1WQ0rbLwCJH0yK
UdaZPL5q7HOFU2Tpy3OgOvPjQ1jUXOfw0ANKuexIC2K0qffeuC/W0GjE8VbaxiJk
feJZDdPgxwA2iiaFV60rBfKaCzBWCxqn+l4L4kvrr+9sBFrOOMC2GA+/kJ5R1lXm
crsq+fgcG0CXLn94eBJAkrPUxRlTDdZqnF8VStvbHwRQEf7fwv6ZlBdvdnIhFHQZ
S0OMUnwjRWVy1lunu/s2L6yqQgj9hYUuc4h4UAS9xTMtzUdBnNTXH7Ao7A/wXIK6
pXGqPlHC69dA8csTMVGAl1I/YaFDYOwFo52iBQLwa3jPu+XuyvicIc1U71VaN7XB
ENINdMLtKInvaVmDib/GY/c1xJdNvOWkSRRLpdMUruDvDomhnU3z/DtWD5GH9lS5
WQsJzh2uiyThe5rhXU/oX3YywWXhS7tu338w19wcE+wlaHCkNG/4QJj0tFAVWbC8
OLNvyLp1JKu0dhc/py09CjrlFHOaGQ0KTRsOEJL3cSM7KlJb5xAiQN1A6KlxEKIM
CJlXzjRbgf3jOnwcXQvANWxOpRoDAxztGRajOcmmjV0GgYzWjiRmqVQ5PpNjksAk
KP7JLH01e1pBZ0n99QbE7qGFA0pPJsgEOlAN2TbjvsozrbttAcFM8ll5koaFK+F/
q7WOQRZSKar0NoSLpTGGy0T06FJGG2RTiPEILuq0xoIH8qrZgGpZHri3F46WFQAB
CEevCx3V0rZDHl/7w5zZnVwNLWetYQY1JC2nv4xLPBNVAyNHJUVAzr4Bjt0zaQXj
nKjF2IwFBCByVqI+xRQuQZrctsYxBRie0m4njBYAOL3aFBRIty2aHoZ8RXGw1rUQ
BO0wgZh3mDWCAiHTVIemehK5f5TI7lJGO2qyaKSH0qOTnLDxSY9l+eF0rzdidRBz
fB3WCH4F2Tc01fg6feMPHocf+eiFHqXRwt/fYT0stR1mXtPV61/aAthW3F5hvvBQ
KZYI563t5BwdE3G4tStKRLs9ECfFNFDXNKK9JLu5YjLEa/UW799mRn0Z+rfLwUV8
xi2ox6yuWeaeREwUca5ywRhg30NhJ/m4uC3KA2aB7kN4d8jrBCT6l+WqTqng/fJO
B4azncSFI0d8CWKveT4b8tuTc0tKZr6PIpgv2RLuQK4a5rrg2+qcC77hsBbwdnQw
JivW/7NEIRMVbHZ1+fTFRzfOdoURlR5FHbyG8HrY47t9DYaT0wKABJZmRQIk+21V
bW/T0Pbl5tMyF76VD5n5FHwv807por1neB7otjaf22FwKi6WemIgRAyqLvmcSWFD
PseEU7Nyhmsva/gvEypHI/Ed2fTpEODtDm9ecyGhkyTN0WGu7mI/70GLbz+szIuV
ZeN/pNBSJpKE0fO81wGQtDp1fP5F5w99yeYNafaJ6nve5HJF/46haAZbv+6vv65f
167A5Dym7kXFH3hjD5LbCNWuM0XZz/ZTt+2lH+Z9vaXDfxrb4Uk4ctyhWRX336zq
HbvdhMmir4B/NCREqVCf2zmUJQSKtMTBxLXGL6b32KiX6AKzsmSHoD7n6M/ZYEXV
q3nbMkvupHSgSGQVj4KJiGtjzEdD3xSdOGun7C8MXrzGYv/SMmnVeWAMkXitfor9
rzRf/FQG++Gv2uYs9ut8F9vPZZluMZTXo0/vHCqXt3xD6S8N8Oq/nAYeBWC4id/M
IMP0A3ZgIaX60htmaedYTSTEamOBSc6OGto/3Zf+J7DcFSrG0lg68uYIfh+ISj2J
RoAFQ23PcUvTr4BMJBcPwMRme91Xs5yvlZQwPO2f5uzo3woxa5ffhIEvlNQR+13N
qipixbBjbRBlJrzt0ttJc3tpGPwpxzP3mXYjicLIe20H2/JxVd+Vr8KfG9LK1cYW
upA+e9TSNZEMq+kHSfJF/ZYSz3gsaQP/isgcj4cEZmitrKG5fREen7t0AoN/jVx6
1D5nonNK9pI2czVkCMQ1ZOoPKIkJhHn9P4qnHAqN89FwRu4vsGZgBuPWp265Bx93
rMiilUCknjnwes/yC/thkZtUVGUnBDgKfjjB4dDPtBdrLNsctY+KTj7uYQ6cWPAL
WaXpnvCr+aGkmZXyvE02Eseu+O0YRaolVrnSvtsCCiUP+v7ndkC7ucnBawPkj0Om
9gJH8u9poCc3E4/tECZYi3vV1GueiFUpaD8eDVSdWEIXxo0Ermcpu1fJFr4MdGIE
BCbLOtqB2iqr3CCSh+Z9Gtno1hesuofM3FHqzEIpQg1ElakE9km1O2huw1ikvgUn
vsr8/kJgEXQ8eemo6Fqc3oyZXH23U+qIStg7psS5C9XVX9zeAp2shqN3h44qG+Lj
oEIqLAtg7QRJBG1+9v0N4hJGz3K6Qq5qwV+v1hPvl6CEpGjEGMEvzjGykqBxZjlj
XgDT1ZHuxzo/pR4mdcVGP6zcDY4lriLA7iUf2z8hPN0HeH5LqT3COSSVPIdvDdhN
pZ9MIbbPknsidQlZLmLNkfgNnD+Cbvu0shxKU4ZcvVKKvZ5YpljBHXqcGC503CrQ
VZuXhwbFYPt27WKpsspAioDZUQbWqKvQnZUn1sQAC8NGQ+wxWVk4EYOvF7xPxG4u
lZ8iRl3G9QVkFfAVv9fNUXVolbszAwq0E/IQCz1Oz3tq3k5wBuBI2irgptK6GHdh
w5lNyArwrgPr+timWQZy9HRQOViNmtDLDl4IePjU28cwq2l6SYwmUFNQwDJaqGOs
OKlIznMQmur8zn2mq/wUY1jjBB7t2+EFCZhpMgZ5Sh1Z2E4SGgJVXUz8OWRVd6ui
3TDZJL3eza9MINewAs7G4wvsnLyA/zlHYCeZeceIc9FrP8xQWgplKszoP6QFUiYy
+Vo/bX8bLRFaQP8nxY0s5arzF9w5cNX65yIopZROrWQtlVm4uxpWvowKaaz11iqd
A9Tkl42y2CjB0XENN09Ajl6c9qW/man8lRZJu1T0j4r/lYg0Eu9CAXJqIRAgZTOz
6HlphiPoV+5ujifouqO0+lH757Sv9pkQLnZuNY/rCenWprYxKD8fLY62aXcR6NoW
5wSGRehYZ5S4otHI44FZ5Ef2Shx6rIlhObUBWfSrWLBLfJd3z+0ZR5bUXisomzJg
I7tbkLPLTJGA5moqfS1yrc6NgX6TJiK1jHddEaxg2vTs9ASOiNiq0jfC0SG1LaZ7
0VMyCUhO6vBqG8ggHvnAwEOLbdcRhxjIEu1saSlbXNhhy/lP8TCWjFTUEergQQQd
RUS0OdU6gVyr4enpdjRWkF42ReMXDVocE8RqWWYnISmQH9OKfzjA2X26ygoOTBpA
64+VRXxeoXQGNuuvxY20F0krGYUIMkojxa346Euqx66yZpRP9YKKalWaDnBkEd2x
+z5ydVOBkmvlZ6ac85CGSBCycvIHHuQHdoLQ3jhCv4vPw/7dDlZKIcMWSzNL2ofv
l2Y3IeEhYJtDy31wegFumKEfK4jV5uKQ9JrIvYHIfcg0lELGPpmKP2M/ihxQ749F
poQRqnNgL7R7rJ91sv+vzckbn1fJ148oppUCDerPwKKjIbGZT9gujqG3/Rvaniz2
bqnlbcAX/if0I6mTNcGRUUXGiPfrkXFfBYYF2Da/poKtVItARDicEn4iEbFLFLFl
N2NmFai08a75uCB2AoBN5idnbG+AWbqFdnwtRb46wzUq7Q7EskGcKnaeGYXmk+Sr
sMNjgqU03qRaIPMsIPOqixln8wAKVTZESavz0azU/LRSC7AT1HAX/S3Plse21T30
wNNL/z0DyZLmWdGprRs14Ecdwmj3RchpGy/SAxtHblhLoCRbOfge6LF3mUqGSQ3a
sjukatvdflVHLmaO/feyf9tjXO+VzumE4vA+LJrXtqI27+3/yyUpYJ/R+1jg7VJh
rla/Nve9ssupmxMokUfX+hV34WnmWlZlG5KvCD4wyu865Xgv+r7+jIiHbmDVKxn+
Nb5KvUmlIchwg5kGE1P+lHybGZfFJAfjBgocQpfxIicQzeaW1eEj6pgAOkuCuhz2
nEH6c7d4oIg3V7eabtuNYEa4VyehBdmuvgR9xdaLyk0gsv22mJSPzn9ae0GRe+Tu
hD/4b/bKgiyrdevkdLkhhYEIzMpfvrfBuLRf03yqwo6H+XADgZJxsIjLtpjwBe/S
SfFHE86tDIJQ1mirIq4tcWuWKuzTz3nKlNrGjImuRG2eh48ZmU8Ua//Ju6z7/eFC
DICbv5fxwg0YFkZsz3k7cXHTyGTk0xyQ0VzyOoPfpb3sPvqOaYJcAFU8dv57Ku+T
qeoyxuep3BO0Crb0iwaNHesAjySIJEkmPEF6izX5EFGoOAF+rMei0EKDPT9Tlp8A
C6o8g0KVS7BYJ+Prm2kJb0vY6J5xESL6s98xBbcRl9xMuxk/7tt2EIrDJsuGOG1Y
rDpNqeJYyiiC4+Ev4tOugfB+liZl+spbjve3CNs3eXqdoSCZT3S3d36ZKzhsl2o/
aVi+lcbq7h3fhy8pW3HssqP8DzqXDB3J4LvwGIs+Loao/Zz84aTkiYbG29w17Oeo
4biT95gX7JqZAiSWVe0BE9Dw9fZBb/c7LKhLkSyk3yXB/ps5uEiXYHyl/Vj9sM7v
91Rn/DthUR48LENsIPJsvTRIUheWG9EW1hTu8UpZcip0twFcMEKEYHEbLJwjIQEW
NGIGoSAYS8WBGQeLfZuZ0orSSUGWPOyfF6GYeJ3cLAYPAVc3KaraUVHVzP8whMrZ
kFW48qCyzzQiYCNJL3HbtPxR2S/Iusr2CSjOnJPATcn37CAa0d9+bcBwd6BKwBp/
xAWeYYRd7yndKc1BmqS5vj91pZRRfEFNz3XA92aXuFvYzdarXGxhegCBL4L+oHzE
CHn0wYVpwwMn8rCZfBlXH+gNBnrJJDjhwyd1Ax26QcWInHkupykKFVxqy60uBh9L
TjPdM1HZc4MVpBncwmVYdREC1DJDzoFHa/ZGQVHENJU9LnwF8hOiIl6SwsvN9aMq
q4usBCKSgMVzpTtqvSnpO7sRlUuhYv2GeuT7Vjh4BAVsASvuRDPkwnZuLtxzJyYW
6sxwMC2OxfitbqZZweRLuyY8Z+mpEzXFdBNoRi+yxhdyn+zclcuLUC4jRyD4O51j
Qa21nU+yb5hLcvfVTn49l41kucBW0GPNlkC2NmDER8ZaK4yHHzg8Ut+pnqyTuHrD
HHEr/3YMekF4T8KXp9b54gRkhQzbdRz00Tv0e8BoiKBt9UGAGwzrsotMv0FtpJ16
OoOVRPM9tlKF77zZ53+pW/Oa6AtKXbuLlB7cifajryWwSd7+0FcftjQfteMbjUQa
bOWk5gVeS1DyxGBCbFHv3geRZpnXdEcTJeTsFwk0rOmtGlKKZbtYNz2oVV8cNEeR
8jcCeuuRAIzLnU+q56cWHvwE++s0jUwDckGFC44V/If8d5FQZL1yPpOUXaNXa2Qw
cMiObNL+4lascNOayMhy7Vu3ayfAtmZn2Li2bNCYnagQKqB6/4TgE2972GZRohp/
2zbqw90pxuIKz58VcFosmDNYNdTAdQwtxXCFau+SaTnkxASPuIIHsFLQYJQhTmnL
PSZFUr1Bb70wAjPP6v+2LEKaPfyy8lK1N10mshIwPAGQiQNNARDWQbKsftQgcxE9
6a7Axl+W8JHsSfQOgWzkJT/a482qFL5qNhpqnY5dblT0Z5Rc+rZjCaNyA1mFwmaa
G3WJqsHQYYFue/7xRxA8yDJV9KUogC+0y3KXZJVP44YfDT22p3z2PK5QliMnC4al
UmB/Fw4PlBJT54KI8xbCx/WJeSf34GxRDGbIU2NecFwntE+1WHlS9v2E3W+jhp0o
jpxNQj1uONteYcafjejJXdxvq17fapIFU4GoblzVx4YJR9j+9YycRQf00xiONNfq
tcnKFMVTN8B5C8aFMDsr7EH2+WrsTTYWn8+lRpdMt8d4hmD9g/SRKToBo3dlXKAe
L1wGP/QUOzUiW8GtjMX+PRJhvcAqY6VTxhH/WgKKfG5mwqwSHud/O9X9M39dypHp
kzgAnMjrq7LyQO8HNgFmkkbIL/P8QSY+f2lyS3H769QiXBFN06P7yVSl+pYLuf+N
BPL3RCzLQbAr0I6k8NCiRD8D9WQZQTfn+SAGv49f8DHmPDv78ILl3olac8O3CBhx
iLYLvWzYyE7cAerrZlYsvL3aNmRfIfhFYMRpmRAUx8iSZIpsdd4JDMiUS9kX+QNc
dqzopYSeBfHX+Ib7ACINMsKz3wKXUQv+00Ew99YMjKLO3SWDdwjRE+OLksOLQGNn
JghcCUCl1/erL/0dzBEdyyr04kf916491p4L9hey1ZeUWmB9eK+Q0eAvd5hFQzUe
FRUo8f/IuDrhBBr+KcXuJ0IRKUsywqUuv/drzr3XWl7vMInNUzme/Y9gsn7JsUi9
FDbepVziSJ2Ko6yZLbOU2EuKtYHdWikrSU1gqFTOI3w+5bsg2CSNHDbbO8rutLsa
rnqtyUp1YsTCAUH7qVGhsCBm3/Kqh/aPAGKVZCblLlu+A5q93wk/V5x48IMran2A
2/grSy86GOAtqRzZTyJMIBBYN5e7ERjlL446HPVSWdQI4+2gHllYjL0WNnYlIWMx
aWDwbQD3yPNn2joZ2jAnJqV0hnatBaMEvSCHpFwBCv74Zihq5buD/aFBVUF031VF
p/G3Zx9pl6meUdVtbhZIEK/+8nSbYFkimveaclCKeH2fv/8sfoqdqyBiFUHC+lD+
GBhCG7JO7ZxcfKblVvR1zpXvRwfWTxrQi07tFDwsAesYp3XOkWxM8tI7ThTX8Zky
DuuTzDmFG7IXVN/MbJnzMTFu09sLg2qgmZX8IaCSmV3Dr/mwtWAQKjDnTWjCZKUW
8k8PW9VWMrZAHn+CqMVAX9T6gbe/i6q69uBQwsb1T35akfOsF6QZQ9rim0D4JCLM
szT4DtHmdcurvLhoUkUW+CqDBrxTACFSFxoBoX6U4QADsi+Rd0Evm7wQt3Bbu1z0
aClNyzLyhlgpAR9BM1k6mSea/7KByQm1OF4Jg4x9vXzABhwsCV+OV2/tgNrU4fN1
fN+7cqDIw07mYaDgaDFT0PifuXkvQ/tg01lr1NeORnnASAAOu/Jtr7YjHqaJksN1
CPt8kQ+5yBc1bT+tU7llSxKOehMc/trFs5RfUspZEec1XhdsD7bIwewyoV+hMFl0
jSuxetB0yM7obltjIhG9KatD+Gs18cMkNfF9chQeadEIUg2h0S476Ug3Y/4b5Y7N
wsi/Zn6cnE40+JgnH9m72wmXQhBv4fQM5S99Gfse71ohCY0lziWYqxiP5R5dUWhj
jgI7htHkVLZA2TzhebuszzuBgyh+GhxlM2DBXlIUTG395JxYoVNZ8rWMZNaWzmoj
C7G6a1hDCikw5SnYVbjEcmRsVcBgCBG6AFZpxmoADU2pBF9ptcqrsG6s72ulI/6z
wL/JRXQEDhC1bHFwXKMGRRo/vrEl2VUjFxbgZqYh/5bGoyh8+Et7IXMT6J8OMbHK
cssyip66ochkR+LWLBZOT3hXh2gsBdwF/D2UZYkdSkLeMk74gNK7rikSRgh8MpKt
073BPKZyGEZCjXI1k7Zci5jDvbwqhFCU2m19+aS8fbir/CY+F5ZMg6UqHnZLvGl4
OvQxkkCMOw7hQ/nx22x5nm2g+uge+C8M2p7GHLdllmiVoEtvHTI2YFMR74GhxoiT
UviAzHDH/K0YKadAhWQRHQ8tzlF9DC857864TquZrRo8D3UFIZBN0HF2ICBUiSg5
rPbT758UwP05yoRSnmH3OKLmIwPwmkvbKiz5I+WMMXl0ASuPIC+UXfM88dJiAV9g
2e69QFa9VehHFx7QoJ7LUJP++SG6hFwA55HB73gvTHruOJxMaj1PQ/9jYnotlc0Q
J5SETePA2PU3EeKhv0FP53c88ZmFbZ0KikPQR6P24OOjMLTx+Ey9ASPozTbV01xb
TKidBHupSFdIQYnftznDBlZ56Du6B6qRTQ/RupBNMDV6o89W+6imaDrDmBZ/BbAK
GBuarJ/I+Ar4/Ru/s/v+mANcnicAyi7sqnUnM6tIC+WDdKAIw7VFTR4Sru4Vi2eL
n5OODA+xPF80Ev3oS+EGsLMsbfDyb6Btzaj8+iKs7jLgvTaQaiI6ILJS5/n7kxLv
lc4zk4wUW+8877fVeX0rTkG+qVa1P0qmdlawLDZoN2I3zvHbQdVZei/C32RDx3/N
rieBr7lsEUAob+A13rEuwxh6foPlCSLK/riXdc2rGN9pQfmE9v7LWRx7QgWzIdoH
W2kn0luVTm1IQ2fxzb4mQG8zIvtoIFdiHScnQbdSAbKHEx7qq0MgtmYyAQNGIzcr
MTzZJol/PYONlQ0XfpyK9sFg0xnzzd1xQ5Gbdkeqvt7EkWS53KFNhh8vF4A7/1He
vg3F99WL9Yy5FtMfRZ3f98yHgKL9/vD9/50Z0ED3HmTM2AL2UCPFJF+ndWIK2Ehg
8osPYH4xEKNDxeklMqFqQFLwP1T88OueMhWgzY/vXGEqWSbvG+4TD4YuQmqG3tS0
h2Nqh78A3pMCj2wBJcA4U345Q8tAhXYiSEP1G57MMYQmZGOfmNcP/PXltY0t81DP
lJbT9LL7Q7WRSQCPQjCF8RL60gCkWB+65jUu5RePemzylEHBSR3WAAKfrCfj1A/Q
RxCMw7AYzWLbMQHfNpO6CrE1EfFFE76HgTd5+n3im7yiHMDniilSKOIqWDuCDfwL
jdifWEiAzgz+3YIMph+oHxLZpA1fGxq+IQ4wqi0zHVphDjGzH5kpPhk+ZrUT99AO
Kw73Ba38H7UZEsyTYRU4rZNcEsODL9gi+5R3FhYN4BBn9kYpFMklrf2rR6Ww8D2n
O/Fj0qXiDrzcWSAIsZpzF3MYWgkV/CMh9oV/FizAl3Q1jJkM/EA0hJ8Mei0hHD3B
n76T00zP+F8s6B6oE6yLviTGNueT+eWOekW6seFCZ44qMm+mZ0DQS7srGpIGKehz
H6nC19sKlqTgLFurFrnECB2tC8FTzeJkQkp05HZMp0FGcv2fofTdr7R9HaCFFpFy
p4iti1nCr64/NxEKXSd2+nC0YVGl2cCOpiDorLmHt0kIRQ4/5+xmy1GFw5Zd/NfM
Lfi1u3HsbUXYVXXRq1IQE9H+NhxtkliuoFxM685FnfRLLL86frmyQVBoVPe6sKZ8
HMYkgjXQBTlWauzIYNgwgc03vUXgQWdjNVloRAw2h1G60FHbCc9Ic9SMfFhaOt8L
KkwMezqTYr2C/oh2Y+o5yia73D2X+kX/rrqaPwuWBEpSkOsobjamDSDmijhOHI0u
NmwjDMmwGCFC2jhGqDD+fKHiyxzekDvUDyaEbAIXAq1obsaVoytdq1Z86+Qh2RWp
OHe6v9sU9YygodbRU41IIonVNbN/EJoKQCSzvNCj4vZqpM70hydP9QdwMzycbdPH
WvwiwG+gfounK+VK4OB+6mivC0rJFOAb0ObOjvlJcsCvd+LZRwQTpp/j29G9A2ma
PTfTkkXhNx7p/+oHWm81iYnUW6wjnkztlApuBJthMStWp2VdqTc+f4GO620+K+AJ
2/u5Hf9+H9DKI1enTv8g6qS1mP8WhYEW+I4ZmxtWb4FFd3/FhK2nTVrq+jpQw2J9
swpUzAcEqzx2VnLvOS+W0NGylSUZlO+77ja54yHaZAr8rxvcQ3KLmn2Wkb+QBj4Z
tRb/YBFnw3CIJF5xlkQMzUfOkZWdm9G8eXr3Rm0ey2rqHPWT66afrhYurq1+G3fn
fTL8NFEg/O80owv16AGk/h8b8YkQkT+TNCsKrDISZum4GwhpMmYw5VdFsNGkWzKL
Jq/yoVA8y1zBKYVOJt0kFVrhxWRHAV/CTYs0n0MHFHpikaIYxwjaAwdoWfSrxwPk
E6nFphu9++YTcxE4u36dKazO+vt737CEPRLtoWUrBxsm+1bqXwcTQ80AP8745+pI
sSq6diooKiQhfWDRF0V94JPZUPIrYFlkqPHoYmQ/M3nq2yBJTrTnw9P+AqKcS3E3
NS5oUsxPNW5zJy6Boyy/OkRYln2RfaQlsV2tdOTF/eRJRbEz90+NxAv/jA0d25wR
JV++qnf2D7eEYen9lrXRgPHe3yoE8wLZg+uwX33zU6bRcVxzGPSF0IJnU96YkSuo
qq7Ghvhvb36zfiiUXIY0WHvia+dVkzk0ZTpbsUyUHfSjXbsa9mJzRWIgUdlCk/fI
JBFt/ArWb3cX2UEZiqBzEdsMisS7XFSALGYRQc5Vznd0OveTVfrL107VWRnMTqW9
b2QeoMabL6N18NBUDHI2LtL0+G5OO4IHpKLIzl2hLWdmH2Y2dxQUye8q3CWEkh/v
xwzZODB97i/e64OjToeR19ag9ARA4TrR8sEwojk+J4Rh6lpvEmhIWlnU1H8bW2d2
BaePhkA00Q9SmxpTiH+hIoS3H25n24hWFNShazndDnPJnrkAi256IgmSB1Z8fhnY
MKKA1pEQcQZmNS37SHE9Nx74m3k0i14DrpuJH1hFlo8Sz04dVNfzP/9jyKHBjq20
HyknZKtknrcAOp6BfRbRzvaEFxY7ffmQEdPcnM/3IQO6dcjZhbf1thRVPL3qkyTx
28PPN/V3EJpRR5wldADYBaygNq/Y0TGVOc/cDOuIUCR1QLAaWjWrHsV5PaNeb6TL
CmJxyBgMnwjw/uBZ0FglZKUztqV+LCkkT5umW3Qg7zOVXEgb36C8IJkVZ1tXJAM0
Vw2MjdhGqJgzMBmi6mNX4yG8/unyERXT87MoCp+DWv4PZXvd6Tv8molO7FJU9hzi
/nAtlcVTnz5Nuu8zCX4UZo7dKYDRBhsPdqee5prVFeqpWqd+B23GdwItWTO1fTdK
d6vujh2C/Ztg/NUU958/i/ax8ypsJ4sJcP8V1OxdjJve71fQ/qm1HAtcIqrXw5KD
KlId6AaN9r9jvmmoFiEpQlNAq9gC8wn0pCOp7hfRsnGaHKPvDFGWJLp/ZMiJssK+
qfTGHCeZ6RtCGh13JYntP1zTHSSxzL5ONJmZ7poWj62nWb+P/QGX1I+2A+OQbdRO
Iq2UD84T9ewnCYLOOhGgAB4pZ9wYeyfPsa7nyqHGPW9mFmJP47HWroMtMUQHv5Vn
QvMwanQ5YoKAeKVieqGS1aeEFPb91bKSNW3ItqPdKuE5l3NqzMCfF1xBfP9HzA9N
F/pGs1hIp7/QK/AkNG2KxsRlD1wypZaughkVQb1jBeQcUjDTcU4EpkktSYRRIq4F
2XXIOrjAWazaKeokvlqaHyj2G53rxcodOLFdhpc3z85CFazohHWPqXTK72dTYor/
DTrxa04Li/GYLTHQ3uFto73g1ZlVrjztQ8+ns92ytkd2DVrBeTJs8AeX1A4zdEcl
6PlVrJIEpbQ9qkJFSUtnJHVwEvB8DwhkuWzpztxkqnIXTN4B/qIHDkwvmiNspTj1
EE+dw1gt2v21du7IPnvR52gBFXMkJJbJFtOQsAm2b4GEsZRIiQRm5ZRzblg7MkjO
tCwMrvKEZ7+2UuBo5FnT01itIc+o6cLnmscxHBPkYnTcIqagY3rBcPfaCQNYnL1R
rKK16LW+iUAtduq9X5ORpbmMwke1araQ2IGIOQ93+QgNyx94kfZaD1rn+7mvmGzj
lTNSSL+cC6xPx6eFnXANEzZn1K1JjwimdbcPsl1/xfgU86vAyTOwAQLZ2NpBYa+N
K7w015pxa9inFhGSL079ZIebQRPMetJZtFX7ZUP6h3e1yKeV3vnaHouQsKt/C5S0
hMJNZh+7y3z99V2k7vba+69JNeEmf5oHJGFMJ4c7Zw0NHpD38sokQOp3yhCJLywu
x1V+J4stW85oVdO+6kzVQkiOjSs9pH6oaeRNR3uPEiEfDO1PgyADoatveXeaBFk7
Wt7AmpluKz6RL6zwyk4aoB1tI6VWQEQStzSG6GDWEvKF0qWwoe39dGBzjSwu+1Fy
GAZeu4ZXHUUH5UD0Wjjh+A/kcVewmOQU72OoD2kNHPivJ/A0aabe3g1SDl3Rl6wA
/gW/LIsZ3SgGlsQiPhIE2SqEMyv2ClnuG2CMxaTSVWtlYlRCWbmehJit67LHZ1HZ
vIbR8wKTlFL3B4vKVf/gcWd0gRKCNRIB1H5kBLABmZ5Q6JZQSE4UXpOFd6v8BhAI
oP+bly6Jhi9/yFdQmTrkNwPf0FKCsD5wMyRTX46p5oF7FmtCKKO3efvfFc0Vmzbr
S5YZtrrGXNJIlhuAGpYxIR36JHNQyaMzcGCKHah6aXDSYuj/PKRY+M2VXv0OAi7W
l5l1RaIK+qGa6lixTfht6n91Z6NG0Uk92SKMJui/VC4A1GrQe58ZKKBEqm6hB+tx
+EYHPs9WwO0KFQPnEcmKaqBxw+yC40gxJub1TNEX6TthKsQ6XpWLI57cYrRttX3U
dwyBm90y+HLQIS72PAGDzhBYfs0XzlI9ghUd1VJSmZfEB98HcKwLAPmaRcxg+qLo
+ZsMHMzB3LlN9LQRsvi5sg1YnLg19J3eJ7cQa3OGSMx6HV8BJCF9pqAND/NGuhXr
JZBz9ZU8HD2hKgRc9WGiRzaT7zXIoOVdS/Vq3XclN6v7VR6x5hNTntaJmUmVkBvM
r0Jr420r+HQZqiiRDbWw72KgrurM10WBmBnIcTjbNLRdmRc4I4SudKR+wFYml5Ud
Ga1DqGeub7E5faT19i3St79DwdEjhxx+OZYp9iUQ1OTNDAFq9nP8L+XScek9QFuu
psSs/0oaAGY4qdpzeSonL3b3OAJBNytUNp7ei/B/4jz9uir4sCfs3FWkTVmTVfEX
44c+tpTfgUwy6VCUzMkeYR11VVbaqLs/xKXex0HgCq65HaUhEK29XMRDmFH5z4I6
irO8JbxOh9GawVghYvFsafomfwVkkGHGacPjNdk94fqLOcXEkOKaub0CYV74Rg6Q
Oct4CfTLk5aq78X2OKNzUxboZuR4hbAvCq8BW0qjXVmAaQZBYLvxznXTGWOpXIRq
X4pK+1zkqghgV5QWPFFSoRCAoiPOfwAp5I0I9hauX90m7CKZgna6zCzv2iU9V1j1
63BQZR9PqVEtWUtsPCfJXI35fKjhK55jtmSAu+EULoT55xLbjZKZMPM9D8rkAVpM
+soK9zVEhL9K635FFUPbUE6p7fj3L6y+kzlRXdrK1ys7/arZWXoZNabs6oDVIzAS
I4V7Ih1UNZCxWAxbbG6GtCJbIz9/rliR6VMoHC0CIm0o9wcjBm25C+uuURZaIoxQ
qh/nnR0gxuCKf5nAAZULDS0T26iLOvhkfaBxZPQ2Fyc8+lJXknM3430jtbLiUaAc
z5lRTPzmSH1cMfOh2yaoRsLvyTm31Sbq0XDIdCOYUplcSsu+efBTp0h5BC10Corc
Xa+ZmF8yuS+Lmbn93nKZGJMmNYbiaFp2CU83fn5Mr6pxGXV3TS/G0GoLPNkpe475
yBt/LP74KMKIptThyLCjneSDdhgh77voCM8v/drpv4Si3UhzGV4lh6Em8P6kTaTr
cto6tIMIbsFgEt+kZPb7jzPBluMaOlEL59SCMTxrObmBtSM/cwhau8JwzheYBHVu
4s4XgUIY+PmsZ2D3ZrKw5fa+HgbyEmhoW+OvSJnLqFsA0NJHnJXzSm9OjB7zNfms
uOX3YWJJkhWPIc4PQW1P/CAYIn3PCDabJfncyUGlM1QG0eRvrRynq82s7/T8VY+x
16nYPyg6hadnZd3ewFi94p2k01GbBHPQLfdl1x+d4y5lt5d9izYUotVGW3FTEcox
OmK1gidEvazdsl2tWoeK7mXxUyWQq394bWTqgA4f9tbSTrnfMkZSWry0P200VAIL
SadUhQ9U/v4+R/blqhzI1vKkXR1ShEqt1k6T8OuYh1rkGFKYSS9kMVAsDmPCpxwx
AbH21lsx4YPykrHRZYU9jErW8zQhR9sTbftE0rTiQaEJLPPkFTVptnrtdpkmZZdg
HGjGIDsL8Tzz6LOT6j+7t8Zh6pT1Q1s2wNJ4WigCpiVgRaqfUot0d/Zvd1UmZqKu
fK08D2GXerX/oIsf/oeTGtpJcGQ7A2vk3S9Jq+h52ttATH+iHUeJ9yImWQbwGfAU
T/iUnB15klcnXBDyKGRk9rxr3uu5QdyAXiICm1lkvHvRLTt/GlJ+A3w9JAfMZkc6
prkBGiUxCxvxHCaS1XmV3NAPyOxV9k6a+MLwRPlj7aslrXU3jGQQ911+v1xn+lMl
X5hBqDVs8ZqyRHv0y78eIi9XsWF/rVyOdKrm3s7G7oaq8Pa0RfFh5Zj5+bhJqVED
5qhzeZZ9yU3v8Q7exa25fTdGwvlYYYT9ST23oVsI47GlbvmPppdIifFUALyefxW1
5C4hHlYW5heT4QBPcWKVGQIUmPnU3clWHoH2QYoRsmE2zNNSMiFDv79ystUVk1Mv
Y/LQW870+S7TReAtCJyRunzvYza2NsJvgHdWbAlsmz/LNQ40t2eIjGdPpZmZxTAd
j4d6QQfng42naZtxBJ75Er5URiU6tOyNW2s/dRZQxdaOdTfRhjnhojP9qiDkXs18
x6Q2zx7D4lAVO0MuZEyM6gZpGEJ8h/wLN7BfbF0cgHn1vE4ttYTtEEnLenXmsSVp
4BSZM59oDN6huJVpxQhAdbh7GrYEgcddIE8EixvqMy1uo3r26swcj24mIqEZ1OTQ
HpxE+4Bof1yujQKxSnNI60FHnrty+AcJakfdk/IOhMUOhng7kiLL5KXO+bqR94r1
u5ZG0zxD4WPaQYoxRqCa+JviG5W+3umC/7ZWO7Z53RYLVw2q9tdin7e2icGbyb8X
gsuHXw5TJFVXX66VTeljAHmJkSrHiFUV857Xc6Rbv26ayXrX8/QBMrbAFm1LQAKK
om+446hjotSAM1fOCiqL+PSm8UkauY05QoGcxdfsbmiNLVEKUMD2Nw6Ti+h2WQYY
eDID/d5W6fSDyUUEVd+T8J7TdmKoCp0A8Wd1Uq8UPkRo9wv0zTYC63bvvmM8T6KC
GCbszmp9c9urZ0I5SCMzedUf1eHUeKMnGm+enHl3FYh9jnroGUcuF8Bedys56IMY
6u2aZO5wh1frVMT4MKrUngiJlZiVj73ATN9imySaJB/Peln5mtFOPYUWNqvscfZ7
NJ5Pl7BGib52VIJQB8UVZCOIK+VtLAEdZuIp8yqq2RGQ9dWRjR6dZuyZ6LpqQ+SP
1MahlK8K7UcaiRtjsTwv+53YZLMjzDzQ+vlz92haGgEyqKX7aAxvoTJrYoNe2qLU
tAfIvY0QwgQuw05Yq5fUnUz5tmI+v+IWQrXYVmAUNx8TRGI4DCJywwvYmwh0T7A5
ibX/r5o9J43q6rHrtpbEP/Jz2yB4x0BUit8qs+206CLwsm7OvDIqYQi4Y9kPteyg
S9WcFjR0dAR1TGJA6Gqug17mKmyGPr915p+yRjH8ng8tvfjGVjmETHfP8Pn2PqAq
HgQw+R+bTiGFwJrpXYfXR+sS4b0hVfUTFHMtCr9j/srDmT3yLNNMnyOXYzOXRZBb
7nHK2zhIIYWaqz2aVmSIpJxdObmBEGFynUAt1ZhRMfB5Q0nJpG9AwLS3AtkFSXFv
DeR0wqkdb2LvrJUktAvyvcoHiIdaseZPGprBXcVTTZRWYvMkN9KePi1Jo6hi7EzM
LT5su37GcXMZlqY4fK1vCZPdER+gBa90+B4In0g1crI=
`pragma protect end_protected
