// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EZNgtYGsQja8Y9bjxTMNqH93rcLzv3e5/PFlGMvmWsEqScswIZqKtquzii1nIt3T
/AzwUGwiM25PryO8/+ZJpF5HOYO3cKQXIh79dTbQ1uXROEvxTgkNygRCt0CWBGs+
5vsJbxtwhvh61H7dtIJP25UXIxX01Beu2KEnkjThYT0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6032)
A9DxZaclFpvUJUffD+QDYbGm/6/ATymc2FCdYWDdd/JFWNEPwZ5Z+/sSgwG/825W
ZBuVpdy0g6KFPEoADyInWSqZxQSHSMGgZECAZf2Eq+sa6M7r431WnZjiJDUG82LL
fa2BMzP11VSSfFxk3fEVmJaOtCg348iOvqANpsUpnQeU4m5xhMZ41Zf3Cpk5z1pe
1HbJFe8RvYBtwzf1yr4xf8RXySTL4YAZWkbYiGn1P0j8oHBnpgz6Je+0iQIV/0jY
WU69s+mHHur/WkZRL7Iki5vLVvXxrAmb+jrSih71pLH7xsnMjjXwEht9xjCaAx4G
GSLt4aG/7BRFv7dkeumQyf12B/o0sdfLP4ytL7gRmIZqhwbsBpZaxkDjF+SWuAy1
VbU2bzfvZxYVpxKk3Dbb8m0wBrFEQFQlFEx+Grp6Hnqrdpmrpc8UqhuAOEuWCyQR
Tmgb2qxyuAHqAlKDC0VytyAMtgIcSDLyktHFebJXhimSmbuSbWdEpsAwPmhX/XmJ
uVr50+Jz7sEnIcailYUzpcQutGIUSNGd+eTkACeZWDoohHiGj1AA3oTgCAe7LMVI
Nqp+dAV8L/FKUmM6Am/JNr8OOoSWUpTGpirMSnQpYWYseZt/M9oElMMHVAEhRjEs
Bf31IXtrpB05PvqT6G4hCOFnNclHvqJE10ktN6iUhZVOrF6P63WV9AIn4kNIxq16
4lFrSgcNkii1c7koJa5h1+P2JxxNCHEfapbHpOQjHBNFCrFOh3M+kOf96nwEoXgz
E7+Qg7wvVqdY8Sxr7xBY3qwNWlWHYyCOGoZEWmru1DSxSr/KNjG5KoZd9tnASlNp
LNf80P31wvIEN0rZdbq+yTj+eujru8ppIT3k3Q4k/RTRnYzEkh6oUT32cNKeQnw3
RNzJP0/XyT5O9K1xuQVs7HAEFrSx40ohlr7xuxx6eB4Q2NVt0CLJLkjevl1Ff639
xFPUlO6a/0211NkfpuPXsUfoSQK6Dg+HI37muIwvssZNSpC3fSN5NKfCd9dH8E5D
ZcqYdx1phrUGhgXnNt8MhVhVvz33kiBayN5+1z7aiLdsYJgBFFscEe1trzACnhy4
bp4aHLBs9/fWZmPiM8tNO2hcUJnr1X9rt5i3OYnPlcU1TQeawbNXJIzFnqHjAcZg
oF8uSLJJdQAbHu1Pv8t7EVxwTvpU1QToTRDNMkyWqj3TtZR+BYYvldw6oyrQ243h
cm6SSR+4zsHs5VsXmUe6t+1eIRrt529lrlfVGVoZaXnxLYFWsWBb6CWbuzGxMCb6
jy6M6Uj1oWjaBw1bSTAHQQyOzQzOixAZ0FrCRvR6qq2DW0TWLW84XR4ar9r3KLv6
IeRdIxYLIVhD8owurH2gV2jURGfrUg6sMczzVibH39m1Z/TggD6y/ygdMydI2NkO
jbsoUexgzjSnP7XCGu3VKQTQCxU8qEfnuWE3qVWlTD14nA8babHvhht1Z3vHDokF
RKp1NtDQaxh+WEoDnniFHadRFFi7sgGCOjXkE0OCQ+eL0p39f9XQmXcOO7G4DLyt
hRP5Q3EVEUFyxewzF4+fKi26DXfUYMeOAyR4NGXpA47RN7mQTrr60uiIfJYUtNqY
yVqqPmVazDsjSF1DwsJmMg2Ts77hsvou0OBMn3LZdxF+hUPMmCRKXoMaIL5V5oTc
zbbHv1vPqHy/jhkfTdmtsA7kO86UQbD5ucwMpP95twBp0UrlxCbIEg4tbXMfxzHn
hlHnfNUQy0R1BPP2fP2SkxtsmBZrPTlLpQbuZdDG4kk5+8xzP6Ve9HJyd8ArIDRG
D8nM80OX/VzZaFydtx/QKLXgR86nGCXMlDKqcIIgk1l96ajP3kS0wOylBD0LiQl9
E0Gta5RoOjncQjzo2UP2rWaGXKGJaNj0SfAtZqn1an0tdBx+RZjL4z3Y4SUlJegk
dGU4pM7/bcNCXu4gLkrkxr+jclHsNIrfbsmO49sr02lID3iNTetUWDPTH2JehaNn
dnsEBVP4QlxfL+ifceUVbzT9Tir2pVYvu/9pskcPEVaJU4NnglzmbTrA/MXhfFKl
z8GleMrfUSSUrPqs5jv62zZfwRxOQ34Qojtkmia8oIBYZKRaDHwV/+fFYPL/T4nr
8Y+VJ0hO5DEb91UMvBWw52Ko92MJBKhp7yA88gtTbuaGaC54ViuClcZIrJKr96Ed
WCoP9oE0wmc4WTbmy21tRYqzDoaUvsk8cnWshYO/GpODoOmk+jtIpISa3d+YkADb
YN3HU1xeirb09B+OKP/uv9lp6FCfGiAsChv/KQAiLSpuTW4w7aApiXwJ48khmEEt
BCI7JdGgL01Gf6iLI4NMNkn0viMeQMfwMOZgf2fJt9BmlF0P7hUQ3A3H34O0FUBa
GHxURVJp75SArL6TMCv219Mfp71/1gRa7KDK0OJs5OsYKULQWWWakE51WF6CmvQc
gAOvCUkdQEtkJIVETIqaqm/c/2YBsbOIk3heBnLGs09au9GW4Sg8ZJ5j2XlX/amK
9m2h/r2vfWpV1+XD1wGmRANSw79fgyik5UPHCrq+lKcey9qPiStqDZ6eKCPUdCqN
6dXREh207krB3UufrDAOMNr8hERTydrQ1oM2BWU2RsNIiqYl5mvfbi2OwqQwfALr
cASn3gLjO+INrgT7vfc2JFMVtuZBHRE4nVLpkpSilqgekiJSUBmHWZjAXpe2OtIr
SdxzJv9A+O36GMFAU63JUD0xCOxJGS+Co7U3g1vL/YSRigu9CmeDW/8LlaVhG+V2
lxXwnBvy3J3nVSr2bSEoVgCqeHaBy7aMPZirK9Xr1oBvjk7SHJcFXhTlV/BojcAE
Or9B5xCOMWZvx0WdRs4Ckph8deCfTwoDTHUGgp9q1i+Zj1Qcnp0VLi3iWjmu9gay
muPL4ideUNZozE8qRSHNDreRKEOJAEAYLUsG65goOVsRtS6Vyi6jp3KVtvkYFJlR
/Hm1Ws89fz31VuWcLinz6pSXLEpksSHnPa8IkuXVdJ1hrL7OUoBspi+LT5ncFYSc
jOYyQyRFvn+VsvVcgy0nOWwmKrtc/Lbi0VFA9RP3zT2EMMIYjbwf4/dgQshiRKVG
6hKmwcgxX8Cy5fvjE3UYrGwxKklDf/zckMn8dbosGz+4w5Pdl4SyWZs/rsuUtJ3M
ErHDyPsVAsmZ37uKKXD9FT26AXtRLEi0xNWNWwlkBiHUGbYChqEHQ4pqjvZgd3iz
5syUVX2whJH22KF4pYCKEHm/pmM8Zu3SMHb1iMay1KU1vptYlcan/eiFuHlGfWcC
hoWLwkL1Ta/MyEhK6faYJQuf85QpczBOIP9wsOX5XQCXRJQ4RC2TDr36W2kFWVKV
pjgFUwoG9sIQy4kwZizLsKvkK+50nwZuFcNFey3Pdm0QwKbTiFSRVXYUy7Mt48j6
NOFmIejPFrKBQ7xKMNChsUX5Ti3NhppvCGrxkd5ar36/gsbb0Yky09rpvDG/nHji
De1t4NdoFwXTktKGT9j8EvEERjDMk5qkc5YIDGxfJ8Gu0r0MjGuS+Oe1n///dK0p
KpuCuRJxAmKO4KzWi0eFcZlW4o/fbwhx28SsSt7/rOm5QlxZFkVFlfuyKd/8MBGr
NKly+BLo//MSe+fB/uJIYbcV666nYDsMmld+wIw4z+vssTVpMjMJjcRBo9WvBAY8
4dCPlwDZXAdsJZJ79wRIXLe2v9w9LDY6hF/hu7oozMdO0/IFFz38xtQW5lfLeviJ
Ko7toPSxtV7++1W+97jt1hHt/dmKw0ixRT5932jpF4N7+RyE0yr+En/RS9l/WV4N
IwK8alwHrm8V8pGcuuCO77BWqnqNVWWQyQtaCJNOlnwisdkq41itw/Opx99glPJp
n98jzXtx6DlcLXMwlLVRDPCxOiz95Uf7ftwDMWDBpVigqHwgmARbHEWo7wz7MEZJ
C9o8kojjmfrhHHLza3i7UqfTJu80EK2DCq4xQc/10F84+0qDzRAumi9wOs2DbR46
CIRq5sx9CdD+D2hl5zwviZW11+UafDFwYGJUC2HdloAvqlv4+X6nQsVF/iEuA+19
JX/3J/IKfjSq8JmgxeQXgoqGAVXiAU27bfNQmqAMQZSfddXyK/cYnl0PjD8Xin8f
A+9MTeUWEK7T0lfuBou5qo0hRjRn0cudobVx6J2r71snNcUsuU+QGEVTTmt5Ln7J
ClloeqqqZOZM5Zdkx0mKX6T2L8kHzHg2T9X1z7ATdUp4fUEH/Ji61P+I30diSyMJ
zuh5+l/j9Zdgt9ML+7hOy5zPkQmWUOmMHUwvu/mA2Cj5BSKJRMHm7Itxqt6KHJ9O
m6rF/w42wK4BYhd8BbKcXzofaHpTvWe0KyxJBjsmMrennsFiu6Ar9A/xrYztq9Gc
CH+OfHjEYYC4dQPWAetK1U+Jt1C5wjDGEWSMgCKtYAVmFmx7Er2YjhzDAvw0ohzd
Hiut2xLun/q2hY+eeHh5L0Vqyf6RKkv378xlTHV+Es+QeaeBIsJNumERJ8FNCm7r
fgHPuaeF9DOkzpQAmpmq78GYyfzbe6pX73q1YMxR5ceCGzbr71afgZrZP00FH9qx
wz0+rh6Y9sIoTnEIXNbQtwlsk4vQ7CEX5SadZ2Nh1cuRltWemUKwMDtFNk+jbOUz
vvEO0w2bKubSoOmXkMLeHEil8CntEiCfx4ykOQ6Qze7FNu5LAKONbaj7o5FRE5sy
u53MC5MvYqY+q+LMfNgjKFyRy6iDdEb0tl+OJzXZzqmjEZ8siwNqtEFEt+DYTfAS
gvJ0e2HQU3wT6oyC0l7of+Pru40kuWikwNlufPN2UmN4aBYQ7RPvHZnLTD8rzZQF
DqzwJQ8gHYDSkEkHBDkaTRgu5gCR5V+8ajKoaz8NZq8EwBeC27RNO2/vwlWtTqRM
wnBdss/97FXwewttO8E7wL3oBR+6WkJCSLr/ll1iJdI7vlKIwfKxLidtXkY3auFT
f7QDJScxSHA9Jh9i2J60ncV/stvqJTRR70lGj42o6UbmbVl9zyNAHl5RL3S0SCYO
fvBoLgMjTlB6+Q2JkTvq0KX3hiUMwujzBkzQdhjgpUgZvFME3eSuJVC4w8gAb+ri
+zAyQfUNp0bkm/apgJw+VtcyZ4OQ5dNTGjM2uF6Z/PgwPDZ5lo/tL4e+H+ee9XCy
XwmXBBMhiPI+DEwWjT70emp4XMFw8yJLgJXFr0mi3wVTQKqhUa+d7bz3jScnIHmD
hvcDbjWQIfpmKdHEVSOUXuhYLE+r3GhTIT+dbr4e6djTBK2hZ2qepuWgR2D9nwps
xz3OUlsJDMkuNEM8jNkR5k6JTePW9uo8vfQUHNYthPhO4TxH08ElJS8fwStW3i4y
FI5oqdWwJHFGL68zYoVkpQ+sHpZmUVE/MemZMxnjGYr/1i4+Iepe3IapTRz6lz2I
ryAH5JQtjrKDSjIZWo0MraVJyxx/hifdA3SOmSg27MsMn3X66f81JeXa1k0sXFRb
vdxCtI3ZMrnG7zQXa2Tj6Qr6iJAxJus2P4SVL4FZl1zxGlsKbXr5cAwy5aByi6zg
vFMlTyV+aupdfxAgeEQ6eOVIsnlKKYlThSR2/dcsWrtsgo9ML+Bz3hRQhuSeACOA
GjYsqNyih8aARaDGrHSe9GJsG5qWlQRjjAx55QFiaG7hxzBbTtC/WPEeJ12XglHq
fnGNw1YElMX+NH/yEoUNQZNZKir+ny7t55fgK13Y6ICQ+6vGNcmlwmVmmZ5fxGFh
V+SaWjAfShqhsvNm/aBKJ0aF2xqNjpXD0yV20+jb7iKDAhFyvaTc/8TpO9FO32pk
d7JKBp+d5swA+EkbMdVrObArsndhhglOVrcNfb9JzRjuItDkGkBp8JWJsF3caYAo
z5lgFsIAGS4ff0/m/xiszHREF6PQX7UOm9RJex3SaxTICt+yp8qucP7P5dBVJASk
fye61M3DRfLTQBjGjlIcKOdz0PISNKYQ+/5+DIqm04wynCoZbykSHI43k1q1Iwa8
JiOrj+R64Rd+zggjIr8/iXUJgjrsnjWSFBl92JWuwTUrt0QHdIDJvI49EPbB7HMx
dD92Lq/1lBa/G2JAjJz1ltjgPzPtB6G6Wbo0LAAnwGhfklyZq0yELhyzt+Cv5zq7
ptOxqGhwO2dULi4qESbWyHMDYKYR6L5LHpoAvJQWj1isTV0kLJuG/uY/JgcCiJpe
nxkxrbqCGDG98d7p6plBqd/MWk+kKCs6l5V29EdMTt+BT5f4MKypAuClSgowzJVX
YYftOZn/vpBK5Q3BC0x2Lxr72ICdiVBGgB1H+r0NooG3g/s6GbvKA5uRdjUNGJ28
7Dz25uniDPreXL4HaGmFGwC5+yQYtdVrw7v2smgWkgUPJuWKxZKCYHs4N33jGinu
2ERPzGBowD2eF5fya/7i44XQGgYz//3NfcVsYsaOanS3I7rViQURYpuIH4gpJZX9
wnGcURgx+xFvIDM+o6LMqjuJ1g7EiLfNOmecb5sAWAov7QYEnRLsdtdjkIg66lBI
3240jlfaahmaxpHZa0OLPPWuAH+LZ37dYHVVyY0MYAY25qywlYjb4v5kfIl1jXbO
X0s1BITaat5YKj70nAV+Pgm0x033L1gnDq9yMfrgPU0o016+UcLFVfMIR1JBrLmX
8oYXTwZhhHLDaldkAg7xJskfCYMYNiNxz7x0CpJ49qXfSAsQw91XxRanKgRg26G8
qmRjZDhh+UlMEjQ4KP4PS3lLwZmH0K0HjudGPNRRiY7bxSnGkoWyUPoZVgClT+39
SkBxdDe6sXENzbO1fWfTQGDX36LR/7mTQFnaFuCoEVcIGGXJ82A/92iMCcwep2oK
UY1IOz1BRm9fESb+nmZ3ygwtX/64KUWagdDMtF/UQFUwmp4fOW4guIESpJ/CdE/k
Xzwm+fKg5rC1uetBOEMmCMS5kJqa9vX4MxRVsvLTF2mSw87Lk6OB73uD8kVeRB+Z
XcCSq2ht86079RBIGfz+uymXDh/ZIuQuwiD45BGx/ZicBuBS6zaRCYuTi2EAJ9kv
srZST/OBdX2kfk3MC9F+zKT29X0kXJOJeVTAr2ETTtiV3CBmjmW6roP+n2cCJdp4
zAFTRsCeGMS+8S0JCHe1sYWfoC1LrHMtEtdyiGVOJ6o3YiqiWJRcvElyiFw8rmW6
NfsucFEtd3SgDROsSqmTtc06wXfcZ3KKWCqIlgDD/c/xvYW7JeW7jEanHKq0hhks
9OBgRoGyYOig8tHB/G5aoQqNjrMZULJ74S6nKBKcVC8NqKi7QNLDNq+sCHHACi2d
pPTRgVJ804d2+jf4ZurHVzIZizwBXrOdOrFUaFX6VG4fY9cZI3Sqm9fHaUbCva46
J2j9t46+P5B5hjaNpHMeDe0zlUQ3ivIktwDRqigvuZRaGyC48bSufu1UgM5eK3wq
mw4gYZlbTgJM5sSBRSBkgfRTlKxNnjneHuf3HGtD2Yr6RVRxr3kCk3QFwzvi4lha
A5KUqmK4d4Q99XxOqF2axCNccpMzIbZCSFs7JJwbWqR1mowfKQqQTfXQO97owEZF
wVg9+Bao/5/0MsD3GPpHffpceRI2bD+Arf3Q/vF8yc229FVtBkf/6MobJsciyAB4
M2qS0B7F/y/Lp5aOmQBhzsYVP7GEY4aZwDyGyZEUA1sH57hzVnwIRG9AI7T3hSJE
7ismA1qYlXc9P5+FYAFl+Ykg2Q4I4rkHB2tP7jJV7n6eXCyun3ACgUX1XwXQn9oo
u0YLV4Ttp0itYCH7QsMebNGl80yhPQ24NG2VCqkA53i2NoiAxEY4+L1VcMMZALuu
PyFLJA7fknnCkasaF7ZPEbZOzJNwTZUSh5Wj/M/zRs2HtRcdATyqJIkWarqOHj4u
TGtl1QXPBPyRQwO2o34DoR3bDDZUBH7mzYkmjwafttJJEugL8mVWnLjmk1jNcipy
OuX567vmpakR+f/8GAEHn8vOf1OWDGx2LPGxyXKsKKL2wcqFTDa3uVMXx6u0YH0n
I6q1RWcy/EqfGljNtIAGFiB1ARKhQT1UY37hjLdrNaSm5VeNJuqf9nN0+7dl/mJY
j6cnk+8SIfncExvx7qzVm4L0t0QuWCRV4DZh0J7SPlc=
`pragma protect end_protected
