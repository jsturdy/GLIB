// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cYeWKobmPjiZ7GUAJXCGi4vc4OG4I2TZjg1ORDcNnTztY2oOKz43AL9TWBA6jlLn
yM4TdgR4jz3HcvHxW2FSGOyt6zw/Pcx83Z8EQi1dnsS5naxRktLUshvWFuxmt/4K
Pa8Y/V7rxXkgETP6Il3ITH8VjomoG/+29Ib3Cs6fKPo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7472)
ICY/x79ZwyJXhXWWYHrX2LkzJRNLJfwvegGfOUSU7quOdfdQkl1FNwprJAmh67p5
JWzNyZTaOWl+26AonVEf9BN4lTfeL/K37PE6KQPcX0uqvsLZweVAF0mrKWMWOwMt
c0upYvmRYaFHO5A6wtwWhLW9e+vw0s2z9C+WJiQH/RcyepByr3bkdr01WBzLXuvM
aGpT3RBnWRIr/k4qeLKzCreuEAs1OBpcbbR7Dq0Itn62qCCX2GzUiIgQr6jb2xEt
OrYZGKxiUodQ/3m4OnVNbFE8NyigHDwyAMzpPWF+lPfm2XQaqk9aoD0fnnTm03BH
d/yV2s3BIK6rAe0eRQJxiqP+k3Lizn3b37NAXgYRG7KxyN3zfTXtH0bmwQUmCvZf
duvdwkLZh4y19PKNGod8d160aF+FJ22JcAEhdRa3LGvIxV/Kzvj3cBGRI4Hkqh5y
KnuqDMC7qIROeS2o8WahWWvI5o+Dl2ui+ZL/KMUyGOB+vcfafa7d1VZkDuAb1qAM
90zrsGkQEx22NSnxsLazM5C7lAwSnVJpoBg1KArQNKvj32d/TpzMGEvA0ZcVSWGU
ZiVcNxLngwdNBJqO1Bync/WjkB1qI7erZOnlOlDXQN1tq1Ai5HciEx5fB7bLKoSO
Y/6X6XFc0dftols9N64rNM0HUvGNKg9ze9vrET4XUQXdOi/17IOPORFcB04x9zgQ
cdeAKyg0vhzCno/ECsEf7dqesrWSXbftsROzffFs61zn3RVOVyHH2uihn7NDszEi
H8ZNdOp37UHt3qu8LR+2bKPiIzKHxhezt4f0TKIvmSQh7iyWp7ER2UyNHfJnuqYb
wfU5rMx7zYwmOY5VrDV++s+SEkQjxXAQHEwwV0Bl4xkR2aXzOgQLjw96dmh+4G2S
vCO9KD3MMfqm7whfs8srVggyJlKiQvQCBB3OOPImDDGTxBVr0Mr4oeiMNn4EuYcK
MYRfGfxLpDUGVfn3tQQVvtysBAKb+4Bs6BpKH8Ymw7Ny8lKCvELalOvU0lSsjLG4
48Z22oP3rWDaxDG2ekjJt0abLNGJ82hNg8VvJmgqzSyTUC3ztVunB+fWhkTvj4kw
zuxetbeCOdzoE9OOqLWNcxH0nuUO+sYCazmCdi5PM0AH01/jo/5WtPURRL4RFjLS
BwDrMkxdV8ckjJygHni1QjXgnf9IGKSBysgDn21kNGO3ur8zJMSqJ9wLQd+BLsSr
to75lUIC+kpwNylrLuUW9q3hneRf2pJn3OWHzUNHiCsSmhX9Lawc76Dm0PFTxfrp
cvNumJk51Y/3d8gmhMsqzN/r9b5r9+Y8Qw48w/tTHsJTKTmDYXiq40srVlx7pf4B
A1plQe1sV8kC4kOEMeyzlFB6oUYsTdAW5UaspUEYfOfOIGP1I6U9OVIcbcs87EpN
cZVe91TgIC1uQW8CJpYpNQWp9LzzkK6dVkf/8hyjXzsXIaUl4ULqdbSoZh+dTrDX
brT3njyoDFXDOWzw88EioBjtQf6CkYsNeS571FHR6T99sKodrVVP9enkru4BTdUK
3wvSRWIp669smH8jRbZ80Y1B45k2PMN5snLsME0O4kvCyKbk8VU9e0X6K6Mvjn29
TyERPEMwGe62Ua9y3bTDW65F1eUjgdLK0vTICoR3sY5jytl23oWZbv93aUTvgozJ
5kGmDvo8XykNirySW6K++E+usbbcJv7Xtw0oBmU2A4F6Uls3WzRGiC8MkPimdVmk
/wD27VF8UORjTJ/A83bx9qTD8NFq0g6ZueHQ3IJ5SzXSUmW8c7AU1z1IqXGnwqEU
l3qc942yCpLGyAf+VH6EvEBgnWTC+UqOI9clUekKPRg8j6J2FWSY9YLcXHB65n4y
/qYritoeMt+Af/SBfhJn9AbVQw8jBqqoKKdrOiLdbYWE9GJOCzQpc1yPO2o1i/6b
fLjTWEP3HegA8NLUIbFFi7xJCtWhZ5WAU5lUPFsv+r+PBBo1HDHuoVRhBwHUCROp
azsDDeN60VupfdO2Hc52kfnix4R4zJv3JLsS1RGjzItvhfcmie5sN2fzO5oZ8Hp6
w+b+9OpdXRHc3Vqo/X+T7HgjutAKyjYLlGdtH6RdYANcjEEQXDJheToveZiyW3Fm
wKpxUyOWsGiIkG1WIuV+7wQxkqnsfpJo0pYqBW6lNlQF/FCa1jvpouqyQkdjvoWp
+oL9APUaHK1UelBgQKyExEa/uIIXmyG0X//IArLcfzkjtraQc0AXlz6KRpQdIhNV
8cGMvBSjadRi8zNECnbi5AxJzGSiixC/13MBUuGgQARNLO8iQTtODgY+wsv4Z38/
nQAe9lJMDwk3s5bC1lu8LBrAa1AlTzt3SKcu4Cbefb5GcHSgrIdAH+W7+xF+uspo
fA8xOk4kVPNSBwnmC2pHvvO8AwAPthTo+nKY4pgixTgfx4AN/erL6kUrU4dpB3Cf
pgDkP1wtZrePoLF7e0S5OA6NIT7UyOgGkNls5jh5jccQrkwdgLWWRB4tRkaWNGcE
KDr/Tot5LT42LYYgVx+HCYQbPUKMA+ywLD8+obkjqx0MP8gzesg8CpZgoFEp9/FS
NfdMeW0VZzOw66ZwaiqenPze3QD+UaPYV59zdBpwJKxGcvT/Na1+UGRRq61yAHXu
QYjaK1EIg9m9lS1zRfgepiX9xrlEnuWEu2xajexRclDlpmvfwelAIXuvdF4OQMWp
qtj47YSBYWta5OZZnw9T2eYg/zIC6DvDWZCg1JdUpmBH/xkrcF7Ok2xqFcv2c1AE
cRDMO9ttCP5QUdVnsKcEo9ocE1stGqxEEcu3L09/dU0KH7D6+cR8FAjzQFhI+dEX
C1+jNAfanlV5XcGPB+AOP5oJeZTD2CK4+4zeDwp5mWXcigquWT6sD/c+aOhEceqo
ZASchcbl35Ir11k1JV7KgrTclwDXE/EtudI8tPnHbqBR9ZDqO2ZxrUgPz3VdTnmj
UX0bP57VNVxr5JKmuygW5u5GcNGYzV5N7v7xPfzB9dgj13DQjknnvLOeWon1Z491
/Vy125aMCMs1uLdOlte2bYBaZxJmcBV6c9wf5kZ1+HxFsm1Z3H4acAy75jKFnLEJ
w/CnI9WmxOthcbL3BxLx5BOTfRXQz8wwUhD3fomNr2T4uftELJnzZE3NPUTFao45
quhVxQ0Dsf0VR6pUkoNEau0yXmrcRjhz8t2iSSEx77NLNoGgwuOkphd7eBhwQ+vt
uFA0pFCrrMpv3mV0qC6B1TrFC9RX4tViY6pMTbWCW3WbTes0qLCS6YGQBEtKt+xN
33rDsl1f/XAz9+dy7W9WUibTEVoZS7CL3ioWWQkLTbSCvlbWtIOCK7f4mwIHuitr
VnCYPJ9MCSi6YulGazBTH/kp3MD451FgOD4p62RIYZQSr3qg3uFo9+QDFBxxyber
XMBd63Q9lDgqkmZ4v9RD+j1XAh9HAQ75CdhwdPx4Qv1KMWIK9ew9AE544qOb1i3x
rIORroKLuAxzSpI6Poi8FYVCUgkF3MhD1UghHVXi+FX19mbZo4pNWZhr4xEfuw0Z
kMU7wlcYL0xdM/BjxuGGCZ07zd9WYYpryKiFoKffgTTp6ycW6YBmoTkjV9bbmVy7
/YXmKM8oBIai0Ww4ybrnzctojSTNnYbe3nGulOjlvy9IGrKOGBGnNVdY9yhe4Jzz
QDLU182Hlh7tlkziEBPNHsLVUydItJb4fuH1GlNCtEuBw1d00MH2eEHoAhdA4sd9
c0/lv+GMsE03v1ROlQccjMbse0/LnxCMfpZbRCM3N+8qK6TadfYiUHv/wdcWEBhJ
Mxpg+zPT2tXC1VGmuiW4tSCGgEI2g1lqa+Rbmxw5+pwJnHR3jjXHpuneSg23Malq
pZRqpbRgr1j2xKVrvBUC8iqwRg0l05QN7kTt2Hlo1ioYnQG1LuGDBMjvLjrA7UAn
6Cnh+Vd4ue/IMbw0uUy0GvF3Xf0FKlkuGiek7EYeUvH5SNfDC9ZHkwaTQs+TL2Or
6p81BqZ2oUAzkxAzBWQp9IPOf5hwvNRlgDHYNPVvhQ9+57UnFapwDRdKp6+JDHMS
fwY15HiKZ9zpo93zsX7lM/AAxg1qUfOfVDSwY/TcSfXuTAKul5n8NvIJMiyKBxj5
9+q6z772Ttq/Fsvay1dWY+pkTsbUkCpwJLqD/Bhmo484nxUaJ4E5xNrgN/msBg9J
hBXyxWXD419p/VLnxtnKp5+grUPsHw3Mkt8cm+JnRAJefuK8SSm/cAcOKPEltn5h
JokcngOuJZPnYBAS3lS04RIcwr7OgKDpdrhGFD85vOmVOHs0iibx56pEX74cTbCE
Agih3EX0IIEhmkHxlI4UzGl0QqpQiI/HS9ncB/6LLUEes1x33qLk8glM1rZcCc1Z
VlsZYtE+5GuccT2MI4yNPWmh2Q+EuxSotxiZyItNYVeFJ0DacQNQb++ICyjsw9T2
LsiHcuVK3PnPz9Cmrg6cnE1nFs2vzZ3VZ9XB8gp4Y0fIjXjGJQXpfqkugoqe9O2S
lTYYEyD4bfkwsSIg0ddqxwNRyYiFEsZMRWUWEB7X8+QQ4gQwkwddxBuI+h4FxVdF
HYR3LCzUlJnTMHDUfkA4fm9HDtTYg6p2/1khCEwz8O94d7M5p+onpLgf2/b/tAVm
Wvqf17h/AMHVamaY6OLUYL+nwhxv2sXCR1r9Wk8yeuf8Png2W43pzDf+We97G1/A
IbUZ0CW658i718ZxjELXbi6rY3EJ0/xenYE83luF4vorvJftf2EbxRfjupyBgjgH
Fw/D34Tu12mMWet8gQX72Id3whbHwOm7l8AdMVJ0D+S9VMfAoHEC9EUvQhDEEeQE
r5xUHgC8DEmp3eN2uN4hUu+ixKMkE9p6wy6WVhb7gqhfArHShxZqTn89m4BuNFGH
xvXETiNmQZhIFLZ1UUWAOhXi7ncoaJsOyVKM08IyvqRmK3M19hXvbPYleXWGun2u
9RgER8F7EYnpqeupIb83Uj6OY8KJ1DXvOrsokPWc72AU3OL9EEu+//U+JCWAqd1x
WqN1ZTJLE/q6rFfMuz3WydDEPEnGod184636mGz+Mub86EPH30xHtnUqLpR7AzoL
zmnuN7hXaJvSL+ahsmA/Ef+eR8IUBcn0oZ86onb/c2iF6jQlRl0Wz9vuFAmpHpki
BFzw1mRX+l2gT/7Qg1J9iumDavo4zTcfyI/pNiie1ATQNc+dcucg5n26n/edcATB
ouHxC3mK6sqNgrXme2vciZDWKPZCia9VujbJADxk9fi0uUt0UdM92eZRfb2LwmsN
53hAH3vRz7CjGKDh4B14svUJWJOO8laUfB6kd0AyhML5tUgBNMM8Da/pHAvih5yU
o5RcFDcVOCBtZVcXRQ2Ve5nTcR+LbS8iQzJiNWF+YleznYxN+IXnOy6/PTipQSem
gKtWdnqxr5s68KCR2f299EwUTRXsg+++d+oHV1FjYZ1haKIXJsRykluUm2eFXlUH
XCXUNwxHN9aKmWYkUCstLVA8KfZOrqs7UE8KjTeuYDeLqo0UuxCBd4zO9WUXo6Nb
+IZvkx92R3hxvp1ju4LG/FCVpWlosqBNeTP+HAKI0LtT9i75ruwqD1+/fWXzX+DH
LkzXK1kuadnkgYzDjt57DD0v+ISFo31hF1dIuKFAJqLjv8IMkHa22A9Fycsi8QNi
Kgc4/Nwg1+RkSsME+TJQfm6r8T0NVLOc3aO4YNfo+b5ZAFkK68wQX7zMd20QhVIv
VRSDrZBCsZxBqlEBgk0Z0gWYjzUea/NDe3zXjkTRsvT+ZdOkQXul0ehMi0PtNcom
cLY/O0SKiatMzOD1qJ6zOgvbZtB4ShK//vazt4Wvh744EWhoX9GZwXDGgNrhkb7Y
ZgHmcHbcORTs+JKaeeFWSw6ftUJuR9FhNgqEmPzfcDzQMxbDy83UiJ4cMhTUTtIj
Yi3vdW4W+senR0TV3XxweTBH871wlmSbHYlwlYX6JB5njb1j2ErMhMq9IOvHTRs6
h5G73fAyPa3aaWbuMyV79uEqlzuEro2EW3PMBNeX9Dy8Gne4cZH/CMt/7OysmHlZ
eHWgFEIPS+Tt7wqSZOt3ToFYn/f7qvujkzxsfX5D3va3ky6WsZ5kw9Ih6xcs6Tqs
qJtNTmD3ZjovK9ufHHZSAadC0IObb1EyG25/tJffmbBemEp+DqFwTdcEMbnSVvmV
Z9Z9DSnkhuw1mKbuxL2scwCMPbMOmvH5sPnTkcKj1vq7Wk580DEvZ8ucc1MfMclI
yJHOBmp3S1BDJxLHUQoSfL9w6Z2f9TA9sXVi5TU1ahYgbqEbvPc2ONkq/nT6B64l
Hi9WiiLlbzhcFKn4m4hjHsUHnr3sNMrmCvz3+VHZzW6ONZQLjBA70fNj3wUV9Aob
6A5k43dPGYedGJ/h9WwoM1mXTPs/WeAJloLyaIKI1gUwvd6FAxNeipfaUGAsSxc2
2pjI5ZlGa4OH2ML77qUHXXufK8J+93ZWR9aNulYov0WilYLGVawSWahtouId3V3g
XSt+UIpDdAmaGpcPqZZ/psyd7oZbY/A5hrfxF9fZfImJHKSH2Z25TAHSwsJNAC8l
nKQU9It7bPO4KuP1KH6qTpsCxV+9I5JmtBEYz7DNmAes5hpa55BJCx7ukVPHsMwu
iyneumsy8xKs9CymWDy9kYgXx+2xSaRyc7NWmplSQSuwLdhXAr2rfTKcVkEDP6C6
0rocxdqVM48pqbDTrkJFGc2FuRK16oTVaNvoqK/yUIrRIsXAKtiYNoigdgPdPbsh
gF5jDWsdFg+qmZ3iRbCN83mFG746dRuth3SZvZC4W8HWZbpT4OJqdUdGfjxZkO5c
a1EDtn3y7NT4ZJAEdHcJzXd2I9/CbJxDiISUQ6mWS0W6fktvB0hSgpNPhOfgyX0b
HYPx8ltmmmGYrXM+uyg48D+4+Hzsu3zTSYtC+aRfE9rFG1LxhntunYNPx0LAua+U
UfW5W6fJH86eQanlKZ0VtJXInMdox8MujeoKXqxEToRfQCtFw1hSS0ijJ8AnwQGa
E/bEenRts8IPxoxcRsXzQJXaobWtBbntJibcIvQWAkeRUhGSUrlkAlJxKbJHkX80
yAjMa2cJwFTmnK4UPPkUC20WDBtET5lFPDJrCddRxbS7hTHJ3hhZ7c+uZ6j6dXj5
eaptMGeo0wRYu0UBwGSsFjc92mETJyxnPsk9ihf46l5HHcTvWRWSiZ1PTgC4cIJB
+YrpF8APQwZvUNUNda73Wun3O8M23gCmCaTY2FgsN16RfP9MW4aqR4S7TYqxqrTP
8ZNdkM8uPU8VrjjX/ZS10E7mpWIyMXg8Q2G3y/doGeIGfZszIxpophNsoCJAroF/
VbL6RutWrcMrT4MoR4yguWF/rMeVb+c+AW4lU8hXFNsecZ0HOe01/flxZ69xudEN
tv5/3Dcd4e31dOEUgMv5FAlPWE7sniPP3QRNrIEFPmgFUmCIban4wrhe3a1lT9KQ
TVGkHX2qDAunZ09pmg+K6yFQzIGppzfFKWwrIGPta1jO9vf3GUc/hPftFbdRPFGQ
KFlAVHbCqvPoIuS00aJ9C7QPTm5anJnDuax8YImdfR0iPF0IClPAIfZ+wgnav1oF
NxVF+Bvrnd5aUPCkWvN7rs0tru1TZl78okMwWexf9Z+GXruwYQAnKfEHTkmgwmF2
PQPeaJ1vB6gjXNsBn3lmhY6cWJvpzkqCJAU6RwI/azfznpRlzvAgUq/0ITqu6qJu
riKlCc5uTLB/aveXToY3Yde5q+t4Hftm96+dmvH/KGx9dWjz6Z7tOBJnlty/FwZa
fmllYvbZGh9n7EPQBEkgzG52Saw++ngVfIcbCxRxWFxe6jQteUV/hHDTOCTo+MLk
1TS6EJ+fTa7dfhMY1vItagdMgXe0zkxlI5NgnI8UisF3sQF+uhDo0ufWM3Yi7jSK
03Mb4Au2JfCwsnoTUGFmFLiA/u/Z3YoKTbqcSUpODMQndN+NTkTS+oew39UdzLIp
QhpgEM9K4w+YxVJZ3LEDG7XKE1ldrB9+BKgTjdBnioX7U1HrGOQpRgNQDfExE+j7
GCOkIlF/SrvJVO/B5vWzAsviv4qmfgcxM0CBtebBineV7A3fA44FjW5M1HanoK6L
bBhGwBTd17V7450fmyBEPmrqHT0CPm3bRlSwpwYoKKP1x1rHrrPNPEgs8MJUEa/h
4Ep2CvYu5bjqOX0NmEtPFrFkLm+jVs5VTcuhrE74NJL2OLSFAi8QSJffN/7YZ9M4
YdBOQBixcagumRNHsHcUODZxdvDFqnbub1/gDvvDiaeLxcB7EthKfe3lf7Zc7fnO
REHNf1NftmMJ3YosQxJ9lYCPBTAvb02NO+pgpqFmEAanL99s72DwgVy61BH026LR
4EWgBgoSAQ7xXS0sSSl/zUmlfGK5w7oe/OVrWR+jxhnhlhTp246DTroLfIrojg8P
BaudS6l7jJqlUCusyjv8sAS2hbNzXKibfxZBwnv0smOjcpyAfu+RiEweWYj91Pu4
IOA2z2VFPtV/gBDp75YD0GBUeNT0dmTJMzKmB2Icf3er3LXuPuFIiZRvYKEJcK3f
r1BUqpfx6JuXXPRTFvWwCiuz7fRUFUMXxhBOsgQznmYduNyyXyzbh9dSq7+X2gbW
+j/dKYBzaQWBCthAq7i7kzTC4n86kUL92toPc2qIP60RyyNPnBZbSIDHuYwr3pjt
glnuoVnzbftj52EOT/cyLMWQoEXh/bRPEz3FSlLUtQBZKrZ3fUE31GT+02XZd5dT
KTIT3pZMgsC7N+uHSyQFdAykJz3MWiHvPflIUwc34XtqWYSUr6/ncHgR4/Q99s0y
AxloD1poskPkDvDSa9T+XLtHBbcikqeNwc7c10LzN75Wl4Np0OKXR6SXaPhVUojS
sK+QGn+UjsXnQCThqeE/WtpeNcR9toaLKv78Jcbu/dDJ4Em1/Wo1t0qLj3R06lkI
hiU3StX9mOVSGO68NDxtcOQBbsFeRtt4L9TQPMCio5IzNShSRplat3+oda/rbLvn
4GsFFG68HBOcU6ON3FktjbNHvOtG6Ylf/grcp6aJ549bljRz3kDSurRxQISG5WMx
5W6DxxOsuMcwaPcPLqHc0E/uu7+PJHZF+zck8whHp75DbcNsOwnRvF0LFw7uNWmd
6AHxmidW0yDirn0/ITrBd+UCm9mWkwGPwEtgHjV0ft2n1q3eTUvh4LX9kQp7OxD8
naqr/6MFUe06PvuYwDXVFx1TOLEcm0FrYaxiNqVtJScr4hsIZQRQH/YQojh/KPIx
L3BnKN9479vjNdBnwOKwXNaTlM8IcTd7bRRGn+c1G21+1iIUG/UyDvIgyo/ZkcpG
l4CPwdodLk7Pq2o5j42pEpvlxW3fcn8cvX3c6dSG7V9cB67k6RrZLEDwiDH83Vgh
JRyp1deUmeiw81K2v6txQVRzQJHnBN3q8lZxPjsDdRUFro0Yq62udjfO8EZ+NCbK
LnEN+PHJPn/e3+iQlwMKT6hFQB9XMTaBEOAZO+ALfeaaQaFaOyC5mqVj5EcMJSwk
LYosDQWWwSmw/J35EO7WRbqZlhHMDNrk8/hxBESlwrX0ATfzXVfKDm61Y1jb05z3
tyqjfdqvGtwPVVjDeAcLnwji4v4AiEPFWCpX3T9zEPsoqO6bkA1GlCGuerZv+b1m
U3AomMVHDmaqQSVnwkpuWF1Agzat1yoiiXHb//zoF8IL4pBw5s21twqqcEUFPWWH
MgQHruq/RZvy1M2KAc9Y1sccGvw7N9gXDMFu/vAI66Tb6z4zs2DNN3gU0hUlP1OM
vGPHsRj70/cJ51ZgUD8xbgv9IZ5l1kJvy4kVbflZOMY+px/SpuDO5YTxUKd9dGc4
/Wz5xn/tB4G1Jbh0M/NWSvq5XeP3Eep2LnHd5IICWMnH9YR/gjfLydeXKZctmyuL
KH/tJvT0yvEzwy1K20YFs40DTyGADHEaywiJ+sZfYlBZ4c14F0ESq1+BhARXrw82
DTMmuyIYRsu9EPRJ7rxqMhKOQGxfo9TwmRtB8fFD17k=
`pragma protect end_protected
