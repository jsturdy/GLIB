// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fFr44X+iNzg6g9Llwefs0M5NR0o58Hhsncbw1zdcQ8q3pRZe7JWHaV0A84u25zJE
+2HOTqm2ikBm20Fq+/J/D59pLDOzYZzvP3MGBTtl09kmksqT8khyo89xAkIoKUME
bbwC424rlNrNVyBKuN+LZQ4e05NZTti2FfJKm3cTRm4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12864)
/rgMS0SQ7YDKqkTpjEX9+FbFrRaT44s5QuonIyTbCvK/MosdbGNleP1Z9tQ2zodk
M/mk1/Pz0b/c8rfjAxn7MkDLY1he+KIxTYHeXifGS0as/qCFRBU9GRl4YZBaUK+O
Rxd2ZdO/6bLYP0VZSj1OEvFyO2zG7L/yeabinZSs0s3dOrKiVCYw0neQg20+L4g2
ITftdgI9q6ayMJ8oNXNhF4UuxmxZzVtUfvCJaNPpGPx9xBicZkQlQ0USof3q8Cri
aHS5hkEZnBM1gf0s/ZHRhnPt1004obze+TdmmEB7vMl7zx3wDivsRCCiiUkHn6aW
WEpdObKHZm0mjgfG6TZiLKB7jabHG2XfEIE9He3zMez9gpsXIbmEOsxFPji5gzpy
8Z8Y8Mda3px0pQO931RwuBztq/a18xWIdzmgqUKjQozNR/xjYl1eRuCVRDbdsHUQ
S1Nmg4mJg/v/jr7XqXV27knoPmuZtjdJhmpCGe8DuVb7yDXCgj2ZodG2MxcmFWet
OUP+qi4KbaX9Yusm6nl7PYbyWCLYzozhBFV6qkU7C2lv3l0k4KwoyxrVz8cLQYBh
mbLVkno9lbINiJWkwEvnhnAPzPK53axBgSSuoW3lq1u9gy0aYJgvqi100nTF21vZ
4BhZblPTtJ8zPDzyixKXpwkiBumXQDoBWSTcf+r//j3jIocA15EkMGwDguiO8fbf
xkl0ONzJYr/f5ulxkBmBuldeyfn8PP5r6AQ2jvwM9eF3Xvzb/1HIOm675h/XY93Y
mdWt7foyvzaOb31JCTWAFYZ6R6Yk9v4u6jTrOfTc54xoLYc+NSBClu6dp9/qJc+W
6OPo9c69u2Mam+5Y5lbDsdfllAzD+LpncY5Iqed0SndYZbVMpKmJrHQorBSRxpeQ
/fHg603+ZA2+Xb1EC7hGtRg4mBcZm0XCik2id+MWlSgt9gRGAhc8Gr6uh2pETwk8
44MOEDdvCqyCU8HAn/hjW+bwCcIJSJE9MaANvCIOiIqCX57DVN6hoKgY/gNmUyqy
wgUuXBpq2yz3hIfivLKA9YDgsVij04mZj9DeORQ+mMPGF8kC3J5WeT6qTd/WJAtU
7PHLGYp7KaDnQHcWRzS2eE7dfbUJwQyYoZ0dWRt/c9VeOl/H/8+T9gX9j1KiYjkf
dXIZhwoOaiAIAjGjCm1tvm2fMuGl3VTeSdXjt9bqGRGsdYvr9ba/UWM/bJfie0SB
1WIqwdaF/TWTpSHguGByeLlDNt4LwBHGS19PCO4KUio123Ibiwb1Uagb+vpIj9yO
0WGf6QEitErwO0n6OMIDndW/3AJB+UeUnJZ7MRtrNyFCYoQE2ZyA0nvaKSbiInvh
HJi3hBwLOLdpJ4DBpcz/Ynw9jOZx8MDrYGZCUr9yirfOF19vGspY+8dITkgM6FR8
veaGfMO02xYoHVpfqLG3M3A0BYPlLpN6DI5G47h8qoYo6Z70mJap4/ZBg3uX9Q5q
5Do4suf/CC8xt97GjfPggq5vA9lfNCUYJR++vLHiQ1OclVsij4YcmearCBfaZe04
BK9RJk0bNI30tEXsXj0CIDtd1tz7Vl8ecQK9eDUIIS7Xcw2lNvGI2ERdnw15GtRJ
wZ5g47ik3UytgOgcJmYpzpB+rtY0WSceJmOX5DkR/2Fqt7+i+cTvW+eqnVPCjEt9
UlAGfwcgTecKDSGGBFDkk7XOI/egutZ1koX+c8VfSIbAWDN2qP3If3KG85bcKNEK
ZoqtCAd9DtyGUXq/NS6f50Lec1AdNTJjkO0EVFKunsClu8R2T40vaIzKbDH8zg0o
FkkqfjGxCH6GI+EDKUTUJQLiPbVSc8dIcoEEtwg5cm9i7o7Xv5XLeGNKQssqoOnF
4ISLXk0z5zVMVCCwjVQntQvCRUu2td+pTwU+r9rMUUjOQ9i4UsgFYsKjZceKPFAj
KtG/fZplxPuCR/k/3LqvpK7fQtYCIOiMm9LchZGPIg9zbCWKpg2fNv/6UgEG6c1r
AlRU/ynkuheOhtoa6FzSk6n1Gzt1W7rkeqVDib08Tav8NK8FCeMKVCzP6u99gbE8
q52DCm0QgX7IA9WL1CQb/zVEKMNFIwNRKEnlWKR3U+LSEUWE/k3OrvRaPICfE8Xp
r5Zta6yRf8u2GlnCtMXbyil7D7MgHhKTWEEqwXEPB3mY5vNslKq/G/yBE+1VowqI
VswbCjAffoeCR6Q/+uTtBNisIXn8s7ltLoSKkaoQ1MHRbETErM7hoEAz1Pc55tHQ
le4OG9g6GQpIV0aEIfv4ZYtsoBL7k8+6eMrYVXMSGHs98plKndmwwE6DatgO07zQ
7+aq5UXYj4VOKNkakQ/ZAf1bWvFvgU6LxHYWnSN6iJIY0bHlqEFUpXWSx5vhHHNs
Hmuv4YPCLmUT493UFZn/1i1OpCuRBJb13vWTNV2a1T+1/ec3CyNjO5tD5PCpBxd9
gAKEnP3Nb7zJ8aTneQbHS/mva0/JS6yqrUbpV8PYuErEl5y8eK28F4OXtV1GkQH3
F3NsmNy89qlbUPKmev+xuIrU/f84e4O7rwP/FLI5hITPQhEtnpkfRm50SOb6urh7
OP26sP94sc9oIiv6M7x4UaNymdwZ/V3Q1KvF15r2tMJKCgtW5k/3qz7z3FUnO3rd
4DDkzl+UWPuwC9vdKOnN6g/O8hbDHPzDPIoMoGr39RudYOnbTC8IBnurH3eitGeC
afFyxw83nWsCkWfsomHLyj2TFlzMAcZnB8eQZg6ch/6b0ubO+uGTTYo3MpCHUmZE
zq6Hllizr7zCYFPQFLc2YGMNIc7naT8Ef9cNzWhv7apv38kVxEu630kdu7WdtNMR
oKqHkauQZWeporrJ+Nn7py1gbDVVARH2dv2KKWTW3/ShUnAuXAX9ex0cyCuAZD0O
WovPEtHoy7R42hFUH3rKxlb5oDl7dbuIQuZCUTgR/r/SrMkd2DhL4FNqSXvvwzUs
Cgsv1uolATPF7Ma2w9azpziQ7szzJINklALIzu8XwA/bzoStB4xhpa5ttKooTYmf
gAgZUrgZghor2xrkQ94RlBkJPzI56mp/5FxosmyadcDJXBmxpIUgXauRjdg2zOoS
K5udtutJTOkUOX1DKC6jx6ffxskNIQ8VylIKJRkTgmo+H3zsYsIqTl5+w+JiLKFH
mrrWkVbt7dyuF9q5XWxyb9Nm9alWKt2F8R201eN9I2bjaJfU5yRVmTKvPK3XPK9X
a5uOJ/R84MrCbYlIFNIDTwnxr9Yd/+Di3sf9oG6BxwQ5cFHDbNQjByt59e3oSER5
dYp6zdMowlJrtzRxjBkmpCr8TDKdcvnuoZMwciGo+V2w1pZYyIFx5ZbIUksNBAi6
w8WplPmJJu+gJnI0jiWWdunyHlzFaYI6ndp6vA8UHgsplj9BHOx4YlqRrmBT7joS
0+1hOxqHkzZSX7Us7BCc4vgBgAlYZ3xYaIp+vLbJHq5OC5wAbgIzMsJdhwvChFBt
KmJH1gzUt7+xxkRo0owby+u4jy9+Y7jXTYcwpkOuRLJhRRy/l+EOXsiAYVbu1xVl
mbej7u0DbKbSb8I28g88utuwMge/5S/XYEMn85Wt8lSeAF1gos+dDn0/J7looSTk
6gDHTyQ9g83WEg+K7AtI0EfnIgzgr5ObGwMft42UUp8WMp+l9plQ2vuRgT5hb5ZL
LmlFxKBXsCleEUg4+5VSw14nSm4K8hSBnX7TaLBYrn3dnKYkBnTqTieJGBi3Sor0
uDwRXsnu5JJva7xcxghsz+HqYBbA9GBAi8RGtamgSCoUIBKd/xwt4yduyBtdEgtt
X6XSmPBw2kBB1sbOzoZJvYP49mB5Fi1IxEG5Rn6q+0xyJkl8VMQn8OuFQADLOfFm
sWY9TzBps8aezG3rD6emoTnPJVdkZRdkVFA7A8ohwbMKcyPlvf5sKWEc4S2Cn8sO
LsKDxzTE250+sFgjHnnJmT22Mf/yCw9ItT4Oe4iQWI7EJXFNvArgG48cYM9OVBHD
DqZdaK6H4G6/zD1DnGA6OrmvEgGqEx8QVM1Uiloc4irL/Qa6o0SxlbyaUxwggElc
zCxJ5jxcog3JGMs0YA70vC2IC9YFGs94o0NJACv7o635kgMSAx5TuGmxumn15y3Q
sN7Wr9b6gtO+cQilXA7L4OR/60/1lFTZ8vPLMOJNtlrLxXczaBkZ3PmsylXc4MnX
1Qi1/gOD1KyicUf3u583CaWi6AasoMo7lq6WIfUpOAgr3EbzxA12otMpPslaDEtE
bBQCEO0Y9cEoE05eRDwemZxA+NGyqNk2R0zzOPnbL+T1WNEtI2AM/+fTlEbhk2XV
V/Oh8wiF+vgliEgvCvpp3nuuRCJbyq016g5t28ShUqRCXrOmk9jldpZfKLs8VrvG
TQrBcWJWSstn9fRvRoIVi8HrSpQCxtGs25sEtGfECjUNRXV50LZrzWvQD0q+r8ld
UnsKSYOdKySlEidxsqBiLCjUQicPLfvFeHgZ20FFOL73Bvspd8Wq4hFW3HZPAO/Q
2VhQkWRQBbACXR9t9zDKNnkbt0WymlEfXBmb+5hsTLEDJyqIvWz66vezkGwQeqKz
EezHHDIPmx4zgYOiV7JByhIaxA6uuRltpr8//Wfj3ngP3O0t7GqlSftPA4vytj1z
U6B4rlmJjI4vwayAZnIaScj9xG1iJgfnZ4jsPXdBjNpQXTMwf9pikTXc3eunpwqS
KKwukp6lQ1ZHU2UM8fLYV+w3X8HGahq0O1rvR5ddsIoerI9TegI4C/cKNNwl7Jxr
KnIQJYMuWcpEZ0m3NlBBF/TYei88jZsYGTHGqpXaG7f7BgNgl9jSFZ9AbjGwm0ON
A2lLdxQM+7HxAddaRN9PvOF0rErw4Z9Q2JhfrEBDjA8Ru2zCNp+/CYMN0g+Sbl2z
VtSiiGTGYzqqbvmL/GdImAI9IESi6DJZzzzV4pBNxVZtiWW5iBGc/YxjqZ00n37m
f3YQZPVjcVeykGi4OxXyCwhPpIs/M/7oSF9zan5/UWp0LhTOfNmiurpYKUA/758G
gcrGXlde6xxmYEZYXk+uSm0UVKaKaZDqkqfM/nbqlLNl21E2WnA8ISeQC68yc+8o
bTi83bKfDXeAT+Hzhs7tugSZxBg1UrSXNevJoiM3b2ualfBgr6XvSmXL6ZhDG+FP
uG0k5dcsQpOc5CFu4KTga3fdjeEeXjDanRIVHOCc6pQYPFXVDZvbI7DPDDGhHrtw
6NFSAlVLAWO4U49FYBhu4ZWuK6EXGLGBOmo4pR0ONcMx5Aj67RNNAoo5NoCRkW8a
BnppLBb5UTRXJMF6IaOboJp1mF+oFEpoZXrJBdPqElVOznOyDvMHxpyY88D+XEZS
gC8xQkGG6WNcRqicuULGhzTTLMyzf7GeLv/HGU8w0pL64Lk7LgWKzEigqxSNWCCH
2nk7WTHS7R0Zm7FOolRZ4j33vfVPD/kujCqtdZ7IRC0twWM30CaqvLkgymf6ejIY
bMik3XGWZOyKhDj9+P0trp1f/Wcfow7regN20Q1eNu8hjLLJZ5aB6FwXKapZ1Ujz
frUrOXBWyFDCSLIGMcUwZ0vzKF8LRfMrJt5CNa7g0BYCRrIJgy1jHc436Usis2QM
BqCe7/1O+Z8iVxeI3IisslcRw3DTmTpUmLzf/U5Mu/YBIjvDrOBYcdlQ24l/0nGf
8ohzlTdqS+L9yQRa5wLbT3+n6i5Qs3slVKY1vsIeN4L9ovfxA+CPV53dXedhEc2i
7eJKxrzNgQXlExfC3mQON+iMBWj0mu0Yr+wjYbtYKQixgjmqMpl47lF6rUCsPieC
6u8lsWjlF/5XhPm8LasyrZLM9DCrE5i0xABc7tqDrQRpwn61xE5zLn3GUqpWJS3Z
I3WJzEbaUWVMkPxFcplrIeHGQUDIRVeuM7CIHv3lhNl0v0A11HalHQHzqqFe66a/
y+FLnfTofu80P0Cnu2OGQd08qa87hpzT1Q4YqB0LhIRG8aqpF7GvP+JNuszhCadq
H+XgTnYqo3rBhONjgT1HY9Zsnab+s/4wvL+miz+bQFfobldyZnfkEhcmMd+Tclfq
r4gUsYzE0HLL5uZJK0DBWYyaVjiOgtpwXd6r7FoqKZ4xxrkEMB1xeneVYsTTeAS+
RNwiJAknUYT2DcB7fPwWAaF52boQu3VYaXHZ9tTiUJSDkZgIJ0hfYkOtHSR3ea8d
cUsOlUrlgLc0mTLGtTXLid5s67Uy1/4jMtaUbREJfaprlKQ7CYBTEUksm8HiXpti
T8nNdvEQYOiprqdO5am70xzBGjA/oPI7bytE6jUQo20/Z58glYiJYuLVPDt0fI6P
6lzk0j5tnPcCrTfCr5CMP2gEQj2rFyUM/sjVFK21ahfwnQZNmMVHi2RcwGbE263N
r5uPeE6aq4d31ichfbTltuNrV1AqSw5lxOOG3TNgo3jmmdnJojZKo8UmuCyKSBzb
lfDdRNkq/0ASqo3ra1QIWbtkMsUxpw26nc+PLmRbrSfXZE2H59H7m/1CY3pRQwSV
+wJkpoN5gAGX6Z+pG+31pMIxLLrOEG/7MaOPerr3tYrPr/BZKBZBAaOefcutIZGq
KFtND8ENCZNY3AqVG13Dqy2+0t2yNOe+Y7Upq+TEoLj1sDH8q0QVUvaN6D+yC2Wn
IY+956vSyecL15yNiMmj0ehDwW3RGRDNKRRMb9NrRZoAB72pIcvFf5Lk3oocx9Jo
zod1uSeLnGSSQW5MuWH0ihyH7oBKBK8y4k4jLs8oRVvQTREhczwkDnV+WCq4oqVv
nytLE2XRYTYJSvG7QTqmLwP/VDlHl3dXIOu7kyYN9FrVeVYd+Up5wvOKY96Q/roi
usvPGZIqJeAFuvnCZDwINc33nYKCExaJ6x9pCY1FEQ6wMhlbisrL6oHhTOUUClVp
4YKIZlolffPE3cyc0eV0KdcgKHe1YS2wMZ3BA7XCCDZQUrWeMjrO8yUlogVXI3jC
Jr9ezRxpy/gSgOZTWqp7mDupW3SCe/a9PF1TyC6uNTYV4UGJdzH9Sxo3H+4eiGcQ
nKhqCE0shILWUvql0NtHtctV1sJ6r11/xPhsrES+Eat4H9rgtNNRd6ivDNiVxEdk
RB5TPBGh+8yXbAtWekaYs43anbGHObWaTz/NMNC1nG6romxIVYMTn3tELVWUryXH
WTq3x951r1rBoxKV7TrXy2NQN03XAUbfrGy3mzMUG1Yauhu4gfckL/swN1hAhymN
Hx4M+3m6W8QJqJw6gZxE/EQlGe1fveXo8/5G5pfiJx9oYzwwaQJPZ2tU24Uq9GYV
xTA2CSZaFSJ7eWJXxaGJT2W9LMzqKQjzGpSlBX5nF37dp26hIvv91CqZF6T4jWg+
ieRnYPgae14ieAu6UdEdZXMi+U4hOoz2GLPk8uaGPO7uGzimQJ1VFL87Qu0vI4hV
AjZ/p6hZNWYCZrUq7s1aMUXp57JK6t5gg9DnrTMlkMU0Vf24ZXg450OBi/LlrssS
LgD00zd9TgGSx+iUpirZXsbFF8Db6Y6XGVw8xrm5DWBXq0jfaCaRLEOdNlnbkIKm
D5pieocYwAWWpVjLDNG4cDMOgJ9jYtM/AyvutvDpN5AlsX5qdNV6NA5VY5yCMSFJ
V9Q6CumFYPebaM4JW5LCk2Hp+scLhGESnYxaWjU6TZWUNw+XWqLrp/JSjb65JclE
Vu3TkV8OFIo6rGGedF01u22mK/784gX7x8fNbNBjBLFNXsxSLyfdVVnAUXuY3+8F
KYRczIMsRHHnTGq+ZtZaE+gUemID8+XkYKKx6bgOaKMvFmDJ/K5pfKjIJLtgSnmo
lLMqbdtuFpqgUoZPS+KU0KqwoO4eS6lzmf5c7OdY+gY2mn/K28++xmlPH77tdwWO
aB3DY2+x6+o7sRxE1HxeOS5XETRrQubNtP/9i+idakTfFI2xlkmoeqjKwGsPQhN9
gpGIuThDsSr6YtqZ6FIpxSW4szWk7o/Q+JKanRckyuAa4D3U806+NUPfHTGBsx0n
3QJZV4/F5MtXH1VA9LJXWy6g47kdyxsZdZYERqFfLraXe4Ncbd8nAb4ot3SCGLwl
eHnIxqPq+PSs0R6js+aPOIFWDJqNAaIKYtbQe6PmS7IjBwTFm4tCNZ5C7lZYElWl
/aJovxSmDeZCjI031x02FC7YYDZlRVP1zwZSX4URjFlyMyniBeKl0sc85dj38fiv
71Cb1JMLRBtU3/O/olH7NEj169SrXuO4IJEMC1L9btwojSC8rFeUQM57vfyHV7at
oLMAoYWX7/HuXnDC5TZX6+y80Zyev1nC6VNwZk+ZnPviuibHm4jFkJ6/4zcpxgqd
siezPSW01GivyglSCXP3cvWRptU8AehG6suHIwV+aoWFqyEBasNnVgJY8EjrAp72
fFUflrsUQ/3aHAn/K9SG/E/ljpWEjbU8o3M76dK+JxmzUvvZFOOkQgdRko12sGBK
vW5YdKXMeqc3RaCn0ungFVyPEr/9kTO/ke1Z9dtek+EObGVYUUvTtYtr3Yk5JtKj
2dtK8PI8Zje8h/GdmzumzujSpT+stGI6PsovMN98ax4No/Y69hYH8HEcG+aL6D2J
cTQdnrW2ogN+MOlpwM+uXE0wlytCU3Qw5986T0gJ7Yh+AjGTOzGc9KwRHADmr9Cc
lFOd8iZbkDKXochuzc6Qi5D3X8Hh3c+zNvf+XcpqkN886yjjFx/yUauonkP3XvnW
ckGWBnDMxyMGf4/uJ3mZMyiXkv28iZExCRffKYm8AExMKmcxpuQbZD+/PB28nqTS
nqUUBi8juStggU7h6KWw9Q3SmC2L4VyJKw0RnpTRLbLYOatjFYWHhbKVyKSKVaIc
vPsV6tnCDdn97DEhWCw5OVdsZxew/LtIEfwgVLXE0A0Waei4bpevxj+AyPCaMjvR
LYkaF9TdBgdcCMZKKx5sEagBvLr6ItnGPGpbTSpthr3grUVw93X0kFEx2euMjv+I
SfpFb0wJ6tmZAY20/t9m7QhNbWaJLtVXFX/GkeDVAmRcmZ9dKNjozdu66bsPcqj9
+kBit8NQJ4DIX5MvT8A/IO7RT5mAXVK2gfKPOXTjoYmSAprM6fcVXzDajcFHMOhU
CVka38dU6tN7wrxh5yvGxFx4sdsxxW4qe2oTokwVMVVrixh5mJw49IeBgUwdRUWo
+57U+2ymvm9ZpPUOZyHRUOpjspQyyEAxrjQdkGrRcp1+G3GYV7WzBnAY71q6y9bI
+A3JeqsHn08JUgorGwyJOkFQYNbRE1eL9BpXpFzBCDqtr5DN7tFG6LkTWb8yMg0d
fUbGm2eV0lPLV2K8ZO5Kz2PsMjhh8kE+4FvvRe+0ChpIvkDdE5HWwzXMWcGPYsW7
6eL6wdcKtv5r6Bh5IGbvSVcuH1FIOlNkbiVwmTmOwfEj6y6PQPPuFugPwc/uLuiZ
sYbtxaq3CSwqYwu7mCZpNaIXLnrJ3R/PdML3jI0X8+NdVjgqOjuz8AHpY66eC3cq
KDhdbzVKUHNEW2+KPwvkPcWnRsZmHJSjBwdqEQUKY+CSjefX+3OvpaaBVylZ3MKG
33qhTSknmdf2ShkjVGsn0wCODIz4xJSno4jDH3J2tbNRY9G5PA3dm9k5wLb22oYn
oA7DYt8QZ2GqiJdFE+32pPKy9laFi4d0TFFbow9XM2aYHPU6mmGqFwk37aQDuwMF
7xjz1Q50fCv8wNdCEohmCYAjlQZq1bNkdnIla6j8NkaFtXG/bS/yFod6KWPDMmiW
2oFFrL65mTL4yew6m1p20Msqown6q78iZJP5MrwbgMSTfDtCHB58cpXZIfk1fdm2
GO1INZFBhYcGswjB5ecRlCFLOuTaFobi76WimF8mz2AiHHwPyimyY6ToT5AbNP/i
5pIaLPkQn7Wo+vakErU7sEfSAh8IR85GF+0E16j4J9DwffMrkQz8l34GBOdOh4+b
1E6ae4I1cjDt39/MqjqWf3hPEGGS83L0Fzi7sIQJzI839uJRr1sOGG8wHKxx3lvt
AfZK0MDIC0IQgMfIinTMBVCrSOrYCiCqzE9bJppxzapXX8QT6Op5PILkG7ustKTL
vBjODoKKB7Nb7W+QW5j7Y0EDqjN+VQJ5sZGh6pnjOag6tqeBHRqQE05PDQvsniKF
t/40XsnAQ5cztv1CcJvSnszguDWx1ZALcSTh686pcquRjXMZr0ZxXuXwVNdgzRcN
y9k7J7ONW3G1fDgGRqvJycgnjmDNp/CLGrB009izSIOjKGZlQ8E/2mL/IwWBX5ti
6vS2sbd5wn2bZvKFE94Zkx2L4NTAByA4rsvdnWY7/k3b9pv7zjf+E7DGfwFCy5xd
d6DY9BIJE0PBKiVoHC8Vy3IuMvgRyMsOHLqWCIVtfnkS13X98THf+HyokBZ9tJFe
e5VKpXCLHaLF5lH7FWJg70HH7xoA1fBXHrG0BFbt3W+Z9mlGyJrg1D+xkEzCG3de
eQW1EVL6MH/h4xsdKh5OHqFD+caymZxyZDgbnT9ZMVGKFPWRXbiUUxLioAEQof6K
1pLrrnBcu3QhqMKpisKzywBz55fFPP0aCI5jBNOs2C1ckTXwH5+cMXCpAnvtZuRI
r0PuvnL+Na53mWbNAuIFnynq6qFrNqB9NRFwzKzHIgGaH8IwaSJ68Xw0Lkt6pDiq
PHAUDWFsNcS0BHBldKrgPN7ebSUgl2KHqWkHy30cx0oAWmzugXtYYJwC5uLpJF/u
iDhLGB+iiQquTzfM5IbzvsLgmz2Wvx6184tCiFb1bb4yUV4mVOImEwuwF6Fo8HxF
VbdkzD/d121Sp7o8oBds7bVT21s2qw5HJ5mVWu62SCRIrL9FwldcoXVWA7SgJgYQ
kaO5pqB9DxVhJaYIrdV/1AgrhwScUNy030o2WI/hidKyMIrmYxzrvcOTx2VJv6yw
mI2qHPukKuv21hddmKnrQ17ABRQGDubsfPgsMTVmwteA28hJbl7g2Kr73hfDNpf+
+XRvxy+NjxqwVYDcyVivtzpMmnghPDe4LTc/M6wBfYAK+z8DHH35ogLuA26go2oU
GDGszRb9R8UYTzR+BiNp4Y9HSKh2eAvAIW2GZ88ypUsouOLBWnY67vjxSasSWNC9
6X8Wkt8sqi6YsW43D/07e+wzXn2a1tPvA/WRG9PF9Q7Gx6QsU3a+lG07X//GQhEX
VNHSKqLhPVYRjhOfjgtPaCgJuGBEMElKvxZJ1bqGc/RNj6Ne0U8F8onAZ+wDiLUw
KKjWWuEeUNJAAXFDZ7raybzj6M5Kmw0x64u4rrqFZ1UNcDSYSKaCKHrMTzd9dZL1
IWebD+CVG8krkFKjHpRmn/AyxCAfD0ZwR0PIke6Q7btsWZ7ByZeYkDMKZe+WrKus
Jo1UbRWqAXdcyLzCCJwUbIEfD1x/0nNrQ8q9/DP0ep/OuiZ+crwN6KbJlIJv4R/F
UDZ0aXYKS0lm/vHHPSKmerrb0gPvF7SCxJ2KeQV3+MVR+vhmdU7hShCMUeojbktd
Xu0QU1tFlEF6jZax6o41OH5u4CXPCiXt24liiKQPu6pPKhOgFNZyc/90XFJ2+BRx
Ccmfqh+GP1A+imyDd/sv9MfHraXyc1y3zgnjYnnhnJk31rVvo8VGspPfYDVUVKa3
Je+M3WdlOlxhfYr9+65A4dC/s8RR+mdpyyYVpSnDz+wg/qqSLjSif5mJRojQXacr
Pq6wPVaiuw30m6CQ+k/vAgHoBsR3vTVjSu+u5w5JarH+dxuw6RLIomVnhHAkMSvc
M1E3novxB5wa0y7/Hkt6vAcvJU2Kt7i9BCn5tuLQkG3V4l4m6nX9+xDQnu2D4ax1
HgXU6kchWbfws08hXgsoTsgeWL4Jn2npQdW9WiMf1l1yNUN8h/pj1Nr4d2GShyYN
BHcsiBy3H3YAtQaU4jsyKFIic4HayimMSwe5zqdIxsM7MoSFL6iBDQmDNtILBvFW
tBbnKeQwwlnGhOZDBjB1yrYvd/pVhJ6sRTDWplcdshO13cS0TIgaDHyL6U+Xm7F9
at6iRYI9brWou2d67Y+lYfzb/cUzrdX81Em1u9R/Xp9MXExqQdlrQt7/yN5SpLZp
qEDExFsWIsquIwQlTSAeb61qdcvhTdwSHBFFxHspATVGshelS/vSjpb77yRCPIBV
fSFkaUP/RXHvQf1NLJwSgtMY1+h4wx44XxdTa1F1VR/98DyeifA2HFsPXTXPf+Ib
m/Oyuc+ZD9tm1Es8dBbUMTtAjdSYCx0Lepu3RiyHD89szlDa4J2MpS+f8wAQZ2o3
uoQacI94efpDcz11C8yiUTq6D3slriRKwbReRyXQu4NCO/kyUPi6DJ7eMdU111uf
2JNH5G8lcf4n5/B0loC0PTKDoIv06Khm763TnaLvJ5ibu3Kwdr0g8nKDpib5yZDB
BnFMdy6szjp3A5TCeMF37c7OkP5CMTI9/e9pDRmt0n1Rpkb7Cn1q2GN1HayKy7dx
gz74S1c7Tvq8l46dFhc/nj35Mj2Vls2UzLtNp352r9Qlj3rsdMlYbfWjDyxmzWSy
0ztkvtS1sH1oBV0e/s7uu7PNFrsXZ60mOcduFLMAyLoFtwTdBtkb1t5qFyZ/DdF7
BEAJNM16dbRYcor7LuFt/HZe2FjwoM4x8zkx9epbgkcnPi/rFm21HXCFSBHJ39LZ
HoXFCyQ42AMdy6O/qzILOd5Uie0Rqk6Cov5sTMWGSiUMbYCey7qmnVChH8Z68/GE
zlY+Sa1nhDCkUIIhDY3TAZJzgscGZHkwaZEYwBWxTTyep8AooScCBmL6LzxKryxj
7Xr563COjC7VGV2cd7UVAyqn9RX5YhwJ+BUvNeD++LKA5w4XdrMTD5LepxECjzjG
qQVa/Z7hM8bBvNz6vDabJqf1WBG7ekkdCBBOYaEXIcdgvNMQYtDskVsjeZlFZvkz
giVtFP2gzL6AevEDcPN+IkobZiuDYWq27d10uyvw3njVDG/OL6o+Vky5gzH+Kg/t
5UgemJ6u7mWNulQrCJHH6itIO0MJ0HY3nUliqOsmK5FQNryrXr0odSHLC6hU2grK
eH20ZfSuajZcbQ3NMbUO+dnZIkZBfMHri9kCF84Pb3jNx9Lk32q9dZ9KjPZLS1Zz
u2Nf/SO0LxQNRMkgqCDeS2u7l2Z6CEVIqSjh9E9rN4gUBAw9Pu6WXxaqyntrsFUn
0MM5XZOkInpwK2jGAn+V2iqS7CTsSCA3uG/P/D9wFuWkoPa2Ai48RYRPpwFqaIft
UK/joD+NT0R+kbHzalROxkSA8Ahczmv+fb/NkLUKUbbdX/t7y7aE7VnARrM7l0Ux
/Ap3DbqtU30bRUvv4Tu5lAFkMOvDL3zBiW5YsBB3FJ11RcaTq9hhLbVMiXBq3SVw
LvXzFIJ5JmzlrzLCeVSaEfGYSAXwHE4FgnTcAAdKP0tK5PryUnMCrqKPxaZcAZO4
vf+esJ6JGmu/3Op6il6jn7lZuYUP7+VwuBkTG8OlLjQGfAVjEQTI9x2jcjTe82ZO
dcXvQzFD+/QGnRuH7ESwukrjzlI6IWLR+cB25AQCx5YZh7W8Ch4KzC7YK9XpIbZK
L/ZVghsh//2u70es84Y/Mir6iM0Ffa7u2otQ4dsukJQ2gunMEqkzkK0YJzY2Xl4T
OyPZRF37dM0BE9IqCgzdxTq7dvXAtNHUpaDj99dBfe8QbjKOOAQkg6tvndbN4H94
ohA3WIoWkB4hoynxnErXF9nvCpp+UGi4PqKTXwVXCZHMcjgHHon4xijodS1NPrLw
CkhKV82pfb9EifHx6d+It7Y1ciRXGH+6MHiODDPdKWzx6YPx2xpcuNtKZukkgwDw
DWLUiyKUoFkhJF/dqVpotQVSHjz1Vu4jlg0oO4RS4fS2NASUvX4gzwY2B9KOZuSU
rqmwe40/89DhRmfKdZYCpXjCsLT8u3RwtQRQb5jJyfnoIGWjuvW5zOXj3VLFuTLj
gmmdEKxH+26ZtbW8YF4F2yutRa7ul6bIi/ArdS4CKJIN9/9GjIi7l6WRVlkJ3Ttt
MgxN6GhuUZpqsiqXkC/RPnWeuvM+YrtU07bFXkAcfiRtNkjc8GC66S7iM8xh4/ff
voUHdOKALenHrE9FDc5cRS4Esaw2SFyiX3gh1iye2LH2t4ZlPWMN/Prlb4zWRsu6
poI/LfPdFkn6yE7eERjO4LYep4554mN5WqtEqhSA675rEWpsIZmGHrWa2p7fVbXt
fEHkq8I/KY2xa+zh67cCPRcRyBHF6lfE2FawsTUF3I8qst3gNDnyw42iYWcAWasY
sr4OuwwGJXXLRz3OxaTRE3ZQnNsqam7H0rrR0YkGXO95JG25s6oZC5n9DopFs2ps
/WLMsjnVfW86JEdLar0UnJIiTzrcKVSG+UVCLbOw7AL1bxENYxrF8I7GD2RjPjqN
l63pt+wkDT0foxtDvCjSKouIVXizo215YtJP8WETnz3zBtzGV+qLS+j8WdPk1Pmq
0IwxtPpZvh8ZElFmjUQKaSQGorSc919NduNTzbmzNlUg0V/v8NtzrjXR5V/xSepz
WRinWGMIhD+WEqCQvHqSQD0vw3oZU6pOZL1UEFwUJMX4bLObUmO7eGAK1+YWTjDn
6YyAIE+BaLc5CO4s37UqolmSHZQVA3b52yFHnsIoal137gt13v6bF151mALDBwcl
Y9e51hWXVoxGy6EjfLXO5QvxMBYRMwzOYXmryTr5eEtoR+Smk9PrK/h4hzwEwkFa
xGCSaHiub4PmlvdIgOP0Xz4JcmV3wFVdZCBFDtwj2CVtZde+oxBMmiTlKs36NEA8
T7euaM/v5oA/P2WSo6VM3LxGAhDSCUQnomrvzf7DUwSL+HDR3MECD+p9kMRjDq+C
OJpNBAKhQA4bL/m0L2Cs0Xp8fhxHj9iQ2qP3aRMhwRGKPTPowrDkcbuBVEQbJkUi
vTalMw9KQHY6xdafMxk9xuTOuj4EtsvZIhEd1XCman70K3f5peFWFHwcFTrf6Lwg
z8xs19GI3VHeRa7dHnrd1Fd8XihiAtWkLtkSQqD1cR5emuBd5kMKYxCdrq8TrSES
8JXwnw7/S6+h8wVVyICqpeFnLaLuwWV1tVureVYbnqVoLAs8LHzEJvg/OBdI43Rv
BwnBTfSDHjFmiq6lM5XguZVq9UGuyq4alYyf3xTCIP+4sNy7VrAUDh4ifd9b4iNI
8C70T+cIieaIPC/VwtmTSmzGOgzYO4HW4/ejzl9gY33J0Mr5g58hcIS2MfLTo5Bd
mkteEmDundd5g141K7aCdJBcMsIgwBub7i4eiLO1aefT073WbpVOXLA0bJRGzCCi
32IhaezQs5wqJn953TxEP6kS3H4dHXq0klAzcRMKYwUDpnuFfiYoWYYjjVNe5hup
k7ABuHeORhBru2lDM6ssKqmEt1W17gOQw3gLJWruyO0ESHicZwE/SADOzK9TNiUO
fYkx9HAcKtfV4V1YPy45L92jQ3irsRfuMv+IQyeMS9jv9EXqFPhaDeOBGRI9UbLB
OxVu0sY93BVs7rR+WeGME9r+ynXvUtvzJrYA9kAr13RubzE93O4+kL+NXA2w/qGq
Q9a6zUFRysZQdlKnho3mz0/dQckq1OYrhudftj7sHAGhY8h4DoT3gCaazqEIvpBY
9c9xwWMqfci6xIgS731/AT55Wwo6Tzur6xr/n4dv1N4dsXKvS1aBdblRXc0ekJ1v
+R6gluxti1uPtFyrvN1vA7SoUmO1qs83HJ1+MckDm+kYedxn9/DRSDQ+GG6fn/vX
Y7g7C5xMlQz/rdg+i5fFtpsvuiLnxjTBy4tQxbLy1rH6hnbV19xLGBSj4Jhy/3cf
IY9RGtH4Ai+VPdVWj3h5YcT+TB3E2cX0q0CE/M8pJVFpQF9i+Lz41H8VcCFTSm8p
aijdqX98csKFcDqHpF+BQIbLyeA2AyuFE+Tq1CZjQe3Z+hHSDxYOsbys5mHkwK3B
OQWNQPH59x6jDHwb21WBDEx0pShgZtyJhc9rbp+4bzvVAxGP7xUELbgcmsBLj/cs
IfsxO4q2PP0C3qD1hkYLYUcB4e+WevAqVd6ONtfJXeUamEDdLXDmq4iQrTO6w6hI
nCRGTK+qODa3vdi2qO6ld+KeeDZe/r+XleaTIzoNt27GxLo6uXkyqfGQ64+v2qUx
uGjDIHhXERomM+rkhkd2R7TXg8wFN6sBw1b7guD3WKMLKb5EHIki5XN+3h3z1WcB
LYBAvf7SLpI4vpVNoQvdIaXwnb/L55DkI1DD5QoYEsWVqHlNpztYMDuBqXYqBP3c
Gx5bWK6ERc+r+NiYuntSX5rwSbRd6GJYJ8vqtrz/vdjPj15Y2FoFEFGTmub1LAC3
vp0S6EVEeHUpjIqHgtfXlm8xO49aHz/r7/4kLmyaL9MXFoVo9Z/8O1RemSaMAwU5
F/YD/CJp8DMIn3EaC+SHyt91g6d+4C/aRQEnMMrMwqezpm/CXIGljcygrpiXwhr6
TyF3wHgx0yg7efBrvRyWqivF85eX/RF6bMrkcjQPYzrz0VmHpvXy/EPqzNU12aFY
V7N3o71L1ZEikbcRmW6Lh1D7VwpOKbrzJO68cHt6oAYO5D9qgKkbV6vDMbYdcRGF
pSIcmQS3Y4StnLt4iWLcGCZFVtHgd8gg3GxrQS2Txvqy/CvXFTBVPONCQdlLufVg
W9wL2OwiluYzeKK7cyPlAKMa7CWEm/4Xof5ZohyJ9ZacoTbJBdHWrkllV3sgz5fh
mqEIaQiSM6n7MihDinJgfs60Zkk/yPPhRnZHgSKA71UhFxu0CJXAP58n5c1GniE8
bHXC5t/ANyED01TotZPGhJ+t9L0smYscWUq+0nWh1aomhuO0xLy5FLhoy9s7f6qL
Huff/FZqttGgVAD8koM3sF+Bz4NbNX7TLoVYwTw36+n5Mc5b1NNxTZMT5xoquaFF
d5+BqrsBEEjKce/BWobK4CLNJYj59r6QxQ41XkTpnVwps2gfT4xbtYQOpwMvSEuT
9ptTV2z/dg6xtDeXAfPcVwobFeiz+9JREXP5gvr6F/zKvJY0+gk0xfCj12cFTp6T
OfRrvDxbYoQuC+QpZWthmZ1KR+lbtjUUOo2YNYHS8C5xw5zIC/XpIOgIWHjTpgtQ
CQYA7F7flRZYHNgQB8+S83c3kfTwCdAxqGihphZ65Z3CphEWYziTE/0SusYuqO9Z
T08q7pBypemgEB57OiBC10NmRUhdyJ/iO/ZzE03DO9IRkGjUlcld9dbnpaF02Oya
Ok1AFCkY5UGSuBaIioBJyDep5bCb8S6EphUSJamZl4npcUNS2tRNQYJ/UM4MYNv/
`pragma protect end_protected
