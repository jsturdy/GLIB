// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ePjSCADNjIjy0L/6MTAm8cKicu6c5zYaL5/8RWT9jKLobeN7sLFOE8MBThxwIDM3
IW/SgB6h7D0nuY48IzaaKqQsF+wyb/9erSRtPh2wXoB3t82HCK/hE4pwaV2WaWOK
ILoSppw/41B4fZaU5kHbew10334FL0Ky23lndouDSUo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30176)
Eb7+DylZ1CJDGon0TAT5YCqr9zAEqGZXwv0icLn6WiYeUWgtkX5iIJW7uxc5EumL
fmBKvJARKp40ozS7jVtZg1Uihdbqm2NZTAF1/H9BIg4cXKTZJ/Ap4W4scGdCRFc6
LvH3zfUgfP0OrwsjRMegv+vzPmP0QZW+7AYQXePTSkMRUUsbf7kPacWhyXff3oPm
m00uzTpg9eiN4FrM5MsYCwQRkM0+piWoNtiR7CAuJKhUi46F+f/PvHS1739sW3KJ
+A5143r8lFv/wGBgasPEcIaOid+5pU+8yeKnw/dGpuWTXm8NCL1Ca1z/VEOjksg1
DmBzel3EJsVQpdXnAFQAgcgzeZtH1C7L6nnKUlNXTDyTAAD+qz2H+qvI1k7UNkEg
pKG4oGowtHKT+bnKPxwX9srhS/9fCeLrbLQzdDgac2wbgvi07pBAmVTeOwByN3Nj
iMNyEHGVyoLaOdVFP8l3bsmDAK8e0ZbF/86HHPfDl51tlvBfjMXNyLWeVMIWW7oE
lqh/cpmrW5AFAfZmgiBP8gSDnXp5wXLfAozrwTzOuYaqxs2sKhN++F1Ft2Jz5LfY
hHcF59qV6SNsoaJ9s+1GLBUGOAOydfyYf/uQPN1WKxDzKpPTDv5/hONczNzfpd9Q
ct62e0rDUUTdywjA2Y8LiTf03y7uqthYgrgTmcgezpXqN9E/C0lZw4SKTuWf2XnP
kOHJIjD08TtHQDV8DRYUGez9/zzdZy44PEblCZH9Y6nVqiA2U4+dkrOPHupAlbbr
ljTgfttFHtILheUt4fqhkH9pHk/3OnwPZPQLhNrothcXz8aMVdqgrXM9lBMIIesX
jHoLrUVH4Qbt7c/xkkc8qcslhBfKxrXZdmyVaYjl1j9KmOqdrOG8Q16DV0c+No3h
2h5Bi8Ipb/URLYKQ1trKYtqP0gVFyo7Kzbb3y0uqi151VpeX9AjDTBqGLPWfL7ND
b4ETSpr2qO/u+wlQpB+xv9CpkwrHXa+AKqCzUDhi0Fmqk/OopaHdCkVdj8OTPrx3
BqsiiU6lJxv+eFANS1oUgujY3vU1j5/b0ehXDvKyEb/741hAyNkbW92HURj78j68
ShWocd5Z/A6kfZ7QXJ2giZ3VXq9CEngduFAioECTdcuewx6wmiXQHoeOl8uVseiO
KzYe7gf2SI5xgeYY/U7KCHeqUtAYvd0ii5IjKT7KQQGm0i6aTMta49G0JCsm8Ih9
bMPwjNfi4RfZOP4O7XBT8T5xPqRNKc9vw0jSSF6bTaymUhAdnVZL6b5AXZNbrNE7
2hLhFzh+/aOwzJf4EQdBdNvZ9qoIki78PlI1B6mNWhtrKqq2BHn/yGqqgEs9iyze
raEvY6xE3rvzuSS2KSHy1tooLyssulpW1pwBkgQPxWSwUv+FRHmR15p8WlSA5GRD
Z1pURKE31tLhpZlX5GuWy7MZQzFburq5uxCWu0xvmesuylEuG9ek3l2MKk+ti3qr
NuThtHZQ3LurBe5jlIzVFFxcgCykG131QIWcVBxaM11zzrOZW700XmnU1LzzzN+q
kMfL4nXFUxWJ3WpY9aLV3n7BBnmPRRR1UA/h7DoYWvtmhu2V9OkX7kpuczJA5wKG
ZvSnzsnPU4cnwy7/w71Ql5jWogzsEr0SAz/CHR1JPAO18xFnktj1Dzslt1YT2IgT
rN2CsYTr/DRI4WWW4COhevYU+jWKUo88Dfr8E3G7uBU9uNnDJU7KIweGkThIGFuI
D2sQuwRF3d2e7GlfgJtEn7PKubqgMQJgRH7pGH/37w05yVhdp2yGSwGqq24I6n1O
g8RbvfsUd4AtrcZfzhNxAyrCPVg3cOL/mcigCwNASKRVjs2GEQHGCrRiC7+p4ePa
1ku20L/Cw/p0azVTlBIAp76fEnmQxPtz0VHLeTHZHaCIRnnCELbxKevvhqym2qDB
wEZwbQfV3f8105Pm/oBfZQVOMUTbDntOJY+5nfQGfhusw0UsaH1RF25eeXhivzsk
7W6cYq8ZYjW2J47yWILIdNbLykqTLlTJxav2r8kptZd8yqvoCzJn93xmcwlss/dU
ceM4+amq9bfVOgjHP7h7WbarSn5DUa3v2H2r6H1ABgo7649L35K4owljIxqFHpon
M2zKhotvW8n9DA1/lfy6McC7BiPGcDwAX3sfypBzXKYwpOwlj4qEc9SDqZ6LLgOF
2AWpIrMZSF3UCr1o4jpUfrJNYXInbzCRAM8V5M7ELE8sjSAY/HSQUcsatHfOXufN
ezyjX4BS/bXW6ibd9jKBUPZEG1FuAPFCsASqwCCgX06GcVKTL7uUFzG9LrbW0zjM
w+AcyG3F7DwQO1UT1kgyO1HqohW3jZ+45WxaYwTmbyLPokd8li7jg2caeK0ZC3JY
THS5Fq7Q5+rBU9ZooXqWOFVwrl4khArwokJPlvCoTip2+5gQbIqO0Z38HX08ZYat
py3zakd2HgN85QHgQ4WNLebuLaHu8Ha0sc4sUsWPEnqIjQCiQfAEvOMmw2Z4vVHS
NEOjJ2ctrIgnLdS8xk0xMoGY3dpfVyxgMv5Fcrt3/Dtw80a1Sox6l6sxLQCA9ofc
R41b7ZRLOTIZIeLCdveqs8AFzmyu9P1AqW5TSpCBKo4tAKQk0cNKZ6oVtLoqUI50
z0+nz5mvvIZcdbE7Jl6+ju5l6/guFiOIgk0oVT4h0eAk+FL6h5GwRx65Uu6xdhD+
MTPSKviXdcKXNkghYsN2joQxRhNwFjdkyg2ATafXqxJC7VWwrMaW6+FUqRUvJiBk
B3j7i2SLcek+spCCFWb+W2ACJqxZG2DZ6qXf4wTO8pniw0mRRgCtngNdY58OFbvf
VBe/XQ15ydmvubD631shNd+fQsXnojIw6jLvgA66LlOcGFJCmKzIlqbiiKN3xS/E
Ixf1W/iQXfYyu+7B5g4OaSrLToYUHdCvgAnYNKToL+5jyUr0/Yugr8Ui4KwQ25Qa
2Xsn/u+CB4BmdWo0uHzlbK/E1mA+Hl0ERxwonVL8Zsnabgdr6AaSRqpsUQcuWXED
rPBWLnuq9HgL7WZG/FiD+Q9DF03FL4AFxva4rbqPnDQUgvyG/lIFu0YBrZIHZRbo
dTtRZreW7c2L2BtT0W+OErR/GblUWhHdcN1LotGazRjr2JKKqiRadOsz55s8DQH9
yRvCmitNXfAtSaqzn4wC7WkXHqXtZ3vDUAU+w0jy7rECrC7lOTwPdOz+b6CDS1px
cNIo6jPdD8OhHs+0xyYrw2M9tr8knVYUrsfmlfDyJbBF4iC7t1x8SlFW5P7XTTUp
tuz892DxsqJMavu/GDwk/sMrhTjokUiquP3kcbgdsXyqftK2s6tlWRvc1iwyCWd7
BKKKsZnyYACUY47uyIRRSxboZFaCFwS793/AQZkVLeTJ1I43dAs3XrqxsYBNKvjs
UKyVQEpyQycSswva4bg1c5BtntBSndryV1v6OPF+y/l2PTLf3kX0LVJEOFJzxRaA
+ZnDKXLc+Qf8dRPv8ph3HDj/zC0iRFr4OtjHo5Pdo0yCpOQu2BKFYJzazYNAMbCj
gvYM7fgLVxJjoQKxCIuLUmT//y1c1MvEZa7R9JGLhFAdZ12JL16K9ND2Cv+q/trA
nGclTAKwbVO1PCT9uOndBZdloXAvx7eNUlAifzGOwNmdyh2myl52QP67LblaPD3f
yEKwmAZXX+7jULAs3NYmi77d1UKr5bSluHsqrd60G8QTdigMjI/u1v5Q1JX1dAtg
vepvAsLqxYgxCsobDaYrw9onoPTnigoXTTJJ1xLyOSMXrEVKiapjRxLUHRT7rL53
CzAY3LA+XTsaj/baY4dMzR5fxmONQ22YNDgSghx1jkQCHd8LV2FS6qR/ClAvoCfM
fUDQoR3/0IQ5m96wVl7CFcqW6HCb/+7vgdaq0OAkvkVCBs6iTFSHscydU2pcYpCj
Ach9xqNBJTJUqGiCB1s84kCJApj39Gv3nClag2qMi5jWdtK+SGAN3TQvpHDLd2pO
LvEq0uGXirZLx1+HhDO/GF0zNZ4pv+ikg/Lzz9owwHMmupv7MQ/v3gBapctqhima
UxfzKHI5XcvNTqQ8CruLAgK5TRiEFytKW31q52pI+Rf4Ut9xtthwpM65zbh24vbL
gbw428wJVce7qTwMP+Eh+HietVj607cUsHLr6VvnUYwY6pydVbgAnCPyp84rMKrq
kTubN0dNiRot7pmVFIU+3F5pyrnmYKqfhmTcSb7RGV4dAQ8zJocZoNawPNGwqpqa
P9HBC179xyff3R6udz+CJCT3rVaFg+pQtCSFu/x+sDL2b4eNZO50cU053n3+TP88
wkmaJRPF9vXt+vTLVVwcqGaal6b1rJKVDU5KGlkuDQ29ct7PR8mI4eQ6O2+F+/vL
6424ketKDvbo7QaHnIf6e+fFc4htk40vCoNdvim9PpvIpkPYlD24Tzgww/5enRbs
LBnnbMzHB5EELngSFF2SCMrMoSW4Ak1IcXthH/vey2jaYwRc7subcPQfz7iNDvoB
SrnPh+4kjmyAc58W9vhPlwqVZ4+F2mCEy4zarKM/6Z1vMzaf4dZ2RoZqm//fNBpl
78kABCIbhFwiYVjHoTlZDkgXEjB3Y6OYl8pE8aIezqICc5nf4tStdOH/Vm9CVNe6
XhNTgiaA/7UipW64JDMrKsxLA13YQtOQRqe/Zsj9w6h9o1aX0qIsryU4/TF1uZ+K
N82Do0FpWh1fiAjxAVUqurH7Lc9YPnQB3aGHp5gkBUhfk0usV7+YnorjdczSV3P3
zZtxq60AjxFragHEULi0LfTO20SA1XbRo6Mrb+D5cSY5Wm9jVteeskqzZAZmvgCS
5OhCzR/B1JPwywhqFTusagh6DlieLjPgv95Wis56Ewu54qc3f/lZlz0jyJfB31Ow
bD2Md8JijGEZpSLQ2gmfyzZ+N5AAFUZ2L5lW7J/BItBEZ1fa9f/RT6KcncoTi966
5GuOZ5KPyO2yPsxvz9WM9VLwRv6BtKlP+03Dnt1CBRpG5qYinaIGBqqwN73vSt5O
9tTSZ1uR13XkIMnDEVG6cDFjPs23pXD++Xmut+aQBXarRu/e3jogIZHqR1a8ImoF
kgP31HdM529kd3LYBlBsog0LATq7AKfTT/Cq4j5BLU1zA7a5hNJxqzSfDdObhzV9
+3eQGRCibebUzEhfQ4SHm9uy7ga00CQP8YqDFXO7PReIDMVyUZdSyXIyRawF6+2z
jT/w/Rxrzg+XiJIuBBmUFCzqI15NxpmIRljbhEfBj2YK1i1LZy0cYdXtucYtnaZM
C/GX76wH/gH4VJHHt0nc1Abs7/JcgzVsOYuO3+OnY2Xe+mjm4YkS4J3KjogbR3Py
zsrc7WbLH8XivUpxwBe50Cugmt5t5nW+eFPyW9ZrKGYQfv7Zy4Xt70FooQinnzXZ
ckngWHoyiXVIkVl83TojAQmPT5I6UkswrS7obqAKWG3yPoSBZGFoSpsx/LbyZqur
kHCSj6ZYptDjwmlKF+03NvzbAbFh3eSAsO7NrILcAXwL0M3nXcRrNxDhGyNfiO/M
MDcTWjuF3BybJiIlDuDXmZcRTOrDGE5oal/2Ar8rmjAJMJa5S+bHwMxce3mEXMzP
A8Mp1tKDOmfjaDlfbdLre/zXxeHfgOE2+EAfDkArQWsmzBS85oxonqLJKi0yDNr1
iF02IMPb1Clq/Mf9uazbgqdmWDlb0Hy5svoLFRstlo31JPcie7zI/k4aniPWc0QW
yUiC0DqB0+5l8OX1WdC365E4KeKtNch0x38r2lOhvYYRyOY6pDvXszQy3lIn1SDx
7Fs/1X+JYSsh7kZlRPkJLgUkOOOREyiDp4lW60eDd3Zv1PtOmdCCj63gFPJmXttF
087/4Iy7Q/gRZ2klqTR7ONhbReiGxMYqTOB4DKK+NGlw/nCL9+UibgBNf0SD2kdY
s5Y3B6jFSxEz8eQB9vb1IzbFWCnvtloQ+FOPj9otTZkmibXvNMuc2xo68HkkrFm9
HRv6XQ9j5Lr3OmImrMTXjofvJvWsoTCVj4sc5fHLzLR0475jgRR5+aqGFyp6xIXs
ANYmsSEhLnUPOIiXEQ6FD+nQ/j6atfxhbHNI0dNdm52yZkGAOBwGkzvHqV7d5T33
TxbfJFBLOS0BbmHZwnYPVKptiQrXa6C3EybGfcjcUfSEvzDCp9Lim6Kf+ocgcr+Y
s6odAixNNiane7ZzwIfbmvbK5BBxRMvM48U77Oy4L6dQxn3xgjultrseSxdj3+57
vh8DlSyGjVIC6w5e2GDR3ouiDP5vaumKpPx7LCe4TLW82HGPY+6VENhQZeArYH68
I9w1PjG61gutpyYMAxkZ+d8kty7Qt2gFkoUjiSYRnoI4b+3pzXrf3CWAc+Fg3POt
E9UDFmEOFpxcTDi9nq8ovXX7+SZdIDjQNoP4ctcXqcDyqgDme6hNj6kzSMoH0VQr
hd4k/i+w7+cwRQV0ekl9OJXJfxbviRNPbTlEJLhUUC3ZkeoeZWaKVVcVNyv7rM7O
USZ1YPf3hplup95G3jjFXD2A3PTUAZ4xU6odJteVO9HlFMnpeaCCnxj6Tl7zV44O
zx2wcxKfnNNyFr6WqIvL0nKO8cBY2JVKCtExeFxTvV2MrJ3Z/AQMviN0zFc8sp1x
txiJhowv9dWdNvXXXUCodS5gPWbZuPwn8Rm7sB3wao8vMayP02bRp5o0mQG31Lrv
L6ur+6XWiIzSQG8oCnHZ4ikXgwn9dsP/l7I01GnwEKT6w+AwuY9bq3e+XSA45dNI
eLgchV4oPFK99EHVQpZwsaXqq2mpak4jScczINRujrlpWFG4S4w0lgz/QdAjSiSc
nN1/E8/rKc49ghuwgaNxhORMOn/g8ozzVClKbFqn/2tL99eByBSRL6QutJ69e6Fh
KyvHL3DMAYWTNP3XZ7jp5FKMP64ZDAmUXDIlsc+DhchSJmPHNxg5HsTLhblzcRev
Vbq5ACQ1Sf7w4aunSFglmfxo7lfeLeXx3kG5cQHSBcdWBtDMaIpJQ63IqsYqBz3F
jYI5VPoopADrtayQgW1vC110AKBuVexOBTls3SPXMrJlWHbIkctdPvVot5MOxliu
AzS5to60j6rfwT78RgkxIUN3dIFhshETvhZUrJgJvPN7vgJVYUD0Enjcl8QjMqte
LguLeEO8za87CbGh1BV1u8fykqfMVZOGjPuUQKK7B1OZHicelGMw6+stJCpiibX8
x9mCtW2ssN01XNR8NwgfGOTFEnMfd/ZTc3b9vSSw38DgaeDaBmTdsXejHdm0X4Za
25mjkWE6oP+S+vTQguX1sMFuzr/A0tUNCFY54MdT/Szh85/FyHOJySIhxn/W/rDN
qalKPC+YMLIj/TuF3FJHK0VoitAie+UbDBe8AZdUUfpTiEYHp/KhsrKn1WqehiaG
SY6RQHdBrCj9KEp6wkZLHIjYNY5w7V9GIysXQnZUiD3zVrHuRMWW1/EyP4jc+ELf
PtbtgejMuga7oCEQqra21B+Yp39oYlLrsuIJ0PLcU8rzQ7weQbntS5v6KtktdL8F
N9rgYj4/ze7liAN4uw3jKLpQQEcAeC2kFWxFJaw5f/NUY1ukWjWDCfXXogZLy9h7
aHjkxWcx2JDWZRAPnahAMLU/P+9d6x/S3f4LD3VvrT/JrHNxd/UMlr9LdP59ojQc
JwgN0qK/KY/ZQ5aENQmZKdRb1U5XDTCg+ImB4bol+pAGZSjQ52SfMBZev9LNTF+i
lUHvUvZhg9DpW9zWSJ7hbfXpW6e+1chCYsXBSuVROF/Mc0mQG5yax2oQdn+F67c9
K0Cbw7QbYgGZiw31TD5zWemkc6RY/J2K8PleDI1E7IWXIHvL8gIX5ilRu9lR1b4F
/MkafPtZFs1hntC+kDX+w/WgQ9eJxx7B49aYvHFeX1rtR/fZMEkoxhXPqYWzmdOb
Pmrx/rhUHF5wdxs9YVi6nxAVQbx2Pew/qb53o9kXraSp859KGDU4qSb10H93XFTL
a0CmyuK9Uh3vK2jOxfBqEce5pZVBQxFVP2BvYhgooRJUz7yO+aerKl3B7FyR2NVk
ta3XSapXonqmAkq2uXpgpMLP/+Ts8H+FAFaYysdwzaxRrItAL5VB58Btz2rSUyhY
q2SUpZTHAOepdSPoUfK17Dap0JNLt6HW8iHNTHpVlYJ/1PFKBkQgjAQAQaez1MnH
cmJ3SEenFUV5DRLs3f2b5YLW3IOqPixLl8zU6lrjOYfr9zGvK79mHSlhH+Gkr8m7
u+tq4WTW1yTex2cB+1ZyppZJ9P0Kechw6UY5iOAz3KYLdhBpRfQJCqfc59WOCgn5
TAYy4Oyp5fZwutn4twFE2468N4aPerLPRkf6ATYOLAvNdn4IghHC+DRSHToDjSXk
AmKTaUS1zq9WpPWLE0gEa98NBz0qXW65ChJsqf2ZgQGe7VKHgPNovfEuJ5pHkxrB
PvwvLyCyQ6pI2m3RVYS+fHT3ab83/BYiPyx/BeYYv8/oGr9JsTK5Wr4+YCs6dgHf
x75lR/+/FML7ch73IfKpAjyceYBy6sp8gTdnPYUknCOn1TMxmiVs6tlNmiS5C/do
mha8etPMiYhikcEfSQ73+H2d/9G6eo5ggxkmYSKD51j1ZNhOJaKBVirKZRfvN8c+
5iJk3VHZVa5JxMzHymtRAznwp4ef5uttsaXuh1B+iagfoUIkQBsBoB13NMlhFF7s
euJZoOqVpXDMHPUK95OY7ghQh3Vt7oswQXWxCSslTXyAZGHwIWlkZITmF9Bg7ui1
YA24ZE94BqybPOz8I2b/gpRvqj1QzaQtFk8Ws5rXlD4gN9ecDt23UP6vFVViWVrl
270MbbYhDB1EDVfWmdTa+FK0h1TTEIQXSTv1c1RahqYRXscCWNAuW1ARwvVCm1uZ
Zdr+d7rIGkUFuMDRn44m+/1Wc9G8WuFU9K/tGhk1spbVD43zIbexv/Viq+O3l3zi
69cDhjOjU/N10q6B3bWoMisaL7dUThCZzESugmGFeTCaCJip+hFjqqYfPgWCJvK7
Wi1lJU9KIZhaiRhd3i3v2s1lqNeO6/0lotAEjl1F4viCi2WeqVyOZrD4rlmjgeBx
rENEzs/9n+VNtKNy5UClHKYnqlQVVoITR9rfgWXrtM2CVB766QIxWyenQsrukJJZ
9LBYM5YCx8voZvRhwaLeY3IdCcCZwHnBtaQicVLQRx29DXfE8+O+wP+6k7n1q5xC
JcNTGB2JBZSJcnQjAXsp4HEcFkkSlJZdn/P+tjgdOJQRl7nEhnuPvwCSMhr4lCy/
CzCxdhzhG410uXIDEcQLX5sgoQi3AAWeNBKJFhzLoa8cWuFhTttGflZTwsYC7+0q
sKk/oo1jXNmVX9x7JW+WIge1+BroobsJcyA9UFKBL4KLT3di6qyuknq6IfZE5Jtc
BZ8Dz4inJ2XFSUd6OahcOx7pD1alRXXTyslGa/ZQVJwoWbA5wEkwdU7m3G2L8Foo
t8c0Z+73oaMg0WxrczPnCYxt/6EmeatpSppCazN7trvea/o252JRzNCm+JBMnhtj
IHZO9XcfufNbJC3ysMnVpn/ccxnAHRfBM2eYA1PPSXugB1OUwAlqFpa+QLRm1xd7
83/CCS25kN0SEKs3AbSsDdQLuGUYH6AmpzrdrtNig6bB8+fRLf1qseHmZMol9wwW
kZqptDAcHKN47NUVX0bKxnz8IQIHXN31tyGwI7p4UJYCtUMQshL1oX2jexX1NTgc
hdbCfKxPs7l8QEF/Rl8a9FHkTtHawNs8ahwKWa5ltNKDModxB2PvfcdmEyqoqwmI
F0eA6Zgciol0VMeLq79YL6IOkrgKwRqutiGLGwE7M1Zl4JGMASFIs1SRJVlJj2yz
XBoi8NsSKx8iuacqGB4DuvD7n8ik+YiOEEQnlT74r/xy0Gl4x0fpTBH0Rk8cMUMg
OLdruI1HX1DHqPtdkTGFacoCfJmPeMrLTrVEuC8P6wXN2jO7hN4oMCc32g94Pjqv
aIQWP+2pbQXE2IlqZ31mf0+O2EWiIu42PloZq+kKJYXePIM8jI3jd5AbGICVtbI9
bpCYxa7XiBUZrgf8Gg1/X/N/xvxRUd9Mtq8ipnie0BsBGdYELHPrRsANx3os8Jpg
KXj5rkM/6dVseruJ7zn64DvhPdVkgtQwuFjJPSGCbmRrZeB8PUKRDNYqrc9njFU1
KfEZNK40R9txTVzFAV+p6swsUXRDBzYsWNa+ro95MH2PXSVURsaoZyAzks/vkSc8
3sLHhIdOIQ67t2HkCfvtWfps2Uw177lliGznJrObzgxbBlg3v9jmS+S96vKBK2L8
eDvc33uk6BJ3gKsOF3qZABWy6NuPcKY6XT6MdNpTzbeJIaiMxYzUoTOYhAsCQUE5
0TK3m99J4s63XKUG3HNhHs8Ex3zcLh9B1II4yxJxIEzBAgYAfn3AmAijmRK9ZoD0
FaqQyLXX0WDavyO1bRCoB+aJdLxPwbRE/JVNwaQc0m+g2gqq/LyUf/Iyvlbi6L0R
oz9aOVhWjRzY/diwljqq1UDyrxuMr/USzq7nTQv4S2vtg+T6e/hhRPxNZPo/3AxX
bKuAttJsJBkkF1TIuXt/S11wycp22WGYmM2Rs8PPtSh2GzHXm4MHNhMBZpYjTNXC
aJ7effHWFFhKToYCNouCPz+6l6sOYgslGNMp87Zgskk6NgDbWXofrgdvpQtjPzgv
25oJed1np4BNNQL/DaGnpT83KoIRPcud7YQEE8x1wREG4DBSEelk69w0AvmiMq3d
XA3LE2TEj/YKNbHV8c56EiuL+nvur8QPs46w6k5/ITUNAiZ0sF2FMWt5sOa08LkQ
lhc2GwPxhuKv9x5B1nN8h0UYVBkRuZ4Z8kBxvryUuhCnt+s+nK8FtiDkq8tgQ2wZ
WkhgIYqcUbfko+kadBHpvnQOnGtDxC1lnA+mrPgm+mBtP9UAf7VHYIw0Wq7XnP3R
0rh3jKY8BfmsJut5I2f8QAFGConTh5TTL8CesQdB5dwOVVCLZixNYb4reB6e+K5Y
lFOov5ZHuc02DKNzcYTBlhQhT4uUDe/wzXQVYNCMu/UvWrhr9M543npA+P5VyVPT
t4HTZIj6nwbbyxWHv9Am4gbesvQt3J+cc6ypaNESqYtI0gBoYXoZHeodlg7PZ0yI
tiC+0j1b2XWOcP6f7pZ+Rruif57EhuSJ3V/jEK6klq6MwJ3E/4jWEaMhAp7kiTPj
4GkXRD2eTn6UCrn5r3LhUHxiEb73sPMAet5IIEHTnQyda9bmT1GObdDeUEVNFpL9
AYM9TkrEdbl1m7acmMiB6axJo5NKCsJ3QoTXWrZM1HHyJ9Wx7OzlbWVEfdxEf6Xp
KlgLufb0UMqxPfXX7/ULmWgg7/iKI6gmNDpGlz8r3On+dlfWUHfyFOfklYOIDLEi
gxKzO8R0gU5YsQxxkqgGQ9kMKeCO+Sa0PcbSBzUHAd8Qv9R2Aomci4giOiprbwoP
PkmPsHEXmg+SGIkUAyE1ps68Tvk1H9zim/eBf55iNRnHbB6Rl+/k0OSa0J23Hpna
bZ4okTVo3iI/OLSv9YplxLVPFcKb4OG0uhfCHP+oxAG9j7nZ734iFEYXyNHcRzWZ
tZ6iu/VaTV7TqKB3fngoWZMvRZA0IIDb4COdULOjvRPkQDMnDIcg5wBYXtLJo7GE
fXRWgudRekE1g73DOgA6oJ3JZ4Iotfn3HqDHFJvDYwK8sH/o7Os5v4Ypwzzfao4q
CLu9YUlmDGXiawyVvMFjruJ7GW0ozjajE2BBqVSTRBiwLOo4jJqVxUhMBzyuiEF9
4GGKygYGxW+yPDWDOxDlwwFZXZYoI//60bfu6VUc7nngYJe5t5Yf4sl+tkQCYnxN
ynmkHorLuTB4Kqew/PoQ4RF+NwBd/cpcHcwUXewz0R2hzX1gkAwWhyXXMKnfhkNF
pQlxL/PlknEozmEYHuDHDvXWzQZ+HO44pvtDWoqtpJDkAMXv+MoTn7fUGbbZlou5
65h2KpgL+7X3iSpbnrrlo/kqMH2VyBCbfHkLpjObs+fIyIYWH0Hir4Zfvl7ZAVrZ
a7bKiu3W9l6hjc5Sc18n/V+Zg/On+4Ct+tSOcJhmvALzNgmRKXvYTcvItvlkD0AA
GrSvQi3yL8zCD6edhtWy5+tk4q37ybk12aJPEDrWcISv/aMxLSJf9hS2OdWIvGbf
8FUSUjopvPeaRS+EDyS7/bAacn8or0j1Bh8nAavA/qXxtFRPJzK8iumNtRoeq+uJ
SympBr1WTBvDQYg+wLrGlrrrd/q2tShSZG8rBX72dYQ438B36SZJcoc6l8gEC1Fw
Lmu3d+qFu0ygsxUk1LZVPiZhVhjtX8F+2kyofUgYDby3otA8S+9YsnwaWVS6TZXS
rtAl0zJBilSCBDFScUj39E7HNBsNSMpC1hX7A5OagTvaaMoCm5fZ2e8/ixpnyu2x
0beEpUyrmGeeWhGsyvW2n6DXFdyCEr+qChTbgMYK7wLEJz66/INplK3QGrjqEvG7
F4ydJgFSF51Bz81ipLB3SswI8gurwITCKMBJZpnwKummpA/n5twMfFAz/oVhIzIz
LcvPB9EPEWYFSzFQo18DH5GVPXoV1+Nau6CyCZG4aYWEt47hM3m5rtF7UVB0u2eQ
cygsWIffxequKjmPCOwBZt9RENkmvAluJ0TcK1ch/KVIuMdn6QAnPoWWLZbjxB7A
INyJgc95sQ/pAhMq4ikycn6R8FaWRKlH4jBSeEpMReeTgGSbhYyHx0w+YaLsTZBn
DaPb5s1ZOosLq3rh1uRB+lY/I3/e05v2PllOAXhQ/mRydi6rHyqOPwQmULxm+pgA
qADOHep4iUrMe7m9s7mjcNkD9ZqAynS6gm5UuQU1BQvLLZP9ZYoL7ESNCSjiaeZV
RoaL9tRFjGcIRAiHMPm33TgVwCeLdgVIn0UCRCo2CEBCWx5LqZhnmn5qpk2eVBPk
LekzKpCVUxTeIjVSI0bnePDdKvuWQPpMRjBD1Iky/qMPSpN7RI/hS7Q7hWxwqSHO
72abKctHcHT4nF5wPhwwYF/IVPJD91HnN+g5zWofs8vQhQTzebJ4p4CJs+tTEbMH
lVixLr7Us0NobH0bVZThGUdwyBd1iXa3osHugPpweJOg1Ahd0A59UXV5+DtSY/Ks
1lrY5wKEi3loU35zYsjUqBJ5MWRV5xvK6Bxk4kvJZXzuo0th7aUM3vyN0Vgw+f1l
0uTPE2DP4xLFVQYhHRbq/ixxXyGo5GzDl9PA3WENweFIETIiPjoxUT1q+9QlhDpv
fNYeSI4Ht2kGJouuG73poCaR5//U4Lab8/eCnDpuHenrJyVz1XygwgCmjooYvxLy
zAlfQkxs2vKaGigM6RgoBGThQhZByRBkv1JWtXXt0iq+mOjHDx/teibNY4vGyZJ0
tTCLIVSC5JaJyiHWm7SIIMXU3pHIo7ODHs3UkU/K8G3epLPQZ9/LAYKl3kO4GQz9
0iUK6P9pWaME+bqg1aDmJR16JkEGlX/j1zJVzEmONifAAOibWRLIBtMFCTcDkomB
6fLyxIIjN+ehAcMF/YHxYD5jpFuPGI3fPKiHvCGjffoeeo9ahGWLjDMQcRcvIVxF
FAyDOPdBKk2sSKMk4A1gC5ulc3cM+itdgCeT8ISKYOvMEeYskCd/rT6UddImhIux
udD89LU6BBYnJRNUlB/eZ/hY6cJuMd48sk4JjG1HDc4/5r2a1j2fi29gJE0a5WhF
lPQwJfdE1RdsC4AvgqsOUj0FFZsHW5sQ+fj4J4O5p6sUEwSiqiv7xMYglB1Ehf1X
UxA8cOwK5d3ZBTlykxNak43t+fQxX2/4D4f6fNbnk9oqvtAc6a1g55/2x3X2Qpmu
KhADOUFr5mgy9dOkXZ7Kbpyu2LyjjWJwii9lf6XQk2xjFFz/67YXpTvF9sP3okyB
m0i+n4530Z8FZ4vPbUFXP/MuyhjCxlbSyfS00PGbb4lhh0ubRdmFKIggiiUwxONB
73UDAtGq4zQ9aY/BaG5cAGvWxl7H+YbHcT5L19lGVIls4fdCoFTB5pG0rIWUb7bB
ZQk+m2fPfGI9PB9leLwvYy0XxR6YgHlrgDwKP7M7haVEjl0M1P2opJroXaMNsJCI
gv0fj6BEcECxnkf6qtmDhrWD5Rx+rtg8zziy0Xoh2Aye4ttHqhFHyJ7CeJZge0Bs
b+NIenyBYXQl+855Q/7pxeHkL6UtcuUCOU3mSDDBdGxQxBlW+08Q/jfH0zgkbpwy
W6IYR38YUQwDZyDHE+3okacF3iQ2KhAHb3o7IfSD1GzJkNMByduRPKFaTQPUWnsB
UfUqPyeOW+cVHdnLOterBe2GyKwgU6Hpr6/p/Oa75OWFFpr3rIAkENL1k8VjE3C9
VATj5OqG05XWAdm6CmN9UqK92+62siBSGokPXN7pVU0m2gXIzhaLJuiqoFg0QnKX
J6FR9XbhqAf1hrqcR+x+gieNjfT2wSD73VX/6jDP6NfQehvfnYJgWFn792W/9bMe
+YoQ4oIDYoR03goJD9QgH0nRx7Re7ns+5ZdBWnFyTBE5pm6Qz2sb+8qtDvSsotH8
gkgEtYfw8+WixUVnyrEWUACOzQl78YA09r3Y4XvBtz+TG7oq61LhOpaUa1F1Mkse
vKOvN0aD9VNv+Ilrkn06NDPTUcrUWycil66fCSYXRXwe5PHDF+ScAckVdz73ZoNp
tguFmvZB4RZ9UQD7G495afScIUOBEeBEHFtNdPL3q1gwJg1eh4S90r2i8a81BaOs
YzK9SYaqe+W+yprkXPmjou/WzYB3LrP2VmTj9WO/le9rYpU+Ov+jckPYMC4+rN1Y
Jp4VzQwGqBUdgKFr/Gyh37LzhUbeKm0o9HO+KQo6gc8VgsP6L5CimFIYMiku9umH
nTvJhNlJHw8PFlXan1W0mZseNknkEIAFmWTGoVLvxj2rqs1GuyWkvLK+6W2Tbgm9
xDRRiNB46nWpxVp2sIBLWI7dhdnx685fJF+tpDdsVJoF4NNrFCUhapcM5Hwfi4Db
serJtaev3opvRV3Kuzle2axmXbYyhjawg1QqsdgIUd5iE7W2zUVe65osWOtdz8lT
SX/dPIvfbRfnjr0ObnKyTkUHdUsO+OwnW1+PIinqpGKtqVYVsDsRulLifa/jPg9V
xi7rzNQy6m42K4/hSA0V+B4dzXrXe0w99WTJA+jNQo4nQT79nzSCgkB5U2Axd7b2
XGJ6BbQoToswttZM5hL/prFqyOHPadVuffMW9lPeJNqZzVzHnGsR3nu6sqOjGvrj
LCMGnXeEXYV391OtRZgP8okLW7ucIakfnrpDH0FfOHl8GQ2ByeyUXpbCRx9UqZot
cIyVC8sbLw1Du2D/n4/G/YqDXwuk0C6GOZE/jMwsR3xN0piO9hBMsfcMbyEjDjwq
W53iHEmBsiimnUi1msOf8ytYfUi6d3t+lGgSTFlCE/dPtMIYxRy67b0tNYmNSeGY
Iwvyx8oim1CIEds0UhCOiinnwNNSPTvuevZWosmczkl9Oid0mtaW4T3ktR2RbJMK
YZK3YABRmlMVE0knl+vz7uWsolAGuKySpMfwzSdH4el41Bfs4ROIKEzmMAdsqxmn
ax6aW0aj5xcfdg35ONEsodh/8JyORmLBv1cZFmhKmqT/LXny5gW5dAkwoS2OCSNl
N+DAuMUopwU3vgvNQ6S576JLny43qdtOejMDkp0n/h1FIx4lDmdA94RB0hddAoqn
bn+l+S8G0oy45/nGs5Y4CGjizjKbyGhLYH54wyprD4eRdaNQdE3iFqLFF9sLMUo/
K3ZRs0GIYf17lokC7nMktjL1/jagpo6f3ABase+FE0vDKt8wG7nqt+Phkhwbf8es
kquio4d5BIKHhwQ3v+DzFEJuDkGSiaYlO1/qmBjhCUCLugZn+hT+5MyOxUvAPg16
o6C9ZT6gv5Z5eBCtL6OmJS5tKig9WxGEoDs+UN6poUHWbQPMRxEPdYgfTU2xqGTB
HO/DJYLjtnUT6VEn5D+VBerz7tPoIVDMmJXgsidvJ0vtMLHbc4ulFTOiBsIbuene
5NhIjcX4E6sWFDmLEeMnZ7UodMQNaqorIgDohTyTxRjUJzq+cOCXcLuYXgAPDyDP
lYNF8XVh0WTdvUgwq0FmEyLnS+IggYsSYM9aPAeMm9Pl5yJWJQUdAJST8mfT9e3z
cyZGkkoMOM0z1RCk+BhXvwJHpkL2xRzpr7y0FKGoTwdm9yIeMN/3z+nyVwNbTyzP
f5gN7YPbfrx7Tq/Qk1j42SvHFIFzcHmbGp0t28Ktjnv7NkbzNblFXJu9gwOxcORn
0ecOy2x8snFGmU00nRiuWjU/nDhjZolvF4CTzORclHbEoAG8hCE9ottn2Y3VQlBu
8pl/gyNPpXOI4lUTL6UZmSBwOO6tlV9MrCtyPcwMErL3A+mRnV6lETImyCMimGZ8
B7v2nsHZoaGxdrD1LZF9zisktkubRVYVrxi+E61SkVRNuLJ/nG76vZQFS+ET4iBf
/ZAXfiXTG/0LG4KsE+0b8u4YPSRPNHk7Khu3CXxaYAbKojke34G/LtDrl28X3a6R
6up8sQLiAZfsfjFuVGEnNRzkJ6lNpvLGnHnVAPXh3y6NgIGg0Ag2yKrP6Sp+AG22
Ug3UMzYF7px0ZlUWTeuwqf5PQZaWQzkIGccyC4ai9amAUHvmRrN93rMan2wt1ViL
kaUfrtkoR7gd/9/tFNmczOUSlXFu6ZE/kiBgfL28Z0UNvpEaJVh75dzIeUQeTQmb
GR33w5zgTmBm3NF9ZDsD4937dt36y47dAmdJ36B1yeEPGeZGAH5cjsROeQ4w+a6Z
a+O54mIQ9qg+ENP2ri26Q/Y2ygeUcmUMg70/B8+3m5f1XVh4bLlEzOmRe2DqXtXg
0QkhVnx8q+/drQ1NaP7Zbv/viLIoWP3wv66Dn+QlbVN0jUTF04dSenWtQcuBTXYn
+w8GihSa9Bu4K8v/4Yb5wCAYIPn8lQSdFxO1M3VRPssbUgomq9QR/L2owB2+W9qb
yXavzX8hHJEAcInuNT0ENNYEPwaX8ZqJeiQoIXUzxO0cAarLSyvQ5mRJwy2ZIxDP
OARNphimtepqch1aXpT5dC86RHyIc0a3+1rOKe0sQUNnZB5qGd5gB0qVcuqirK/7
98nT7SiR3zIZ1PVVd6r7hKlvbL6WqdCrjtY45G1QCCgJWwHVPp+W90G/LsiRaWmB
JG7E06aUz96nypF07PHtPP/0mqPaCXjfe+g4H8QPgytoGmL3BBh5+rWd/l5aj/81
zmY0djeM043T1ToH4iQn/SPWeIhMCkS9NzqeKIXjXFnejJ55tlDKZLvcWQuo9nWS
eLp0il0hOEHPyK+zSc/2TYdrP2A4hytM2krZuObksACTai3BgZR3bQ/IuceYeaI6
pjcCs+kenlGtYd3AZetlw9SmjhdrZ6fFN656NvmZxAU6Mzdvq2MRRXiE0TVFBUmT
+VE+I2MngoU0tXvL0DmAaH9l2wF1sbv88yBwRoW4KUthC1iMakPNLHrlx3zvhBul
9Q47FaNpuK0m7G+QRlO+JX2HZZUkQnhnC/Xo1VSK8uttrnnxeKyGh1MWTSnCpAbe
C+PYA8l4jotPKv+tY+cjiMJjVIpqyvYmGDgWGmsriGFMPuzycWRX86ukE4IQJCrg
/ujOlUtWwsMIWhEdICqzEO5AnujQ5OhqXqTE7rHqi2V1+pgfTMrha8Pv7YYKHr5u
DK9C0U6PmH/8iQ6btFq93i8/Hbz3UXhwT5dGBoOqkjNiQNyLOv7szlC5n8E+xBbJ
5Wwue5SgIxFMqw3vd2i700aAnfjyE1+CsYllEVoCsdLlVbvwoMz1WKn7syxQPqG+
WhlAnFbDi8xWUef7TiWlPdhWEDgESsbgOwUA8wLmY0Un7lY8opUJE5tJa7UU5Qso
6+wO1NXNFT9rahk6SUFsSNWJn07VzlPaeXv8Ifbdnca4N6S6AKDXIMartNqq/qcc
enl/GkVNJzhrgP5hrWGB7EHyTV+jZUsm/MN/dh5DUrUqZ0XyotqvUmwEmaOEcDSL
+vMxUDnkcnrWQetq2LYqeRYftFnZ6fVi6qYEx6az6A+qfL4zYYjsUSsRPxOoC2WH
e78x/Wd2d3iGnkYpLHFAkiMGeulKkq17HPXCtovrdfBfxk/TvPe4/HleJ8qNKhYC
tjUAjJqew89/X6KCW71IiBPaLC9ll6+efxI56EghD01AfQKYRiy1XcV4w6hJ+O7u
Cex5dXIRHNW30f2cmsOtGkR7DQdtCGbSsROY4uASc+l1n8Kd57g7dnntuuP4Mx1t
Enq00zG10nP10Fcy0fXtCcd93yOnvAZdEyZaoqkcXayJtWi1TTFLgGDbnI8Pj0b8
ILivNes2B73uoIXm8S+kKWMCqeoWmu46G+gjfcYnSCUnuqNoNy69C6qw33LyivbC
sXPTPqk+owmGkhdUEgNfLKjxbUW/E9tLdFKyevTNMRtNui4Lw2ybaPXWF95fTfwa
LZA6BRVoG7w+Eda0QYUlRdLSJFtXgoMUjm6rtdSxIUVD75OvJylzmHP34xtKoQ6t
jAgV47X/lx010pnuZmR8yUXvd1vtL7Uf3S7mFAGGaymlFQTKa7ivlb3RNiolmWd1
5MCacq/sC15x7M331vy4Py2i0kMqQCylEMfd6hlyDt8GIV9mVmk3H+nMyxNyAanr
LKKLTNkszA0gfFr+Gpt7qnmbWydAViCVs32DQICLD6j+UnY6LsVjc64n5vG92yrR
0gQ0ShKtD39HxbdmWZcqcPp++S07CFqbOwdPXX7VFaxfZzChCa/2/Tcjp5NLAUwo
hQAM25N/7895ik2L6Wi1OKwmLxd0ytuRmQKsiJz/o0HfLH04fw7SyK3/4LuN8+sU
N/3ACeVjOH2/4iWG+hw47GU5eH2lG0vy1M+PyKElpPTUjlt6wd6gE+vQrycJdKdG
Xo2blCkDLK9nnOWSnLkLUj4zPSf+ychViV1Yv+tv3i1/AY4k0c57uitjNCZE/A2M
LkPcjOQld6d5GxSgmaB/B/lAaHs6m+JpRwrap/po/AGZWTwcxVG7l8JDU4f7fHJy
y24z5J8jgQB5O94T+WeqWN/E0c1AtBqo8jDh+HQ6uD60h8gQyL+b1ej7E3BReCw3
8kNsmM2jbAT4f4BB+pGkiSG0y9wE9jffJ2PzKvyQJVecEHW5koiP58FbX1PL3Dq9
cSfNBo0j5+CgcLZfUS2uKw3Ki+4TeqWCt79ddbpl65HGTwlYculqwexQNWnCxRdv
t8+ZXAe3u0tLqQWX44b21UDU+lbysk0aj3/S1RHtlrBiTewcc9UWxbaFMzeNoB5G
rN2rvxc+YFbv21Wr4NiFWqlphy9hWN1fiTd3zFM89EV1/rTp10RO0VCnMhOlTqK4
y6a6yLrTVASgRuQSa6+jDZZ+5deFnYOJaF2Fy1PZ9Bb6JbNoLFXMvj0E/KYCFaXL
ARXFZgNPKhd9a40xkFUffSmwFf+WW1ZCrMbmCoLW5k765sBeGhfT5d95rdnMvm2Z
gKquPW2eQck/7vlo/dX3uTax/b193RVZET3ISIHwgpDZIforK8T2kBKDoEhh9LKM
JAtljts3VGVrKnttecamxHntgS1Vf2WvHQcegb00MLsvQZdK9ktvV5ys1M53HdWh
kFWJnm4foVpPWYClZFwzDGY06lrc0aouiv+cDcYnsGyOYNpwia6C73c4YkVIKoK4
eMC+85bfLiOA252fkr6MUZ/53XrWsY+5o4cdxV7yg8wqySv81NSbYMVCzhxBKO0u
32V6ZymA3emBhRrzSsS5UXYwVDb+QFV8TDtGH84UkpWTVsV65WzcqYcPX9JeSui7
beY5FuZiGjMYLJnM6AIJTe0Us7eMRCWJ8gtVe0CI03R1W249exrJQ+YBDFLt9gT2
yL6pb2zX/+HV5Oi0qrDyTui5U8eoRhE2ZQBYc5NwXdDLBqTTkqRYI4O830D3eFZa
3Q2+hNqkcP7XlC6kz3fs7JJe5L6FhLKmhM1DwMH3vCqYGh2Xq2UwW2G0Qtgorwlj
c2X866o4sf7kAJh7PFcy2VN1kZIT0a/UzjbT9JsPWS13xhor/rqJuAai3xoDOwfk
pnSTDCDFQBjHvoxa5OslwRcIbU8xdKlw2sypTnPcbJnb8CQ5o2S+AxVQJBfcrmKm
gkDt2jOLnB+aNAw5t/aIShucYUdH0oYLC9sRuV3dDbbHRCnhVT86TICcA5lxQtHk
QVUN2cQMEm3+lDQQ5KJhZJcKGXsjFEVYlh7JYLpG6+gFdKPZ1AB44JnNrTo3a4q6
Mnjpalr9iuynJ1B+vGUWML7sOX16xgAeh+/5Exfcq0SOuYXCaDKbL+owWU4D3nj0
lctKqd9WitTBGbfp9EKI6+fqoQmoZn8lhC5fYsgG/LPjIiPrguwblvP7YpsICXA6
FA+vvZx/0a2KT1VGFnoUzf52+DCCgyy4OVuF0s5C9FhXPeu8S5+v2ABkd8+//a7l
3VHTZtQEpe4x2ODEAvavpkhYDUnNySaLEB4TmGAky1CEdxWy/C4JCIE2TXPpQuQ3
Tv6KDrygDF9Z+Czb2Dw4aHGf55+CtduPH6U/HgS4h1xD0nb3VJhNr8M6nEa1O0T7
qAXr6iNB34Z27VXt1dTY5LgVoHkEDMsxS2f2wdNAmKbrnAemXiEVA6ZuOIhfNcZI
eSdPKTeS9edQN8kMzn33iAcSsTSA4muc2tbL7zlXB7vWJ4HBab+7JproCp6C30Oy
dRpU0wpopXq/H4siJIGbYKYFwxguzHPsxBYqWB4eAcn0tkFzGJFWuJkPLwIqPBm/
ZdIXrlEVvSbofOEr4skgeFHt1VYjMzsFKt26xifdiiWWeNZJXsbQMBh25+m4pOcn
KiwbU2B7eUrIHbxt8ISDQ+DKnYCVjYJpvgwvHBItKkKpTfpjj/pQwTKaqAR7GeKM
Ds2XGhjtb+fnCh28ct6bNwLQnJO1F9RtUam7Ii9I705hP57xIyfrFrlt8Hb5No3z
gF7na5De5QnH9dn5Rewqwn5qjWW6gi/jyB61FTa+QR9rWMkXM+B/ASb1TwfPQoF3
Bw7xP4pKzfBP7cv+EqT/GqJtg36G9fGP9Dt8jNFOqKoD+Z+F/qQ+/egkF+pHeNvm
cQPLiuDrw/3nOOtTxHFw4TbBg7QqYG3B7FJkTZeJa7ZMZYF8KlYufNEAeGBxXR2A
iA2TukTRD3CzLOiYxDhz7l8Cew/J2LMQXwQAoZfSRc/wzPzxlssMAo3gO1m379RL
ALGOW3SZOmquAabyh3/ALvTwZ6Mo5PIkVEhLnxYX0ByUWwEomC9c6LpT6/76HGsK
cb/yRwP98ccnbe8MoYz5tAUq6FVLOuu0Hm4kOvYpBcfeKZ5SpxNMvBcHH6qR9CFA
uJh/tVThM5kCl0bcBHuMskDBwto5u36tBSFj8/r15JnnofZqfRKWkQYME23HzKtt
d3BRD1K23Jiu5xPVgocnqmVz9ueWHqFHQWp5Fbrk4st3lWdlL5cyZa7ezTUmT+76
NpgttbOS2JBg9GqBRmO7iF36bCN2VsCeDeuZXx3/1MB3zS8jmXYCzsDzK6jRGmMu
9maWSdjW/0NTotuoaZYLo1Vg4k+LorTjXPH58kCoeo6/Lo6FB5BoxLzEzAkSDnD7
0dRjRG71H0a13Qum41VGOfLm6i46UzxJnQvpziLub29aEzTl2Bre8Y8NyAsDYE6p
Ib23WxrQE1Tpui8zENSyajaMG69MENvEipTV6CccQ0iaLBHfM4ouymUOqTY+Iz8I
XYmWLB+6aPmtkEAMgMRYLoLUENadq8MILUQHwThU0jY+f5NLRTaxVAtFHaN2uIUP
zFnWQvnL8fTQu3EbbTRehb70MRAJFD0l5DQX2GhQXymEiCa1Aq375D0R1zxhQrdE
bPcFuBQVLXZfTdYsRYeWKGNM54gxN+Sy0uV6udDnZrLW/f0ttkVU+oQ+yzfu869c
24V432F2+9T65gXR8r7trJeZgddb3GpEREymgHNHpQCT6SQL8CaVi0BrQUrSKsTM
A3vUl7B5VAZRuY8FQAVtfdZt1tNFDdpNVYW7Cy+A7+ejpT4b7IR0uoLP3Az0eJAN
eU1S8g8Gzft2cn+BuIsX97u0eCea8FdrI+JQJpomcucJjvK+/aAKMZLvnM8CE8vI
M1oVjRXn/uK76Vo4lA76pfEGc/aVoyQr73F45/Z3jUj0FAdF2EGb2NS67tA+YHcR
ipBrZGXwtnEuBg55Z03Q1uY3fiNpjmgTruhuhOC1GCYL38OSj+E9BFsGNy9GXuMW
AC1rL5lqhR8nK1N3xHE+X4B9nR4Xeskv1gCQplrvivfGpLWkg6T6ZCWsd4+gDNJq
EZW6DxLGcYJ2LWK7Dpwovz0PGw584qHwOH+W1Kte0dP53ebF2UbFmfrsRwRPwYI7
Wfw8u6Ue5WP62aovEaBNBmzpu5JwfxJtBPo6FQrH9q0Hr14aITb4zmliluexHS2o
g1As4fjCd2y26CNBgHJx9ZV+ACCMCchr9AD3lRtfcUKTwitteEmd61IXYsmIU2XD
cbIV7FT4ByvP0gRtzB5KdcGKwMJxUi7kzPE6yuvEcazEktGsSRyvkZTw8nX63LNI
v7f6a6mNWXCWOC+eTZhRW/3e/m5ceDpUtyF7XcQxJ+K/S6YWpy3IBa5y08m/tFUW
KftrXpRJ274XwdI6pRB3O/btUBD/+aBI4o7zxfMQVkKzqFuZiD6c3ix1GlSZ6HI0
gJOcsEWyvciyyJ+nbOzS1tetCgZZWK1pNQZPSqlKsDn/rdKMteHmjaVccQt3DhJN
Gw+WBSarA50nvrCaYgdePBXJikfgKIsvyhuHNLQ90AtNc/akIcL4+c8PiRO8HuMG
oQGCrLPLe5qIjArFp7AugLGC7OpTNvvush5B2tBI4ef0abqdh60xC4J8EJCphAg2
YsieekMLv89RSkt+WDitigkNebx4Mrl/PMw7qXzOD/6QpHFJbGrGHrSmnoLD3avs
7INGIQvXfeq66lxHUgc1By7aYpRoGA7ZXRVI0d+EOR75hhNLpXbCNaGtt7RnucZE
Xnzc93sTIsZ4q5rWywuaF5io4PEG3ufAV3/KmoBUrIk0g2dZdxx0MWj4GZPgb0Wf
Acf0+GJByPDMHBlh2lHKMNHk601yuPXgDm5Z2Oo799Vv1b4qQViImzZm2O/fgYHC
BADMu1WKzItZWFUABWcnl3HwVy7BMKEIFfAe5IXb9UhlZZaVbhbzCS5YUK4xlcO4
ke7WOMId3GwjscgoQg6zYa3+WXvCOGjpYP0lwS3G2HhoxKl4QFoGVDY/W53nl8c/
zezgL3o3ZwC0ft1LGKwnxMgL2TlK1u/b4UmLL1KE1lLywc0RIlNyr79G1kLHPEaG
pnkK9vWH7PZTaWs36aalYhqKhiGHIxfaKxbiZoU2qAbJWVv9RkVwqWDIHeZtmHZa
K+6y3rppzNezduE2SogyGRyczIA7PObJlwKsrBtUGp4z0fwBoyle43hOqABWxU9x
Hp239rJumY8nQmPeFDDUeGwFtum3NxJOroftvrZaUTPooZ78HWzXoBT0aJMLy9Av
edhZtKLhZGqdVAK+PRLAThC1C8kkjqy9dr/1ZamNM7w4jZeu4A3OKcHwuFd0oVa3
cpZUWg1rI8FfrZEpKzr587qRa3fP6x+JfiwYZHVev39TAdC79VoCLJN6U5eS4pLl
SKY8oRmDgWN+DJ6wbv6Ow9u95xz/9v1qC2rvmZ81WInQDHr5LIANyIqk5gTFofeU
Ohw79JQOsRzHLJ5fM+cEz0IOC4pvmxqEv7d0aY3crmvfQ0Anyk8GTGwyH6PSjKmQ
7BtYHn2nBJA3aV2x1r2sx/fRu57omnPHsZxGYtBznGARNE60b2DWxY4tz73MBtIP
faehewvmWo96Mwhbvl6TLOjyI5J86sr5RzULpzIhzXB0xRs5P0lDoRNfie6hWsfE
uPJZR+v2uVJQ12hs7uaBJZON6KyVSlla9jzGnj4yV6wgXLMvxlmw2vgnxsxYXOvh
Hvv5/O8F7mHULxcNVGiGYnqEagTlRBVHV2yXL8icDpWW3Wnsk8DSJSlY27ilNa3Z
YBqkbD76N9gJoUbS5qErExKZp9fDdSn/MJOeTUG1noMTxXw5BBWFrGBUMZ4Fm1N3
i7qIFvQ47adogMXeltRjsLdi4NiaSO4uttBJ7ll8A5phF4uI3BQQJEI090dXtTeo
ty8w8L0drgYpAJISbHDbGej9VaIA+ssldKSpbxU2+y2vBdSU5INN+4ee8HnLhpTN
Xb4UI2u8ody6PK8vx68SPFxZYEEeJlxCH0EfKaQkVOhAamKB7W9ZFn5B87bVr4S3
cbsjUWupWYOJi8nTW0o91UhlTfc335P5IwpoN+jBIjAkYW2/SwiXvnQkBs3H+Jat
7/7p1m865tlYV3WIDoHw1mFLJxfAF8y+Deyi8AuIhF0VWvTqkSaFxC5PcmTilU7I
Oe/Bv8YhjxrYnGqAZr9jjlBU/O+wxrLm+oglx5NvzxwgglqZTq2ub7kyPjdkQoHp
GMm0qCrONdpFUv9P0MZ51tZn896+IGTDWyLyT285m3JzcyByCRwPRhwwvLEnSIUY
n4u0DNta3+EI/qOYMBJTKB+Zbo9pr9ZrSRzSKVtJ5ZDSeApaZrwwJ/y4GVwtrENs
Emc0RT876LqXfE9HtvfAwN/S6KCtzH0KNUtqMkww4JLtud89jADTw7Dzx0JMaNg0
+c/Y8j5NYH9a07VwPiURUf+UhepLsrTM1cFCPNujLt9s7sKZzhxENe2c7X9ir+9v
arzyFF+bLUql/XFnOCBFSeh3wmzWoGxEm1c9vm3R2DfyKh4e5vQ4Ap+95mbdJ8ZL
DpXG4hTniDBeZYIBcAYexp+pRZvFFbhYwflOsBdvDd8s0MYOQ3tuiwx3WE3NZEfG
fFsDQHDz2k++DhfO6kf5yewW1zycT6Bw55EbgZ8qv1FfWv8wjiB0pb2wBerUdCRx
5UctB2xEx9Spzi1uxf4/MGHBBtFyRKcoO32bWQ1fX8Za8uA2DJhdEQCInKOnRcYp
3WfBA6srHGtva3VcUOG3KemkxkD1ZNR8Fu8XIMv4plJ3Arl4R5GFLgOTMCfHLnd6
HELlokobhekiNXCHVFm0QM3YwJAiAzF2C3ILblVEJWcrERlHso1DAbtcvftbejw9
xBqmqj50hCjMyWEwDsHsbZBombwZliI9XFygm406474JIq4buuDViY/Y87+PO2Yy
anxpKa+S3BN+Km6u/w7hDds33Pna9kXyUcpH+VmFmEo1/YiMMCJTnvDfDMG+YVbd
wXxIflM9DpQ6dGe10C19taxj1k1ez19W54fYyV4hyJFyDb2MWGg6UzuSg4ySCZC0
Cc7UyW+WjFvwMddFV0wfkaoOESfY57ye6Yv1IEMognwWAa8ZW3RkR6i7XHDdVOzP
H73JJKHCZR8bIkygtcmDSncvBjrSnZu/rf7TTK4gLLNkqOpbTpegMMA/uxnoCQ0F
k9X5pX544PtMR0NsNncsoSx7oU0WpMzL5xYxV7PwMRyn0U2EDjV1NhTfJryd1932
1itK5tKniHKV91Z3240uM8Cp3IEFDTWMybMYRSzroI1odJNyw55HWJxHOAjHZ2OH
HBYvRja9289HZt3r08fyO9IUZQ5b0g+X8tsiPuKf2flClVJVYN+tat7B0DKcyUOi
mH6qZkvj9h7vgNKl5SMfKUIMfwjpzadM8mfHZAs2lTLkjISrw1oURBwIbfg6y1AU
DNF4IFSapnD9daCflZ9BskC2eCqx4E43t7/w2VxFYlTULiU8EM1TSb8jYSKzp73H
wl4znXrE7/eY7jsXwzRQ4HqDDgaw9U+y72KMpgKkEeZeZaZA15GGVImlmsRH7jSD
qWUhF0c9yl8ZiXgOb0bRrhqG6xI+9Groa4UsMGvhZmyzDiB7S6WgBBxUwpfKLl9b
PYAGlN62gBgE9f1tpTiI7Nvc4SoHvRZaj0VSplYffN2W3f9M9XruYTvidhp8ttyB
CB6w+sfH6aIMbaNi9Gfy6duQewgBRSvwXY3eg9yZiLtQYYls5eSWNXUTgWIHNHTm
yQlNaosnrlCdBMjXnwOxzn9mZIE12/19AoF96SYRZtLOOyMTaUKqvoEQvvZ9+k0K
PEw3nu7lK3gKrdH5ScPljA/07JoPx4+AV1WluehTU5KQ7ticKPsIbwBzGIz7zoEq
0sITecYvO8UuQYDiqHcJKxQRUV+u7wpDrIdXzUzQTpyh0WGbdKy3wO6ioENsto1U
xSubQk4X7ZC/sXTArx21IT9eS1s0NwOS6ubR4vE3gWcanY0VUkZSY0ObLkYK/aYx
dRxizXFjmbWNRP2eP2fmE8pMesJ+/u22Saxb0NkYNXGHmZSqYNVixiHsasJcxaW5
JfkRVKgZssF94Et2Fgn/1jWj5yT6Gv8ju6W0bHRYxRJXeKiqB8lBvcvKLRf31MB5
yrJKwMjEDZVEz8qIaCaN6LDELUaJj5sAgHRYkKz8qmjUjNOGEcpRYilglC+eVXBD
L5RtMV7EfGLEAZgESNI7FARY3iwRvsWMOARHFRpHzMVIR3Y5tnOvIBiRutiqmzql
Iaf9w5d/Wu8iY26wLB9yEGDBbkzXLC1IZeQfVtFQRwa7Z6Ym2xbiFcjoZCYLjUgZ
NHztjihkJCGyo6ityAUY6ken+8Hhpf8R7PPpeAw4fkubwnZNYU06XSM/6vKxayBa
23TXlwPe+xIhDH239U7qqej2g/waVdm18jT8JOhPBGTeJMz5ErCLQ+5z+uxCvXsz
KTR6jCTQg0O9gutmJ8opwizJqCZsdwnJE6fWaVU29OiNddvADJ7P5ZzBz54PHIFs
oFDO7rO/rQ+GDHhw/b+8dLbo3UxDCOqIYWNk5OrXqfHUTlbvi6eTpsvr2SXfrgCo
o3miJbc5RBDW0Vx7PN7ZyfaKlGfsDiXZsXUFF4NqvNfKBIvSBKQt/bVTH+5nw2CO
rsQGuTYl3SHneK7Ll+11WKv18NaOeDPA08/kgLc20EScDuhahmU6pwuaNlzcvPay
SpPuiThgFPB5fXengJe2zhMGenmaFeA5v9MKNO3kdNPdqmMG3u+gI2SYySZReP9M
P4/dtR4X+AWaUbCQwcQw9R1mw4+EAGzbXtpn+iRNPTGgq8dph+vhs5IZJEI01kDR
EhDi9a5sRkeSkrSy5SU6MlwFa6ZoX0rKf4539j2wlx4hejwiO6GF0F/hqTY/RrYT
eRu5iiAOln4hE4k3q2kFYonBla9nZaCdX5yTlUS3U+ZL4jTtMTbW41sAYBlXOaXf
SxqIGFqVvrtzDNlqGWaz0YUzwy69dc63WxFgPycDP6AQ3qwA91ck3mIvtW20whZx
ONpdfOtXQDvw0VGduJDSSElRS72XVgaf3/m+LAyO1UbNfcipV0S1TxrQY/onQXHu
CefQM2rWY6aDojSeU9RYNdgfR1AtjzfhaVAcDv1wN6YgHGCqyya1qHf86LMpwNYc
Yi+SBnvsGr4hYsZ3p/MoQNOCsLY17KtjXvHOUY/BsU2pQm8ge8FLyTijKxY0ISmh
2Xt3rT3WNiZ0F7R6xQirVD8s+QS+w1EoIIvk5RZZTiZCppgeGVIaAFnUr2qWng5K
nkxfLPUV9q0rSCMNs3OIxYllK+MKDTlBCtelZlI2cITSy+m1zs4sxUuYPzln9BNm
lIr5j1gJTi3Msm79TrQvBRw3cYSpiBbFYf0za+c/uiWPOVmjeIxsFQEb1cE78dBG
tsXaHGQBJ9q2n5aMRjxo+qBrhCTPoph5mEax1w+/dLVNk5P9/7fQe/ccqHgR62PC
x7qeK8Wf9IZJ/KRkYROni3mIwdZKwDpbLwGx4NALTKQ19cW65uaLcoevUx8UeaMR
UPmNWrt8jtJxd5vZ46/rhRw1dfYPy9iunoA4q4XzStvY5PApXbVqu+noRG68cOP/
ify29O64DYfs4nd/ETVuZQPdndVqtU6YVGnXF3kVUKs7uXzrEpxEhrNyTTT7R7oz
Rlg5PDRNKWUNQYiTBcZvO8NKh9dQGs3CVFcU/v+KsIUnErnI/qfkJeNBmHaiDldL
Q3If+NYn7gAtRyl4wi7HX1bytRHFfwC7fa685coJxy36faJxcj4OwJWi7jjmP3JB
DqA/zVlx7WCe/vKqnRcZmBvV9TZNGZu6OTkYjoIClp5gek4mids/XnnAe6Tg9TqS
Y+qQgh9pM2bZmcOFYFnx2uWiG1sJ8g6KoGdKJ6/CqOyud3pTSF9Zs+6Hx0XKbkHu
NEf9rS7CKUaNMxu8YexSTUqztYnlkrOHGWEY3oyR5+eHVOUt74ByjR8//v1YFeMk
JsjUyfVAqUUc+zQ+7DoOQQnoUo2eFpaqE84yFch1yc0VBqnXgrmY+R1LoVrQ1bhT
OCz+QJZ44rulL27j6IkhL3AA+1HLsBto37pWrCqyDz+aDXu42Lx98hSj/VsgRtp2
Nd+kVn3OGfZLKT/WDCtK+Gu0dAUjwI1QWh5WZCLF8PQOvuXX5CNeqQtlORjZbuhe
vu66qu7iop7A3hU18RCzsjY1RUPUlKmoQ0hNZl2TQRPzUosuDZ9skLTfeVH5nNCe
gNL+fBr5Ymu1uwThQs1NfKvKVCEy4ElGhjwRa8H3xc1Tm9md9n+94eFZ5VIDn646
duxfb/p9iiXK8GIZ7B4a3UJnzt9CwfpR64tGDCYSa7cTotAa8f6IuzHpHkMiWO+3
nHiO0ElQQ68E6CROrl/vVIB4b1niW8pc/UoU8vqFmGwouPM+6xI1xK/EGGJxHAbb
QTeSkSogSXoQ9W6wYF1d6MvoVJ0YRnj2LlAGHTqHpSFFsS/XVYysqWiRS3DvjdoV
mDn7XHoA4hwpR8t20hkGUiPVUwQ5702Eo3riwVytzC4mNE47pGNsKBjqpvQYeEbI
AU4m2KvB0nUHfx0y/WMIhnMMNIRfpljb5arOlaEQ1ubbIiV9kSvcGCMH0RMZoCRO
VhTqnmAiL+fSr9Wt3OWTwdaqSm5nOmtVrxDDhQ5j48cACI5lGLtFbh/Rrc5l2PT0
6wsal/hcdEKZ0Ko/s5YMKtAkYp4OSJ3QlaYdVRWoSdsBJyiFWcBuE6+54w8h9Aoi
lzoNFXkHMLV9c9+MkD/bqf+JUmXrHs6Mkeh8kwwMDFysXuIBSGxXrMKAHYEY3mUI
11Tbau/sIJrHtTudSsm/Byl+Dj2SQBrFiFKO9gCbE2500oGI05by9pJkgCxmGeMp
npIxvwuYS8bPkroET5aJ0N01U9JfdIWoZszR6xZ8wTsPzI/hYQL28NFnUhcuWWPs
NdFRcaiMeEhQMjuH4NjLTcxmF18Q5UQpVZup5Buss4GA5yqOVJmtz8NHIzUvOqv9
oVVB7R5k2APdyK17O+qWlpFX/nF3ZZWOGG2eRHxL7aA7nLA3kOYAKbVBCWIfwN4d
TxlvZNEdvxjnnGNpUnPhaDI2iwlQrwJR0BANmj1kLG0hcEwf31B3Sy3kUa6gcKfs
EzVRj+MeWl3Zac9YTgtkWzunu/MiHVkZ9fWyisnzpT3zY/dLeEgnnnlD8uVgkbtn
/BugYu3x7x7lf442VqsPQMb6wdfiWydr88LudPonIGVtfNXRbyqiEG6lX5ObGO3X
/7FaFPV/qIxQ4fXTDisj2Z8PVYLtoqxE4f1kCmkgVN0pRKYbZEoToD1PCUll7tdv
R5g94QsRRm/n870mtTrpnpeZKwJ93aO8Sv/LZPAxKiCDY6bye8O4Qv5Xwx/+OkoC
0eO4lIQ2cns6X3GqsmhkxColLiOJqfuIGswvbsSIOc5I/ngRZ5/L1c6ne5/fKNUB
cnVC1rkLgKhTZf64k0kzJa/KNnOSOmN+SJEechoFnl9EjhOg/cVvbbZc8IXOi64Y
wjxhoglUpeR1qBxkz8wTX2mc0NTF4dRVNqUCC9f6PYblNM0F634GJrkk35vMNY0f
FmesBdEgXRLELLI2un/WQnpc7BJZEuUYkjptr8ATrn9ASxtX4WpHLY0xZejlJQ2q
dTvLV7wB1+7ModZQhYmSJ0qxkMRWbJtGkHdk+9HkO3vvI/B6hE5zlL4ApNx21N5G
wXu5aRpDC7yL3gbjqxIVfXEeRqBmXh/BSKPpAkEn9w3xLEmPQa23/znmqrbhvXEw
Uanoqmu12ujrYT6sg/I36AnGVpFw3gNVwPV2iJsFyOr/8QPpBX9jYtjwIa89I7iy
y0/n4Y7zZ6kXQ9/3QSM5behEpIQ2otx/bmRQ20PHFAO5nAs+HArga6rfgn+HlRYy
HE3r3+uZ4W3l83oO4N4VXJYE+qPFWhFXkP1px0Q+8N5QpqHp90cNrcJQWZmDX4eI
H9dsrgNSjYNRVagrqXsvRQ6A1t0KcrAIQEa6+O9aiuaWzd+lvQXmEbD+oXcC0A6v
izk4Y4iIJ9RVAdjpIjIlLFk9LHsUrHHWsW6vmQ+Q66jmRQnxJ9iYsfwbaAgFFW6b
X6/dFndvXaO65UR7l4+yzfDoCj5QehcczA1b1M/VI35vL8B1eUKKjkPS9y6qX/qn
81KZZyhZBOGWCGIjdQbESzW1jd/SDPhvPaf75G+uDfaYeeeK4AAirwqxHcxfkAMx
PzQde1wEzeE2FGBTbRLdQ8oWNvJDJnUgzSjrP0ZDKT6tyGb7NmsLFQCdTiHkbXo0
7EsNawP4RX0s+obRyzJ/MOP2E7M62Sdej0+rk0EaCXjsDPIJCephpfBn5ZB3tNSG
2jlNlMhYZyG7Lfcy2EMYA3cWUaDCBzOiza0x+50HNEFgc2ItQFyKSuDNpDOmJrpZ
eeE4b6N1tfd2Do3Qgo+n4f1goH6mn9On4TGZmfz89VTJ+WRQY6jjl01MovtpmGm2
hGGHo6HV/OGA3127lhYbTsZVzIWaBgCXO4Gus6SP+nbTB5G26VL3VHbf+wGTZVuw
+c3Tz1EmQOhUxLxm1TbUg0RnXYEl/i0F07Dp1PIrU5V3JTCV/BTth/qoqOzLF+4x
uaG6ZPT1CnRG1jiupEo0AiIlioKbPiG+KwS1j5oJRVzD5GrHAlZXRUpVEjaWTTOh
w48m5GVZCN7xCsrJT8jgudryZvQ3uuJNr410S5AFziTUf10wXFjnmutAWrcuxDvC
jjLMTrI/U13ep4XhtEHlNeM1Sjf6sQptM+kxI6+MhovyHbtuhGew+FbV9MgEwPBN
Mzwysg2qcyKDTJniHv8bUfWJX/YjN0eWq6dJD9LyONR7OLhKP8IQqbzdyZYcLRUK
Q/T4tcF1vnb3QWmWAZ5jnZ4QYSriW0MMpSO48mcPS3fllewl0XTLqJv2k9GfIUMc
isJxocu0l6BniERhwmHGndEe4gNXRtycn3diuuys1ItSvaip0YpL33QpZ6/KtgvZ
+R2LZmkE7MjdFskij8sWwuCcYXgQQ+iiXzfzGviYKZuo+7AReuxWszU69abhq9LG
/lbVE1rA1adiI2XEmrttzvADDnO4BgcZP2mFfNNc6DdwQXjMwqkGD4ugXFPOrW8a
19Vk38n6YkihZdKowrsSWeCFXyliPLIdPvcZf7zAxDQoSVJrXsAaO/cQ/5IgEqeQ
IRIh4RFJnfsBbrc/6STHE3/LxdB/fMjZk3AAswO1Gd9V79tUAZesm3y3md4ETclH
04sLk6BKFVPixfhICrjMm6oTsvEvCXpX8qJHgyJFxuRn2VfBuB95GrW2l7D7s8CQ
vuIoT5pDAWAF0US2yYt01GHd8ZxUTBT88RfWt/s/t3qIymH2IwtFG2DnfzXOEq3h
SBzWjhsEjr3NxMbJeEQFeARge8j+ssPXelyv/MU3BZjhHRA533iNQZRsoeJPTFFU
1DTS36TOUmB5tWHPHNqinib2HxbvZ4YRxd6CpgdZNORswvNXRE6Q0Q5Qjn7z5+3/
Fz5zFlR/xKEWrbYwJEvddiInpIdEbcJtuHgpgUeNPbj33A72ukPyd6mwJh2VRvhu
MvBiecAfP1+PuyURLcPl61qVagLd2qkufs6gEMDRuDzaulRuFzgoLmYMRxD+SB7s
kDZkNsEwaKXeBBojUxZa8tIauqNp0Z/wGmBFBY+xTEKK0l1zMW/rNkDorwwha2d7
w1WLBHH7MC3jQkHtWnz/FCYILcmdjA9no0SEkSErgxbXJljtXGRCxNyg8ShOuVxa
mpsKe0W6E53Vwy68yOy4ESYaSVGhFWVD7YLEdn6NOxOO1mhWUfURtK7ATjZ1W92o
xXcXMZCySPw2hHwn5NaCc4avMQuSKfHQdPvaXh+W0U0/fgXwIjbHIq9mm/ZYd7Kx
LmDSVkp+W+0y2AiTDmF02sLoYxFJKv95lCEWq65+bsWcule9HZdG6HmMeg/wmW7B
S9yadNWJwuFHcKayg8U/19GgAlRyUrFm+qod+tc+MU+qYGpPTugOm9kSriuCJozH
wgj8YyRi1WJAjGpqpXXixSOfbfBZSGwk9ONEhOXgHl7FzZ8q/FRZE4uZM1J427hM
Sgh3hSqi+34YB0Pxoip8qOKPqGHquityicDoczEXlDleo5IZTq6dn4CZTzxb80sg
B9xg8i26PYr0bbCgSWMq+za82qczmF2MLcyxrGazLdMYJRQ0tLKwHPmwkCi3byOO
fZqqsQW1ZCiPyCGh9TKdl0KgAEtDGWQ6ipfgQxqIiFtHfVclXoCshAzCxK0xbX1+
XCpt823lX+3uo911D1wJysSQOAHnS/A39cUo6Irr1lcd3Ij75vnCzECa1T7940NF
gtdO++i54iktKyN/ov68vj6acSAcMKpA0LqgZkYfRfTbjllWJBVBw5BRAYgKggcf
p8wG3lAtrXEh8cNhF9d8Mi+CKu7PS0cq1PDYmIqLPuDEjHAwO/WXK8IU1xeEcBje
VI35Darh8Qrc2bV79JgdGajq7ztAbDgYvkj//gKZ7AbjMMi5MctsxFwIa7SVIZ84
GBzwGm9o6DD9u03FQ38TpUQCQBknw9wX8B3iKI2QI40CySeVtD6bBhU8mEND4Mia
YjmhhIO4H6GewO4SkMmY9asZO8EnHKfspC/raSciDekgiFq032sWf9QP4Hr4JRb+
Q+CEmhD8gCDFN6O4APPwSBAd6dC2FxIbjAPEG2bDLdlb0lm/ZxJbo8ZLv5HXL/lY
qA9FOy0sXEpNt4ItndsQ0dTMOTRPbppKs8LWFRllPTT0wboFnzxVbWK4X+7MNOV6
V3HMH7PsKnC9A5f8h40WqZqQ91IEpTpsgKGaJz6n2CtYb5JPfchQdK4Gcbvv387p
gISoJ1VVSDEFrMR555G+nBdCUhJtkZpyWSsV3SIwEVGtFsM03xNOgJY3yVk8707N
DXZ7+HlOIobsjcA52Moc19zN2BRMqEFhF85iQsvdOo+eoGm4eGaoaEgz44enhxNu
9Se/DyxqU9CTQlzeNabSlvY0fASECARUs52pZCHYV5eZth2BDtupxIIUBj3tOwr5
hi1RdCYUgDMReaL/FyKCnuq+A3RIAUHfJB/tt5cuL3xqtLys3aPqX5PZba9UvRkh
YWpV0ZHCgHoirSKnBYCmuyLmW8enoIWWy/mhKYrbzNUiQOFu+gm/dgPcRt6SMdgu
GT/iK46hTZRduzAKcSS5zce0vT2RuEan96NmpK0GzFvdhzr9ygZ6p0XhOK+hJaSc
XRjIov9+Ice2VgSzCx8JGMsl9nx8hkt3hoR7XgIZr4MN25xokvRdfFDaSAgjg+u7
jKXFkPJHb1J8zY2r6q7EJSMEAHnySxkLha+REU3Vc+Pu+wzpw8xY4eJeUUNr63yk
pmbijApssuGttF4N7NU2NzHXRhOVc8JkBE6P2vECHSs5gMDULqurVZOnb9K0u+pZ
XaBGBFaPMEKlHebnDdneVe+P8OUU+HW7gBIPzLyIFAz9Dr7QwSQah9u/dGq1god8
1oyXyBMpAHA8O2EU4Z7KAkkt/39WAObbQ6Y/uDpDMM0e1cXH9HknYfrzjw8vPiRP
OSCENeR1rWlZtLES0yHu6Uf1sch0vhInL6QeaFLhPz5Rrk38tc+fnL+u1AOkvnjy
vcHyY1CeDzCzMAzc0RxxpLUR11lUl0yjkl6ivBk6qL6VW04Q0ao8GpUL4aQuyVUn
YqcHWs0zxKRE1H7gvjecDbeAhTyQeiKoxnGsmgDi0fHrKRzsiRmVrfKIuRBhBaBW
dcgGnXZANyIbhNfPT5URlvLVQcBzOUBO6bSLUakF2/ARNgQueXlF5nAUKUKKXTIQ
uvfAklshFWyqmrf6QBfgl6fYTkkgsXNzw08B+GM7MA3nLRb3p1rPHicVS9h+5ma3
LOkRsUpLcqoBck5sCJB4a7A4/SG7PbK7CpC0hh9zYl/udG9R4RmXoEv74+Jpir8/
kCw3uoAKxCq3NrMoNpBW/rKqLMD8vTQBo3mEGXooaeubqGDZN4xpvp+blsO+vXQk
+j/TVsuCoxHDstc60v4skbT+4PEmpu46QkNXtBpOF4epi0STKv54dOsbAK3Jhaze
NrgY+SriEIqeNvUUR2lYAjzJmzX8azSMHe5TIldvpuDdiSBgWdPuk3QSC1UjJZiN
k+bgfekvaTc3ZCaa3sOijkxFcGtTtF9e6TwO8yE1eXCUt8MwcpCr5NH3nKI9rOKB
5f1pc0E+6W4vdfS/nUKJMQYZ1KtAklmbFQDlRqaJHeYBoCh0D5YpqzYUiL5phcOO
pRbqGg9p5kvkZZJQj3SfT8HgdvoRnlsc61z5KTWbYcBA3W8eu8Ee8DCGwhBDGBgp
6HzqcXELfCUHdizsAW7g5SnbOM1haEZ5uDSPYNhcphXXQu9IgCRbLktbg7TE5HRi
6+ZLc8owWVQ3grWDz/wuMbVqtuu2Ku/Ka0a3KfHarQJIOXHZt9YcgS7F3C0SdKqN
9FCy+b+CxSseH5Xlq+IFCaSzJyPzd/ezUKPotwV3hpRsvHjoJjh7b1ZkQP3I68eD
elqNhqCOdYIrT+u4HqT969uCoHvcU5yHByxlHRz2pP7aTgodRI0RsN1FmaHviqB4
5sJ8atTzuwmtdMfe/IDJlIN4pguOVvw4TV8evE0z2aya7yXG1S9z+1V4SU1l2d6X
6+ykS93EtYpLVS+5R2SjOsBX+uctPd/tPg1841Thja3UkJBo4rjIuJj8K+xU7JiB
nhNSfBGJUJNQsE1YhQkJNgR1jTbQbgakLkYk2pMwscRmgyfQlzXCfQazMElCQSY4
BYOH0nmF0pRGTfVHITKJvGPWfFqjKwMDJ8B8terRY0Qx0XigYsQGrkQdnmnSUSJd
h/PTcK8FVPr39o8qIZZnfXsN+xYDnDOrjaws9er1qc3x/wQ15tygDU9BDbUnmGO2
WLOgEcdhtrNtzw19oRnwg5wnuC4uLVq4oh78EkMUrceQ4prJUXmaHQlWAhiycYn7
UYpIsvR0Iv2pnEculeUyLc9N4o1kLXvbMPEIVzR6VYm73f+GpUinpKVyZV3rq0H5
BIsSAIOmDKZoxO/L2g8mhSqg6+FOEVw3MghYMJ2qco7mvhdAThY56x5LW2J364hC
YlDV+1Uo3hnDV+JCgEAYaR7D2FK+3AwOF4Xvsj9qZI9xczC6XOTzLcc5UhQAGolx
djHqkxJ4uUFSPONHfrghh88CjJCzU3vfHRzlA209oQIiiydmOYkIuGE5KvNVb6WQ
oHkr9IHWPxLvcHN30ubHo0htNNTjY3vwI8S+W0x6j8O1N7ggDQamPPc2GrFINJSX
ssznK5izNpPppI5Em02r8m0FWFLYSVci/hnL5msL6B1EJASu+LpblbDowIM8Asx+
psFZOrp9UOgeQ5UDiSkJd6f6rMx2zcJizxTnHabUoESjn67UJbwY6z4GTWBB1NMc
AiJcY+wZzPkvaNbhNsWN9r8EP7Rj537DJFZq4GAeAnxQGBIPr2zKHhe37DxLNnDf
8VbwoJh1nUJ9yWx/jn4bIGIjFLIN+SBsWJmCTgNfC8c2KQqfX+GPnv0bpRCR2DY/
0WpT9ld+X1dKGlEJcLRsr9F3v2e9i/bZSnJen9e9xPBWaLOgsa2tDq3w/SCrdwY1
LhjDF3xw6VzrMUaHMe8qs17xOsgYWag+ULP0g4gG6ogsJ1RmecrPBdHJuxT+Wz9u
uORlImM857dXjnju2TqIYbNzOLT4fDuRllgVmZVjYqa6s7G1RocuxVl3EcdsaJ9D
7hlZ5hQE4MF5sBsh5w/6K3XKeJUvnKr8iulmPwDHP/IVzPQCF+ZNvd8FSEtxOBC2
yfHOvDApt2+DZrZsJejW11xmYgzjidMJfAqzIWcDGHdwFUoxye1c7JHVEMjbFiJm
tlucQbRbSsMvkzb8hTVPS8Sdq2j+NZHSG9pmnyOkA9PrDb0TX5Gs7nGGkOEgsyme
xgGAJoM0QzVyF1thy0SRrTsK0JL8FXZ9kocYkbNHDqZVHcfigZv5OaomyJa7q1Cx
zD2U2Ru1n20YRHBYUtVVj75Z9rlwa8/FL2Uv5JExDbIwtF4HQT0FFTOl/eDqjYEn
kDRbzVLeyYfTUAYZdejwIplNPOISFfe8BL6uU8tepE+M3K+9pAnphMJUbfLMsmdZ
2tc6nEhmF9e7HxIZ3wOLqu4S/RS+4v6e9+xqKhMcRT/QbWuEixgQT1idCAD8qkE6
QroBrKLGh/mXR+u1SqOBuTpj7hqv99t+M36ya/GHHXRFb9cgaEyoZffa47ojriqM
WsEWHakIx18xac/osQz24TH+U9Peq2KdzZMePVLB1zxpsjcGyRJTXdcKCl6Hd8eY
3EgyJGXTx294Le1pSg3SfaSwO0iacxchdo1H18/8JErW48MgrDB5hD5c4A5k1Ji8
6Rrc2Qe3AFszNtALt+jHjYSj58QRTVhS9z7CdkNelWzn9US7/jW/+H6/YnDcyr0z
Ljn9S0TaVk/1FnUaLiJuGf8r0q++J6eloVgMHj0rNk1Y8M0sfSqUnPKUl6NTyV5m
o/ioIksnlJ+4Ka7DXAHglKT1BKioZcDlV8GusEMukalk1vhLpuO9it91gtFYi8b3
uuejX60DJwlPkbbFK8vcoL59vKxH0+hOGverWLDLALXMR9A9h32Pr8CgHv6Nx3Ss
MmUAjeYFqw90xy6ki6HpQzm8lgXQveuIvdmQSCaapd0iqfS+XQt7xaDgjo+ozZiU
4+wVJyRDKPWvt+yy6O2FbwaHn58INGYed1nIyiQHKJJhZRhKhcWCQrFKp5fdTaQh
fUoWOZAeGSVJ4c/ez5aP1n0392RDTPDpRrt9FvozrUKgz0TR1FiHguO82DaN5gsR
7L877Pqc7/uKeR5X3FV9tH3E/zjhltR0Zepg1/aDtnrmq3oDWH7kI8s9llmx/J1f
oUEC4WaeSVd5rxVbPxSDo/j6cWpetw0AQfptT6/qas0yCZh/wY8ZC0AD7BGl/R4C
mwvMa7in+kjRy97cil1eVeL/ikVw56f8zwBNZbQyH3FrxJVITHaYmWr0tvzWE4Qg
MoJB1RhyK6nSaDtffWmLWnY4l3iVqHpS2e7G7cvbKmWkR1FdKaYO9OogKLFlgq80
jYIbl8DcpHWEt5yWzuK+rbsFpCss14Z/WzEqwOsJ5u9/cTsomnycY4j6X3JHfcKV
q7fOi6LexX/6FDfZaZULwoKfU2USTcv5yXUaAVEgv+/aW0o9n/zqhSpZtyzATB1D
vwjxRp7nl8AGnqdYpJ3OrGnltm+CeD3ODcp4TlE4utWY/CymrU9UGElAkO1jlEHT
e2FfzMXYNAI/W+BuAHleusZm9XDKy7EhvZOmqtONEHS5rIOvymjKba8ojDqA0BUK
ADX8E3ZLkipGO2xM0tse+VXoxfVvRJEzzigJUc9soL678xN5v8yLPXq3U/3tTkwt
JDG8fslgG97SII6CwnZ1hU+PEdymzfBnIycKdVeh4gaZbkyATvv3GsVyl4iYhcYb
wZzTmLK5IF4+k6nEtVdEF/CjeZKAOfwVWmKlb844CbkPkPe0RO5iMSBNVg8HxqKS
VMeuLymWlBFQ00MuN4GI7ALthkn+tTVO+Hut1ChfhCZ/ANiLfkjWRYSjxh5psk/G
x+viXXZTCW6dOgqe8Abs9yTDO9W12lGkG6jL0x8Tef/ShTa2mSMC/mhYyI4YVLgM
+DcpzYDx1KejOJV+qqpTonI/iFoTF6I4ei+ncdVGgjoBmeiZlFE/kHs7m9LuT4Bb
dbvTjADu6yHwOSmM4ikzIH0K2gFkt+khrs3RNee9pq8WKI4pNOmqU57yB+di/OB+
xfFSj763u0cI2+wJfWAYon6fVfhm/Y5vf5Z0YI+sBkUjuOTKygh10G4ouDoxtMjw
glr24XA7NjI3JIghT2QdrdcxwwVdYh6fMVOc+11RxR3UG8QV0DfQKZQ8L2Irf/pQ
YbgsqHb0605UyvDyOuwjFTpH68BIV1aFoGJt+rVCN48B9WUDI5uo8s8V7elFENsk
JaWk73ezjtkuGE40wUDZwl13eQnHucK3Ygr+u+XNg5MxeT8wNHjjFrqIToJrFhWI
Ayc4nG7tJfI2gAcTlIpnDgUfaYjx139THe/mvBMaSPUDKlAa3mSmvr3LslrczDuL
DTYWnTy8QsS7tgr/b/SvojbJpiK+9lbXOQhLJt3LgvlJOAz2V5lTGqfxhdVDfoIl
92xbWh53vpnNfY4ojlMV5c8WbdtcbowCSJWcpZxbicQDPkAetc7Ap2ki6mhp754E
eTvtgHGtxm//Rzw9Qfd2fdVkabtgZf+hsgNTVPVW/FV8rYYkNYm7DeTYkWSpEWOT
BWI2NJ0jpNx3Mr/yfkEWVzh6Z8+VvjZdeaqrLpqjMH/pc9aEJ7opWjOUcbhEaGen
xqPCQhBmKJ67L7SPwbs60HDyd46+GemX2jDxsc8b6qiRYCVaMH8o7S1aN2UJlFlr
3J5rWXn+DzEoToEYV/QHj7M0qqZYXX4ZGv89mqDj7awvB9THaZslVV7fsIsWumdc
B1OCivrGiflF8LYNot3fmrjN25OsITzcbrXBXPqLjUdSXMT62yEwfbBPdWzVdZts
yQK6VVgkhyBdEmH9y6LFVqYPfzX2A4xLqV0Q8+Qo5tXxXbFZ5VflPmZrJTagWF5q
bL7sZUhlUp7S/WBN1xKZGTycRFdOTqAv+iIbt5h2/wQcQOxsrVxMxSaJl9UDEOU1
9xJaIwAYTY+axT/JcPb/ppilkdpd2LJ6AgB2kknEu9xp8FEd2wEwo0g1Y7mLKK0M
XFU7NcQJVzddpMbcUg4Gh+AHWhsHMs4pMg2LqPQZJXr1zd4VMncU/L5+qUThB6EO
avfQOZmbe4eKd1090C7gsbMyhAEVGpoxw7p+Tf6pwlGVrL8jDoNsJObDvTEjigcB
/mSIOCR+Igs3ioZFPZ4C3MUTB7hJGI6v1w5CNr42TTkkckvJ57C6xioYp3eDUTbi
EzFaUAIkA2NqlsQxb5RuRcuchZ2tAnNSLYdlF45EwctpLJFVJQ4q0OmBWtmNoD99
2m5X6MlSArmp+4vQMuwVEikRkqkLIk3LRpxK3t6e2/3Lwr5mm55gwGyENl3lkRYI
r8oiFfzBy3KIasuY9hIbB+ZeSNHpjRhLEbzD1iDh3XbKgVAwyyUU7IY0XT41xWh+
drm7Tf63yfLKD9TVm2Z0TkxGOxN8Q4XyrtVWY6VZ9LinVek/9TJjSacntOrN4AoI
H45OeHlQ0BWkbaLAYLsNUftSx/PJ7cp6mu1GnRvhLHZNvdxQrydiQg0G+f/QNST2
n4iA9m3zAYo/6WNyn6m2r8crx5Fn/FRVWdryz6+dEhHJoIl83wkhZsOsGkFsJha3
nx7Q175CbmskZsiHpMkmDHB9OSy4OUyFFtmOSaCjObvd6bodUfVUbRw5iDh+jy1x
YthmWMvyk5kfOQJ03w4DqSlhKcKnWnXSkiPOcz1JYhM15pbTLOoQpCJWVRL7GBhW
WH9JHcVrI78t2thrbC+1T09BgV7xMYwZ2qn4RIU49UEt+KuJys21i/+bKljTxSt3
xmGS6fQ+hQbvN6V6PGC8njhGr6T1GC2E1zprcsuEfn43IMD6aDRutpwuFOpNzLtb
/rCEOO2/4wHTx7147eMAuBSLvH/HwaxuBYC7icQC8dYiJL5CZ+6lK39Iejt1+rsc
+VqSLqeIBJpq2AdaiqLV0LVYEdhyXMYWx3eTFPIRkeMXqcqQZYMd4/Tx0cTFHKNM
orKl/ADAKgDSL7HwU+MfLY3v+Nbafw+OlNYSQP0EM2RPC/pf65HdYGEkoR5XzIMP
4nFbGLKNlvxKlpjxSw5+KmcEUz0TRf4UdKaVk1QXS4V5ORef7BUnMedZonGrqpfm
RN4p62fy6og+LgGbxNXpA2rfScRCvy++faNV8qVBloeiqr9+mFU4vKvXHpDGgBdJ
XS3wrpHONy7nXoxqTZK5CFF9y+XDJTf1I7WHAc4ozHZvQ265qMvDTivBb0tbkhbh
0uzvH3tPkOoYyM/hBJynmrpG8r5bCn5+aB5gFo2dnlFgDDvzHnq8/vGJIwVkhXHB
SoyVxUS8Slh3mQkX6eGap+vQL43ZGK3wi14dlg7GHgM=
`pragma protect end_protected
