// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UChZWi/xXNilEqrb4HXqJL1+jcIbC+qQvQH6evziRXT1skh25j3PcXBd+GdtKwSZ
YlZZA6vO9Keo/t7eT80OLdhz/oaUy21ZzTN0z0mCi+bRmF9ouMl8XAo1jqdEtVJI
h/YZ3tzfuYZHKG6H/R2RcbvNj0BshsL/hFts/Sq6Wp0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12768)
Lzi1vy+eNbNTqHxQwN1wjYrOJbb54ORYiY3W+nJD71lO6BRLmRSqTPW4qv3pY2pW
UZd+RenuyfqxP2ItGFYyz0g5RkTotxK/rkdKcE4FN69Grk2WVhER/uHXi4wxNqie
FRdlAlq6LRWuyh+hKYvP7dt+k3p1/r/VzRh45RmIjlR6RNMfFHtRW8+Tx8SSrWmX
xAXAtberz9CVLO3qHd9sSOTqFsurSKlopJePPxQW/bP5LOUy9x9GOiRTY3QEK6jq
7wXnlEPCop2QKskHChhDNKmb4Wda8yf4OH70wIf9W70vEbNo7u3CheqtwA/xR0lR
R9/hWt2CJvJKAhd/PrYva5ORjt/ED0qHv965o8q2d7yBCMeapdhMLOHrGzCXsRkr
VAuP8gk4VzD1lrCSWFjxdrGZMdGh6MmDcKDjpZnln6PKbIPQz1WQ1fwa4Ihbjv1k
1/tlSW3xNsl6OyYQEv+32vuSIkx2r8luRyRcfjup7Ccezh12R/FDA/hu6ayEWxEZ
eP6gMgoKUoEuV8YoWj9clulUQNUk4oTh3P6TDZMgUaKVFbDvIBwiRB85G9ARnqDO
zjtZChHockcpjxRlZe7EOuDe+PeIx4App10JrDfmk5SVBJTh6c6DYpePXDWUdv6D
yvrjSO+77Xx2mbeZbGF2FWr6d/wTpFo913xhmC0o4SLpH06jaPgZc5VYym6koE0U
so2Bs3Yw82J2zmtPL51c79Ann51U6UnFk3zWYCS61ck4r53XoSOlIXQpv3w1D7vS
35UCa2sg2Ytvi+SB+yeUI+SS+pNM9HhcR84G1KrMqF+bAHZKzIeT6UFpZ61n+RaK
gakdQOCJKxugOVUnra3K5OGuzFGWIiFajb8gVern+ucFzQkoI5ZSZ4muLKB22gwR
K+4H055xkOqLqBfnD6koqFHbfpYGL9ITxc5XJAQ+X7XErn0UjTFNoLclUqn5/jJa
oXsYyxQ7JYMHuKJmi5yCPpqCfwusXbP79w4d2kiff921Zhm21e7MXH2YVC/bKIMp
ysxpX1BYtGcdHg/i0zyloaUXV9mRrwhHwDbqhYZch6W5c3TgQlUOKhT9cfoXoO8e
wnQOSpwaeN26dTXP49GFehWz6pDULHe1Z0OZiQvx+QFylmiB0RVYChzkCC2QI3Eh
3ZoaB3W7GYQedK1vV19pMbZAKupDdO/QE+/gRAQy5tvIo0eu77XeY85gsRCTMlFJ
veq7cwrmvUDGMMQW3DbQs223UOUChXtJ6bpgObFCVKcTDg/fJ6C0pSsuPXBq/Bbr
vxvpZwWbIeeJfcEUTGDnUo+dJ6tWFYyN9KhoKJb/2UdgrRTZ4wiUMcGZat2kjpkm
pyIB976gB+nioF8ORxD8FRT+fQODnfy4WzBKEHcu73Jd6Fq7Uq0pBZ2MlrUwU4B1
oAx83owUckukK/M869gESJKyWprFMCgbZ8/mUzWI0scMQITi+8Zr7YHu3audxjhD
1saPKrt1AxNZP1xKNDEnWjlUx4/Urbh7YDnCq/NF0OoGL/ePULyn8M0lxutaw61x
UvAZdb4UL0OiYl56XFVyzJCGExE9UdUowr7jS2UTTQ/Z+GGqNp7VYwkmNZNHqt/F
4AMsOdUxac0mkVXPmvRbtlUVt67xoU0HV1q3QsVpijhyN1q7gK96VuGPfm5N6HBv
maA79mtsRtmxSooUudSb7WVWOHQYYQkzEi3yOgsD87514enxreW2RwRFjQ5OQC/2
bi00b9nfDivW5GcQAt2HehrrGlF1uVky0H0WMC9T24tBiMTN551BF+Bq5oiEcwZo
SBS/c1eG+fCAfETDhta0AGcRQibe218X7KNUQyB+gW220c9CDRjoSbvqtRKrRkx3
fLsxIiDC6JL4Evr/aBUwvm7roylqQgpr0V8YSOgv799+QgpSYlcZi/G9RteYIyhh
8r93lrBj3uJ+kR0NjmtMMBgYGJdxwSyb/onbO5vslaKlMuXUi6Nc/hl0MQH/xVH4
6vEi2jbWx44nmY1TrUq3eDlHYQAQAJ5Lo3OOtaQW2b+UzywtX8dA/+l8G6/iWcOI
G3/LS6+QJozvcl+cO9ciY5JMLyehPmqmg4GW3OwApz0hWmPC6vd/Wctius3T71Ty
bALH12hjZ7ZrMxC8lRuvFYjYU/417o8ZUGu6VRnz0+1bviXsLrDJEaxoRuhMEQWc
KE0mwJcNL0nPErAveu+TD/7nbqH6g/I8YFOHpvjpLB1vHCmV8aDJ6x0cTg8c+XaK
o9zic3Kpgx4jdK8/dkVlOjGxiQ+FoaQfhJ9JPb7tusf+Zyt0Jmy7aTSIdLDTAOnU
zEOb+GJRECA6pvS+iX1oRjKvLH8pa5alEsP/6JYTJDEQpHtXfferOeZDrXQKuGkC
Er219p8dyI+73EsBfle9D5lxZCJQGDkVMEMcCRDpTXeadNj3+9W7UMlgQfVh0Vo7
RGvP5qMuz+FxMuxWOKQLuOzfWfjwzqAUoKKW9lyvk6GV+Iwm8RWS8LsHlNnmTBYd
X0TmVIDDGmmL5EGywI3GvS54YBydNikn5XDPRpWGhChFLgoupiypkkeL5tZhyXI8
Gs5N0NWD4nLLZXoLdYtSYm2jePmP3FcW5d8/F/qBMUTAnYjVb44ukTjKXRisSUf4
Th+hrs7+Ej2jNgML9/R058bmPmMZV9+RNcGz7gV4avGoFQujBkt/oS8xD0M6SSEo
S9oe6X1qAeFBjEpCgV2rPg+eayAbJ0JZVbzkLRsotnP9J7N/W6Uu6BtXWXcgJW9g
SMLFRfjt8/2rfi+BqdFvwrYSH+m4Lw0PrOTOt481kz//kzOuxiv6qMi+5hLPJ2fJ
+CnxIEphf3ojsBChdjZ58CUWlbP3bavst60lteltwDtphypTv0M7/ZfEzZ6w6UMf
4fSNgjRC6bVjtTB6vlmTB5dx5S7rxhN+JQjuJZBAZWN2O+Z2q0gVUJULz6J90PxM
GSeQjm9NhoE1SCdCs0on3T0YSzYbQXOjkivE0elzTrHXywQvQPolPkxuunLnES31
8x/l8R1ejLN0KlvvCqPLBp3GKXbn/DscSHvL1mwyoCe9mv1ScT5tE/7tsCmyOGsC
Lir1klnsFVHTfKrnmTPWTjEu9MZjbuphFOTE4gnFq/tJcCsDFe9ZNiGdRflkvr5a
KGJJxXzfjwIMW6DfgCj9zVjbVAFjvdAX9ZLFNUKr2j+UV1VKWN8Oro7Z9obHhi+p
j7eTv3ZWQuHncEl0JHYe02tapMnmaIS91ZdWXvYeTRazOD1XzmFDdgADe+U7IZAN
ZbQAE5uystgxNbic50YnbPn3fbUbEZZrnVz0v0sLeYmc3voNUNwKznrep4/gm7bM
idsLpz5G9UrpwuHk7C0jG0ASyb01wgtX1GVTU7vBgjqD/R+mOEVcKZlJW2Zn6IX3
O33k9cYzKs6sm0OD1iBFGtR72Muom2+8yfDDPihmIEGJ+v84gtO0xElMHDhBX2tm
SuRcH4E+Emwy5jRPe4a9ra9NBTBoP0xvZx1RIXmp4cy5ogF/DBsORMsXTsENUp14
bF6Abhk/AEVsIUZC1NIz35c2khs7uI+xnSQMkiDlud1W4KtJy1hmIMqNtSlNC99h
ifx1f8CGUbQtm4Zg2bUKpZ5qNjuO+kICbg+bni/orK7eAnB2Ra4BkOx1UAYS2E51
QnWmA/urMH00rmrv27fCGVBC7q4sKvFVYTJisrQJjH3e56CpteQ9vJF8Bwo5uLPF
dVstoFLiEbGVLREJycmqQoBYaBx1gIQSEEsDQBjB5kcAtVEAakvPIYcraFqILpKF
wk6aGUmIcDeHcu5cY5b59t3g50+TOWQgcN3LEQEOE6sDhxubFfTIxbTkPitrY5Q3
lFt5QMOzKfna62y6m4MXoCB8V2NGoNeddQM8YOvwQoTkE9nmKN+HBjBYCZ6FFcZF
qQUwzUBybiMgv2YFfTV0KxE55fpD0d/UEHyeh6JZK9+9/QwMLr6mfI0lyacobirP
YPehIzyACDL1hShiUoOZm+GUVvRL3FYEIpFl2VEn/eVvo+EN4VzT6a3kHj2KuA2o
hTFPesaDw30az5B6kM1o4HDpdnKZM+Odq4F0vcnuIhhOYD2U7P4jvrr0LyhZpAJt
iU6ZOg1pyPkrHiF6H24fqXvRzgdJ3UIaR0x+MzoOurRYaBmJAwlYi+PZKmX4515O
khAag/B00mJe1XgdGVoJcetygV7uhg0IX3lt0ZmhiJevtuqab6v4IptUsFC2p70v
3ZVfm072unWSeIpsdG1nxQtxFrbH9ohF/ABPKwKZNXTKiheozBbzcSQaXL97YcZB
U2JZ7QetGOE73D42hNtep4pq3j37YuSMGEGiX6LAJME/rYBZn66NsfeFA9R4giWO
8/83i0PDez/WNHuKDYgpQiTyaWGVPRHdDdjwQnhejKwQyUEaBTxz9leOImL6UdE/
m27hvA13s+xv31I2SZMWDqNEJhwDW7cEn6/I18gRH7go7eyHZkUcv+BApbBtYK1q
MlUg6yC4UjJDSd8DPg46gGx5dncpmlc9UGG6NuC0/GbHFKnzzCLMKG83pol6dIj1
2Gz6FSsynW9Ghey1mPdWpvVxpsZGprwz4pMep3z8O7MzYnUQdrJDJwz+69wp1yJQ
GBOPJtHYKHRtXJeTcSVG1d/kC0wdcU8Gn2WH3fpIAcRmTZ6pPIjcISw2/Y71+14r
l6UwAH++evQQGb71XJcwdwrgSGCI/0bUPg/FlGhy0750dZCjDFo5jKOxG3Omj83h
LedR6pOO917KoEjbs+kx5wQoS1xeDS25FEm/YeWwLus8cio0lMowshKb02jOM2Vx
WZ+OHKRoVzYzBEv5SX2zDRcAL3+dJ6S7cCebCzY4D9rRV+IvLjtuEP1YN4bz1lI5
AT/lXfNahrkUPBBvbMmU2hb/vfQ5tdS8H+W7u4RxURraBEhwfuSkcNpV83QlLgys
SjMtP80iFQVoFw0cIrYymMRFT0zOo57xp58/FoYZ5Eq3AEYfCzRMA1yqdfZf227P
HRCS3jOOUTGHdfIr+fzNnrugyNz63kcYjDQJ3isNdesEmGmSl4dZKMRxY9FvBl45
ufDeMkD5wLPwyDRBMJ9V3opXbWHHpgiTL5ahH1Uj4c1E49c7TPD+mXisWe3bcjzM
paXNoNcqSzUu77TiowuaP9SgXfltNv6dUqURC8NgPiDETH+bWotZfExAW2AnPPNM
l0Hv0vcAqzvATfCSVUNd6woDswgwQ5VZcUHTOI5ALrfHI9PqM4XlSEiHbEgL6jA7
+4DtV71vN0mX/T4fdKZ9nSDbygIg9h7qePILqysEFi/EXt+w32dRbxovPR9QEwXn
0l0Ehy1Y3KRfcJcNRVUOPEJmfR/5aFiEze92HtmeDanJ1BSNDEJfauIQmHbWSM8H
whHCox2C98VgX6+nNPzVbPkLShKBUZEMuEbZyKANwS8OmfbZYpSdrbcx1VVSam/K
V+TvEdjACtjIHBkJZ1pxDQ50HkhlRTpD491D0y3+619Wju47CIpk0oGtB881yYzN
nkywFHrTGJMsj4YLqJWhDH34t7Fr9pUnG2NJmFSELyAb7JrxtSs+qSwlYtY17SfC
NioUUA7VsbgKf06rxuVyYm5OhVIMka9xYEqzCk2U8KjyhEiShYkehkBaLAQrLT6G
ZoJAUEWZfhiPax8m4IQgPzXwKE8CeOgTeTnH1eyFASstujQCJ/hew5TOvmV7VNsU
7N7diTQ+TAz0nA+zVmKVEx9RaJKVRe0ZPMlFiljzY4tdAlV1lyx3oETFsi3b05Zl
TX0yazPL3eIA7Wt4W95fc1o4TTTejQu7Byu6pdQWH3fQ3eyMwliQyuloSMT3c086
YkMFyt/vttyJckIQYDODFIum76PHe7BOveCV5k2YJNKwYUOJsN0MwACbEVWklkkL
SPov0u/ZjVZ92G17A7VRGlxSwLbLnqmvjn2DskEjwVi3v26aLbyeI12ooVzq/GDt
2vSO7GW9egoSdzd4K38tEl2g/3mBobla5Sbg9g13z3wY8BOAxPR5UFFOOLxsw6Qs
apgY4zZrNtBjj7WaFnctZ5jNC8fqIjc1re94wHLRSdlH3jZrjZCkFGyItD1ew2WC
iIb9JkTrcKYxDHsXajfvOfGZxKJcqAK9GVro749KoMm1VMx0Mf5T0dDdcoLiusLR
qs1QzubJ5rhRTVGQErZeq1RziS01JOOJyL68StZnySgYdJNJUnHnJvv9u4oM/uuE
GDLpPuKs0GevqOb2IgcD6hR4tMauAygxF0HfZePRGxSxo29VoVhLfQYTmnLDITKd
Yof0cGYP0b7/Ht2zGwVcesQEw0Kf3k83liw7irwP3ekHjJdCsZIWwZzWjGbq423r
vJjQFCYh5olcOAwfPYj7Dfnp+qpmksvHEiUfxDex4PyOizJm8giQ4Elr7NAn9Trw
HXhDemt86DRbqJ7HnigylORRlA/PofXSkgFI7fYP/flz1gsdtXMYbQjgWVZd8pVD
zgwXuDuD7GCaZSPEJMF3w5NUMRJb7Mrpmb50DqAXLb1rAeac09yJ9r/DBcCeccQ5
oOBNsNSb2NmdMHYuuHugXGUZV3VAMrn+GkskTsiDzd2VinOleJniIzPO368NqP5M
ntzdK71FEE5E202tWpAdv/X4NOcpYdTz5fNBqKi0K0tKQkPcr0Ds6NG5D7b8R5s2
A8x5z+5VHK4ock1xmDf2AJrdZSzG7LxuDm7N8x7Q7qM/gA+G0JOvqFINF8jiAYfI
p5bItWUwbM72mTaMWEOPblur1AdHVeDAKWI5Qrf/r2fMPnsFSz+7+8ogMMt4Ng/7
A0Twxjw5u06TNVuSnyXg7LNA9YeMP1HkHkzR8VkIGGol4ev5cPdjmc7681r00a4o
SISEDQPa8s5XUcyZijF91SdufmK3CqqgvCdOieIJCP8RN7drmYHZsCb062RshoOB
AE3Oo9732i9NLNAXSohYJV32WyZ4eNfvwQqdsflRHtZ0nQjoktYa7schlecMzGDf
atM8+kebVJWCvCqXO1cZOHUwPji3lS0lgnek8Af2erv0qBmzaHfZG/DxcmB1oGrr
JOOzVL41oOQYHHH1kt7WHGSu8lUpwCgTAQqyBL5KuMthEaa527HbLM9iyOCzKGkH
psfFUXL9I9gFyb65mc5RPm+PFWc2Q3PqXa5g1+4yK63u7W+jATARdo1fsxSvamSq
VOTFf2Io1cno0Rf77+1LWjzGLY/sm/YJIv/+bpzpVj/GS/S2gKUN7fgJkgbR/wud
ij7aEP4oaw0ZytKHkhGqnXuarkzjm9n5SIB6jgJn/bbiA13pHC1koZhuHUJNPv8k
6OFEMnmJ4iJQCZr+J9YmqqLBLAahlYw0hXleKYWJrzLdz8fA2R1xWafIsczd2GKv
tO5lbnEvcrGkycskQk/Wl/BuJ0dpUULfJbxSAMHAia4aMkqvCWV7ERcoMOhXTx1+
GxJPzNaagBM8a2xhWUkhG4OQ9N4lGomGvnoWd/ifBT1xP88SqhLHjI3q2WbN6F7o
IfEFFjmq4b0ex86diQGr+FjdZDjZEHnVvHMU7mEdbU/wsZ4aH0PFjoANL+KiG8dz
nKuR/99Rxk7edDqCFHBacLRxglsULp94kWMCZwFGA2e1AuE2alZyYIAnt4qpK6s4
1XYTHVWBCTm5SeaFoH0LjywoulKjDPSlNZqwOkEW7m7tjNfNeK/Nw/QDZmBJop9j
fqGZhc9AHaksIqiocvMG4D3sjOIHxCWFkFjw9Co1RJMz1B/4F+6tHx1/iJtOpq7L
tr3iuDHXhgfuJTnxPkQy60H4ug+voNT+/0j09gNJtryXJ2mHxK7N5RbabqpH5W77
X83fD8OJY2x3UZt3FKm+vzop0cPxkjocE3mwsCDX4Bi/DchzAZFs3eJr9cN6SD6F
FS8W1oR6S6HgBIQGSOvUqXYCfOlaVQqJ+XJG1wSses3FRutwiJmMZ3EsX0y7cVlD
v0eMRhZITk0Ikpk1jU9cHZ4VUBZsuQq19IdcX8NekM/VPlN9EzvdcbT6fkDD3l6c
gT9JjcJOt3kpnMIwSjpEimtEFqWaVEQeri7bIyWBIE/n4Ox0LQxIPItTZv3iGhNS
ApzCAiHbzIS6W9Cny2IoNpuDQHY3Lyrn2a/f83F9BOgWivlRNlda3W/wcst5pPmF
OJ18KhovDgmwiB3NWwwuo+vHbwgT4JqF62bnBA5SrU1yXyAoTeLtqhFnodQ0NOQ9
4BjVGtyk9FGGJqYlw/WJduR4iFFEnO3z3rxs460LXzoXSdwuanfLalOjh9uAwvpv
aDpF+4YBkhBAeZe8aYvAtHfIchh1N4OqucL/cRtpv7JznrqXWcUZ4SEJDhUTp0HU
A1/fazEKOxgkvPyuEMQm3kkupXSrMRqlpy2c84zKy3EUDvVnaEzPKuqnL8+yoAVL
Rlm4Js9X0oFmGDO23LBgStBGuS8MX6yWtPgXEmKBTbXh8Q3p2vuqORGHTMnh2bsR
iUIH7TsO4HhqMfAfNf00Yjxdy8xmp8uVoDBTlByxk5L1B268AT0aWAjc0TFGpxfx
15++qPY0KAm++Y/nuBx80RoRjDQUAClT0guXl3OGIZmP5R4cL4O1GL9C2Di7WNAS
F87SWbjncS5hlfGal+JIV235+cOxHcvZ1y2DFTvTM/nDEcReWopUCeVkfG+n23If
Qc4Cd7fF3JblbaEnOuqkAcSGugAOW+D5NUeG89H+/2/sWKihD6SoawhAREFNaDic
oW66IliX784q0WwaAkwJLFIgBrIMby9Fr2SmV2D3K7flXksq8LPBTPTdHtQapgHS
uqzUHAMyR7vtgB2itnZGGRO+Vo9vYN/QvfYWELpze78FMe7iE0pqAmKS00RXJpUC
Z6Arb/psYbFB35Y/2+0EaLuz9SDM9MgfzB/cvnHk3JyRNKobu03ne40klGddfQom
cJ/zVoAwpvMtFybf2ZVbDOGVBXiyb098q6LWELzwNfkDqqbBY3yCJUBDP+H/LwUJ
d2rhOIeYA1lC5ygzCc2zBu1vquyhMTV0Gq6MQc2HGD3yXepl+zGeyPBrf46V9p4J
To5IL+82Wua5u6FqXJd/26EJvI9Km4kyZdKzXeHD15l6M+YXlnFv7N1udSz5IfxE
DCQ/PwXU2pKHhIvH9xAGjO9VamYEMOze1m2gRf2c8b596POFzj8tOZSgwC2smJbu
dIyi20bKNSsDjyiQZ/yOYWTTM1KW7raGuUHUZ5/iSZ9eWKXgL1z9JomQeRkOUvBp
0ZnbRS5vgYrUC9ycC9FzbySsdW/pxMJqRY/hLz/pLu4An+Bs8QVnDuoqggs/UmTA
mW6e5tAJWM7xHMWSLpenxFFkUFcv6WRxoA7mUqaL6HlCAg8dtj5Kbx1m1noVzE6I
tM3bxAAI/U6GeeDcuSprLYYZzxjwZICz6Iu1PISiKv6iNv+VH0Jpc1tKC3qytzd2
c9/1BfN6Ro2c4k/PG21c4dVNTrBN4BFFHE6oO5D2NLHULK0s/khN8nTpE/QYL0YP
TuDpYNKsa/hQHSQohN7UsH+OrOudEZzxXUFsvB3cpYLP8bLC/2iwtsi+IHXh7Z6K
Mu5QSl00nK5APRYkor18u4Av9Ilq+mUzeecSSkM9QO17vONP9nIOXlyHGcg2/vVg
EOcozEJFUTGDbNIwSaX8uAQiyX2n0Q3FJeIXVPn0915ge3VGglBhi/ZinY+7GdqP
cdkHrnpmXYmQLjWI3strfWG/9FPwRF85IpC7U1vb/2DEZ8WKyR7tnrZFDd1mNHMA
pfpImwYgo+N6ijlACcahTodKj11x/VVx3+AryKou0d0ofT6FZlx5460HGqgMQIiZ
MxiK9bR7/F0inu/E6gGT7jEofEgV4D+P9cGn9mbPJHm5+zIs3J3jh0AhqZMTyy0U
krJydzvBKIyw8+5TBRVDS68eaG40TXW8O8lj+5xbVH1mg7+cwsr0wwRT6JcTkE0g
7oQ8JVV4YfntaafLAbu6gzTB+r3wStGRU2TjF4f5Z4BmSb5Q1Y2sCNGGDqHxnrfq
xyXvOU9dD4VQEiaLj3Oaelz9GTGtyNC27nXHAba72+COPjloJvMyS9sDKw7xJBNx
lTftlhvkMILnddqf0+pSdHzqaL+S/2cxO0gbqbYczSGX28ft+DGzU1NhDStq8m5S
4vM48srlluo+egn5QMstb+3MAFnCMUhF3dUHcEkem11rDbYxiVG/Xts/fmEVSkwV
fdA+PWNaDZrh3mj4Yi8SeEei/+GaFTMiW8CkMkdPuHv/kcD5EVeI9AGhjaFkAVrU
Uh7wC0liO1+2gJPss1FhOS2N3yBtmAW/mj68EwRgprHUc/K4qmgrTAvj3ylpe0b9
4M2dGNpBSTJetTHE5NO1C7uHx63r8ylJS7STDPK9DAuEMPFzn9N7W5YQIohn1Me4
6XkRmDQdVxQ0oybLN6Qy58N3adPGwysy07LR8nhKVVHyd7Zsrq8YGI8jh5DEZcvt
/ZIRyzblB4kksZ/PUk4YJ+YX0+ZI5Je2LQkCw1AUankz+O7YcEWGZnUP4V5e0O6f
hJNBhycYmiQoFJKp0L4+NUukWD8UPH6In/J2MaN+FzNXIh5zgT7WEJLWAeriFeBM
LtpqsV3dGAz4NLSzwx9lTeKUEZj6QHXl9fIEKRE4UqeQ0K0UFbbDb5h+iUOn7jKp
CqmXsLKbA4FbEiWGyXGkfc1lXFyqiIuD4upbmBTYZGsCjphsSF0PC9G8i7XgfOuj
povt6r7J0p0Dsy00nc/9kFr9pFZ6AA9PInD5hbI46S3BwwRCldEc3T3lpXsePwGy
8+5BhBLxJE3kSB9OXiNHDkxwL/ltvcX0iSHvPFM3PXK6eXzXFBSusPulJlP7OQLa
MMghi2YHErlad4owV8/0A4OfTPTQEFTeKo6wn5qPtWSzqrkyCsR81CERII48k0YC
X54RDd53/nFbgLmdK92aayrnVUx9M9H9cLgrk054BQqHJrGgnAyQMclrmIFGpezj
PAe1B7VI+vVAGZI+DnyFrrSGJ8pSK7ysZkWobNy4OKSRlgmcrnv/R6KkqolKP/4l
CbNqwPyTzOuWyrdFnAHyQhUiqJFHG0++xFfQSNYsbq8q3rusmTGgsNXsR4US6PjH
Z6evaRRV3Gv+TGlRzh4Ccjd3CeyZ0vk/sqNciBgQSNlpQ5Y6vvHabZAAjRC4YPj1
dt9yBfFDzsjhWFwME13Kxoth64pkJBEAN+q48EB/+54wB5ktJ+mCTZn/cVgfg0Bv
kX8MGhhZeI29Hk9kIMbO3TfW6Hxs6DJHF43E3mL5Stzil/BZjPfviUVMvJwVHUII
6+xCsTiC/dPBE1LMPL1gur5OUCZIwpcaneoTJHuH+7XCo9eyG8fUwghOByg5L8Xp
8zc8gQnYCNlqQxlZVkWb4Y4G7+odAyIZI3U7yrDD9q3n8HYL7ppb9cYhIMJ9vdm9
GfqCKMstS5Z1rxal2zzlBern7WrbmYu/Lj2lgzPjqMp/8IZGJP6L9kesNVFv5VgB
YyM7t0ajQWV9fbRj7lZv5L3dbkYpMPHZCFfok9vuc2ziooVPgJw7EeLATkG1AhNP
rR1gdSp8DisVI2hX+1SPzNj0/ZFGBuE0NMXmZNRh0ADLdooeWik4F3QikMsk2cYs
ZLS4eZWe+80VrqajZqy9Mw9VSLTU3N/P6ELn/NsCDFSVc8Mnq9oRhRgnXTwMhEuq
rtgKpiCElqK7aQBX1oEV+KsSWTWB1CoYW7RmVkCB/bbwz0EnuMfJfqencR+r5O8y
m/N5BxoXIOZdYp1BrbTBknGbdiCBfsSOgbZQlEsUVqSgUHbvZc9AezPVUW3Hnc2v
Jn2d83bkaxlM02gyzjaqs33tFKLsMpUrRGUBIMeUKkb37k04PgPo8M9NlwPip1h3
McvCJycOwE3/GUDlvfR9aK19DAFMdlsEwBzmZtrCe83+WI5s+fJB24RJbv65VZV6
PKvkxTJdGAqHK0XO6BBGOEYoJ7c4BrdfFAgXqMtx/NVZKKd6/k+eIYvDnZJNdKOg
B+GU4OykZ9rkqwx/MRL89oveu8OjJlF5qyhDChQwr/+SqEKp3ioNnBZ2xz117dMB
k+BgJQN4GjxBLM1Bo/tJV1eE+PILVjl735Aq4bo0Kvk+GF5Xkj+Cg2XNJiBqCEbh
5B1dngZATLRnIIk1g2dwouFO2zsHorqvdBuY71EKnnu9l2RZFwhR46BCxNcGKp5f
lr84c5dEj12ul5ceXO/5/q4z/B05zDOvX6Oh4CnfvgpDnu1t5zUlNAhYNX1+8Yhr
gWVszj8KPK7ojUkXd0XNoGcOpaJpERlgK1vrrgP5loTh7Ffu0/9F7pHB3HB//Rp+
xweCMHB56yqUTpimyuswyYJxF/U0eBPGrbOCs9ryueabDKpOiFi+ZijeQN8tEIjz
ug7m/nGPc+Omq5BFnAUmmWHHds5Opw1+epWiUtTOxGAkMhbp8FrVCYZVswjKbVbb
j+LIuuBMmbRH3qmAakw88K8VXhjoH7R8+o3cXZGM0VHKuvZhEKKZ8Qlz+iu4lXAh
dyV5Lj04oJvd8pPeQbx992YlGW132wgAADh88Yy0CPCKvA15GIZnOXl6YRmqf8m1
XjgKW0wnLfjLC5Q29lxtggwHRz9P67hH24N+Rm2QmrDWcvZJRVmGgPWbufwp4ca8
W6uc8jG9ukPLkHF2cbAx0mRgkum55TLTD5RnD8t2R8yzk79cFhqFVXyQ3dalI1qV
X4TBa3R1J6gBHlzKs4sPaNyIesD0zQHJStq8O9KJhmrgztzx+f8S0tsa/TEyKTQd
NhWvusn8a+mCr0MKtWOtgWryW/9xJs3qmurRHba0ZnSzLUf0L8vJ9i7brBZoVf3H
+UgbngxxEEuvOZRBKESvdIW17pOZGqq7I37yvUYJstufGxd575GVmunyq7pCiTen
SsnwH6dbPNT5JXxovfLAuBT3bSNUkx7ZEtH+DsmoCovCmrOLmMTpBj+gG7sz8u8Q
U0hM1iCu2+Ng8fBcTeibaqp1JcDOotqQPHv55lWe0l+Vvrq+hNPwxMDCWQzvTo8E
qhz9iunugMOtLkm9/8Ap75oot+VrhN4hp//tiS8vde3lv1ajJNTL96dolnSQhEtC
0vydxvwgjU9cWTE9UejUEVZrWb+aWVjeI6EBRzGi3UzejcmGXy//E+SdBRPVJ/rN
7Drfo/hv4/vd/OEo/5AaHsuSnBfUpOJW8+FQmpPUIbbjL1i0G/geYRigQWO2uzhO
xJhgfT311DmcVK8Y8teF6zHNPR7vagFRE1MI23Wwz+r/Af5/58NNR6+Q2wzBqxkR
aODW/jKoBByvccCg4iKAB5US1T4hdrruqm/FHOfezV1gIN1Ik5UbdRKdeDuXaoUl
G2imH6voylb/v5q+w/M6CS34cwm7qqaRgTEkMZQ6LIqH4O8nLIezXbxFCl6tBF9d
ApykxSrlaowHX3uR8EnxiINQXCCHt39hA7UKiaYynMCgUirsHZpCE2iDPbn+1bYi
tgeMyehhfKcMboktavLUdKnOssaNX+qKrfIrY7xtEvrHxFxJuUFyjohFx1QczDss
TE6gRfOG5wmuF4j5RDqWLGDL/GhpvVakUDLMur1ZUFPovG0mKzEys9S8mPDnOdQx
mTUbtNM6RwX1VikkTYBss4RLtw3APaCvoXyaZhS/LP5OAGWBeIlkK7ijuhvZkhie
N4C1lZjW/9KkglCR5kLg9AIg2cdsnqeMRxsKCa5QkPgK0HONJ63Q3TyazDyXevzu
xDAzABfiHRSMVDW5cwTqxKE2rOaAms7OnlEBlhxTTtxyny7Q6oY3SJr7hZqVk6jr
NwD2VZVYE+bQGqQzl+lxnVAFzXfBFFWOpoIMViy25q3LGurQ0+8cNNFKNS0HYWNg
iDv79LkXchTVIP/fjLg+U9Uu8kMURL9DlAPeSoCzoCTIdPsfEAY3y3PJimYAKmT5
befjA6FUDfDGXHnsOepenJD+ePwoWgtEmUY0wgn1pOFxUyB4ZiC4OZYIcSQm8pDC
xBLIuxu2t0MUYPHGfqe4HffrLgQURUoi7xAITM/8pTBIov/gaXjGfJlNTzGVEsNe
4j2NnI7YLz1MBn7Woz/Y8jAnFpTnr8JMTS5UDYZusDSOMnqKQ2msw5h8+5e910R6
1bI+Yljm1imZO2uFOUPXHGKVnCdqAuyBETBlOcC0zbU6DH9RMKKnV8fmFm0LGza5
P4UT7sPalrFhEMMu1GRCQ2CWizHKtjR2+Kvg8p4biI0OaBEG7xvNUAw5tojvxZfK
bHTMyzVOseGyMRLK48NPIOSwHlzxGQ8kns3wUr2rCIcs7X9lKhA9zVY3foFZKwsR
KKUqmYIo3MEp2hLJmw33aYWTAwHZhBbXJzu60kMb6RDM53Yy4m1KgLKDZKBWl4kE
ZGq/RDEzc+FvtRaCK34Z9D15SfM5q9Oeu9Aa0i/mzEWrT68M8d1XVm41kvS6LkVo
SZ75kp7yPj+jwE7178BwsJkrlzkbb8aCF+cimxdYjjVUSo2IyApG7FE339TNS6z1
WTXZ7qqgAUBvbFlXZ3IaOy0exOHltouocCpiKjZ2bDHl1atBfOoDFsJNoWx7CkFQ
PWAvhUnrbb09JgDixLaN0EyOKg39Bf0HqPpRQIuSvma+sCwv6KX5Lkwx3VRizKCg
PvEbldvjBoZo908mXkSzN5Uh9LEunsD+oxHPltzrFAEj0Vj/bz6J58gUF71EcqwM
gs/nLVzXjZWfYOjpW2kjaIlRNtWpuqmijg0sy0QNWGos9TiQ4mV9Y1vOkFh4pI9I
sUZv++CE5OKnK36N6UKNNufXVWWJxPWAo2uckcAqdnqbX5VZQeQvnKFCZOtB7WMi
xfG8I14h/qaT07IBi5pnKMARRxWw2YmX3wLlQnx6kFiSopPTceRvNX7cFYeY42ZF
LjRCWyHzU4VpJnBjnT8y/a8eA46tXd6UaiI+yNxpDnmKsRBqcXTMmsJ3qdVWSEsT
91Pqh1H8/S9O5/bfrPvziyBESO2gN5viALsjM6IFiX3gE+3zybEI7soOSIGmriFt
44P4AeitvBuCo3NWtBf7Bg/MtlfBZZCkeNfQ8kse/+9xFoLwccvNy9OopwuOktMt
Pmmm4gZsZGD1zSeUyFpE1+e2Mp7/xPKGc2YQhbrvt3Y9T4iGcFEvQY9YDEmiO5Y2
kxRrscbqvySg3Ku8X6flxtmn2T0VL1xXeh6SBQGDy3zPUxSYWbZBwQspFPyjTM4k
snlFZL0nACdByTc45HivQJsuDE1KJv6bECLVzi2lPs8DjBJExLLB6oY1L84GO6L7
LOH79mFGLzMtE09VL7h6jFtcxe0pGkZUKhZu04QfnuRr3RuOFS/etQzvY+85CBJ1
t5+lzJAoL4bmXNHcMFVd5XOry0nLCNhg23eJgN6ygzWsTs5hxasSEq3H8u+1qO2Y
Z5WwJNcow0P7PLX4bbC2arRzO1jwIIFsY92iyhVNB9FdCyPqcsQZ+ZsRLOgLCshr
GdImtnkKpioj/FBVVOnCXLjYcH+HMywQtCfxlU0z6r6qSqJfbnDEw71mHq7FArNJ
vomSBJhmy136+EpqV7rae0PEVP6iMgutaIbL3nPxc8p7ickqH4XiCpYuolf1Ln8j
v1QYmdWpe0IGlNeah1WjOV9u8ZcBQQTF0xiEU7/J/gNrBLqeeJB4+rrGeMiksHpN
3ypvq8gnajgfliRAth3AZsJd6kQBQDu6GrUhl2W2RrxbKDASGv2+BaG0nmgsFVOl
L22yUT5rbg2JUrbn7ELd62Qy6i2qfGSulG0bmjKHR6YueAmwjbkASkh02EZL6Bdh
MhkyDdCrPBtyzbVxK0NqD+s8SxlMj9gqdfbNDijuuaXWc4q+f/PkdrTlvxNELrV9
coPP2TJCT9vVJhWqX2cH6OpIterCTSwe49bNgP/jzfkAvdFsz1fyBwT8Qk6QNur4
swVhifhKo65Qx3d0t0vEwJondewwNg4e0BfEGH2nh4fkLE+EXFXry4g4/Qx/CkQS
CBThLUqtJN+1iYlDXeI3jYFzmj3v2CKtIu+WaPC9ekzzwvXSz616qkKugGMaQEj1
8sUmzs/KwcstTe+zb/8EpIzkcOxKUcfiPVQBDoLADr+/qKg5P3jhxmjOjhK62ryl
aRZtloOl5BXSpqr5Q3A4Zk/QGGX5pxEXzII5DJY/UjPAFMztF2VZlEdRjwbloD2R
XTSprkpKdLygpst0oAhVgQc3MI2LsUULBgwJPh6aQyJ4/lOJnHnL4RuKb62zy3BW
1iiNl4qvJ4fLHoSLXIECVKzUBgPMfRquSKrSezwIv2QDOYK57/WEhZqcIT1zdViG
R0jyHUdFhn8z9xxOCTOGWwkiecqmopqFixWoqI2MoAA0aoLjkw3o08aUXDuSSan1
Ey/H2anoWXrdv8V523mYq5tKD5NH4mGUYdgBU7j5XBkw+lz0wGSVnRy5/SfdFS2G
H/pM91hQ29oLHdjxRIb2AsGRxKhCYiE/eAZsul+4hun3DHRFublIpwdrPQfnS+oi
kE7eS66VdBdo6fSwmkbpj/2YJU9j9irf+xYJh57tENyS9n5QttRn1CN3gfuRQCQ5
CvVmneUKynUMRcNgGk9DJfeaih7PsTWaYJOxbGERoBXGV2wKDhzjLlf5dbolG1JN
4bxq0qhxRRBl02zuDxqokw+5zGKCoGOBPN7p9d0Flq4iHrEGBuwVDvRi/T1OC/ZI
IWE4O2vmma+gHD7hsxD3X/7RfWU5pgGavxFx3AqvkRz3AhFzbp2luk1veFYuNe/t
1irzGBUR3++dqYLylPgN5cEcICGrXm91MZnGsJybkM3Tu/WOIwGLSj+hxNVfmkye
KyeaVm3gF7DjazUPYLoy8E1M2wp37/kS8gNZ7H+pU2aJ9imd1h9J5EonBMvKlgtt
eo2TYEwNfoyeTVpkTwTY3mva0bUt2obW/3m8XWSy1SIm/RbkoerIh9ohZ2lnEGAs
h21EPfPjGm7PPm+FoE2mA92GYYeoaf1FSK8GpoIJx2RaCfbmk9iAZC6p4aiQXSzH
9RENrh+V/4dNGb7cD341a41l4nbt05SSNpqxE4qdw/IEVaVoWf8Twm2v6iCxiMpG
`pragma protect end_protected
