// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aE1uie7Z2HxAwOM7ma1TPVy6D/gJS51CPwZ2Mu06l4Ci8D5yyKhaRPzY10bGDL6C
wsDTzAASciDPppRKV2BLEsc8z4iR1Y7JAZQHZcI1wb8ffYFoPalcBQJ5FZsRitMS
bRXdycPFiyKQ6D+eKFnuy/4RslonVzcV3IzuuYFjwCw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33248)
dyEOPmZ/5utIE/n+6l1uZkPSx9++pi4xoH4yf3zqO4kpgfEU7AG4FyERZ5y83qYS
oPzlMdwsJ7iBxtdozYdMi41Z5iH3p7PnZyJUa9Yue/5IlJUuSojBFS7C5v+s9uan
UWILUaTci3dr1oPZmXrKVpKvK0t8EAa/t7e1r56et6o5QbWWScURQT9v/OXAMnZW
Kqwyp+46mPd7C3EO58q4BcXEwNrmevFubtf3f6NZz6aX0Ivb00DG+vNmlNle0OM1
lTCXdirRRgThJgdcF+LfYG6q9TcYusich69EBRY+5uuvq2Zrb1HbmFABbI3I1i1C
37FR9Wa0I5TznPuTr3EtEGaVbVp1BvZjnH0c4qDVthMP91dg8iNbQwzQZ7DBmrZ7
4EYuBO/8z80OJuQNmywCkI8WqqSt8Qmftwe/aBCKfJj1q9NjGVW5Cp4Ey+viTjQ8
ilBRjW0UQSg4SHqlLHw9cpKel9Yk3Ono5ZR6DezALE6tPTQQMJ6y13scCai7hjhS
UwfluW8+vG5pobUmEUySRxWc5E/NjvaK3MBfEuzRuEe10YdXSZ1azALDYNt8SZWt
qvT/X1SYroZDfEkvYtupo/k1UZTPGEYHu/TBDZHd4hs2I56LF+ZC6JUWsYEad5BR
4QSnnbrTI2Y6p0RTbjYiD8bcl8lAX521u4XJZWGodO0qA7ukcHi5V36ajn/lK3mU
uWp2PMC0ZUEnQEdrrmukPkCvGN1feGP8ld5z15dQSDR5IbGv1ZYXdzOsFd5W533A
TsVzTPy8xsMe/Yx4/+BK+Z68s4nyzsqNUxFXo5Z0zZRaJCjKSpYyib6rQy7FAX8L
FYFzfREItgu8tLlUYWLC5bIuG/gL7hMvi52cTY7E+ntEW3Ohevs1Nfsel3QRhuTQ
PDr6smene1Cs4IFucGNT1xYBHP2CD/7PX14I0ZxVOGpTa53txiOKg7E4EO5dYtud
a5wRCq1RcoxmXKUfZFbWj4UgNvI9W1S6hW9aAm7DTJIyLHbK3SqLfXmBNpSNNqlS
w9lAH95D68/NcaaiQxf71dAOh3OUMPKIaMCSpeg/GfarGrxO3TzBUViNU4jhAbva
f82+uLvfUFcUFB1tHgXdR3SZn8U0KIdjf67O+LCTvDL5wOHXnxaChBF4kU7h9Z3G
GC0wqkHNRVGN6T3Hy8n3LLA28LoDN9r5hkjdmaYmwWTbCgckq1w+3ziS5SYrhmIR
4sj+ze5bRk4BDXuFxMsYy4F1Ith93yJTrT9g4KRvKN9XWisPTVIFgqyvBvjuJq/A
Z26cXLqP+NCbyIEO23FYnbVIUyIBEz/ZQE0hFNpfvdGVVCCVfdSn4Hv490cdlgwh
KIOiMp17zfthyX1OAm/AOVFA9Hrq/Qhb8Yvd2u8rDj3Y3x9jrf1p1iJSo2L1YTul
hj5952oVwRQtzzg2dqX+8stcKH2sOPDbTj9jOJSXMw83JG3ZC4FxblR6YLdwDzQs
3U1bX3oz6pwWDa+uIyD00ihHtSSYCHQbS4R47cY8+cJV0D7ueSSKvpOmjE6EFYWW
AznRcBhO1o5xo3JEexm736T05lkvBmGO5SJgSxSnqRedt8c0kM+BVEtqXuDseqyH
LCHDv1NvGQnYmDC/5nWVLvXxDdHVOyV1f8CtgMYgisV4Iwsfn9aL4JsCV1tFYBwr
B5GNxn+qO2wBWoX6FbP+BfVGtvJ70hr7TWt6sB+/EnjoWq69S+0fcB8GaM0G7B2m
lpjgRXdRY7E9pdaiTpzpTwXSqXxoB4lmFlTAyL7bcQdjTnfR3R2igVRWa/YYjaAH
0kDnaWdLFTMvP2kVUBWy3NvfO/YusvMnuDVLx5syifGSCnyMSgUH2qo1uPTviuUM
ITtd77nx+xCB7SmDDAsJTzxiuTLBUx0icmbTEbdmDJ4YIoAzMkKijrE8TUWpH1rb
CLHJzvraGkVTJjqfvbpiOihc2p9EQ39JsXzCVCOs1nvWPfOn6tfYB+L3CvSYVK0X
Sw9lRYr0WaASEoQfxlLrr0BWjbS/llShBtB5kqaxyWsUZKyKvzu5xTYJtsfsBMY5
OBNIXtj540Jq87ushviHJAEzuYbcf3OYQkRhbnhVDbCQgwFapbgg0hYrYRauLyJz
41cD90KvSZQCVUgiU8luy9kTkWmYhXCeNfKp5MjweXC2BS9m4F3d86uk+9IGn1UP
Y3gc18htcIEd63n9IBS49WCVrnjTCiVQBwgCWSljAxXLCOTTsVGrrLQ1N4/TVwEq
s4E/6WVnfQ1RkuFaPbM/c15w8lE4rzz4CuPZnpnP1b0+aXCBFBMb+Ra6gqV2/IXg
XlcVSc6H95SPVbQlaBuPz8CPsNQl1Jd+snlCu3E36g+Nsp8F+maPAT2aj1JpB2Wa
f+UhaVl1O5SYBNvvNFyHB1QqajLVha/beP+XgEytmqZzi1zACrZQWeYgiB2zwrou
D8C0AUJ1dNSiGOEFv4x26M+Z3pblifUDMGzIpb/H9KKr80bZ2T9OGXPUY5OfmbXT
MclEWkuSgbax2UN+WI1XEh6xJGyIDsWJPdrWk/AGfU9vJuFZQCifDDrUZX/ytKCy
ibFyuXu+2NAbqWNrJhybz5O5o1/WFPZLy4uGu8OapdRSL5OWG/2WGiKp9KZJE1+0
m6BD2PKLxIIL8HRazOb5W53VThwJMTcF8BFg1Mk1QNPonteO6dn8uUjChUDzrKjO
oAkaG9iHeDrbZWlmtbcHugLpDCgQysVS60JDaVm18IJNMhlWrvGJVdoUZUjpxAn+
lRFUGbJq5YetJC728htkUVKtjHqCiaJPoYorKUHqv2vAahiBDRJrbFxsqUsDk2Yh
npBCaKPRbHVPNJ5iFG38AmbBiwTPapdHgK4CBPaaVukKaXBterEgJkqL/+FTP2Fw
S8UicpiSKIsvxrasNqyrDSdbR6ZwQp5GmEWY3Xx6fKRiU0tXZ0H6PGpbsoLmQNHb
2nH/Pk6RvOxLuMs32HdRoGvcSY2Pmx+1eKooTUrmP1NX0oLbAS/xEZ28SVFZRYRf
TdmMHoe7CeVZ8sEj4RIZKazjypxbTa/XduElwunKDRxKHHJhDYBwPDk97o48yvTS
HtRRIoR6sPydMLoTaccUJH2hgFt73XaznZH/Bjg4/4BCELFgePapks4Xl328Xrcr
XAK7k51cKEIgItUL4jQpOe6stju8Kw5BmY/9/1cZklX7m2jthZQr7GHmdkGpogC5
plrbaVMrX9AADYNFageyMCFgJ2DRmJdEkNFHSqwzin6HzHLg3Oez9vTpbCJEZvWM
UGXFAFtDZCEr4TGGo8njhvOaveTVi12odEQG4q+rnPwCdqmdzlY5BP1ZNYEJrFv0
wM4Wc5gjWn5H8lw7C4fKe3Hj3IMDRkEKDc0ZjvVAsQqelOPS+PlkDRHiqiseuLBf
KZdv63cncMjktfWbKftVJPJ8AP3mUzUUi0tAlNQrMpCd1h9x7oGmmPw47CPdRy9C
Se79clBcV9MamzW0mUYV8RftsltRJ3zE9ECTkANLW15umb7foc08K63SU0nazjgh
xKsReNrflefK+uqVH2KP5OsKfzz0q7c/GbtIBCC4PxGbK/r2msVMpiTcml7rwPWK
UbiO+94JI8/Mu4CSh7vklIn4FLLIxVNpKy9ehBMacfcuuThrVd04ndlmrRUYDhVC
8VkC42CZ+ktHu2Wa41oz41Ot6/1/N95ZvSNKcfFmzadbOV2EHM3AvznN9ixlR5xt
jxMrzgmFSZ+CRxUmukMP33NIWhKlV9FO1PqRD89DCiszPDKklMH+g64Mla1EA0gd
JPtnS2WqL8wH0FigNLiDBHhUeOrc3hQWpS7s6HAoNrNIUi9YPAZdn0O4VRGWZixH
rQxlm0hIppaSOQ8LKHEllM/k/HI23c52al63nfnUniXHfjqHPmTTThbiXHFaaTow
yLW+/o2IuYC+J6gnq4wxBu1sHfpGZ0IV05bWvEfsqQcDGDT8posIyebS96KXxOt/
aaarXns1wZxUw/8CYrL5ir3xJLkBYfaZ/L9iu1dVd8QoZB1ad4b4MxivqoZhVkwG
YBOVedNOy1yh8NZFhJTmlwdvkeIWQUJpKZp8ros3TIVfZrKTt+UxBtnqJ7YKA5Ov
hudB7AB0sI30yWlv26G6IhUdoS4/f26ig8UPV6WAQ6duWGuC0YvYDkL8momIGtRh
znnPu/eMgImr7tp6xsrhuL/E13lpnHfVFumvIPK/4bdMzFNLMJYTfZ7/TXv8CqVr
NICTvkzMehd9Xk1S664ilTg4W+ZzkXWUAKyUhkxo1kmZxf1ExtwAiXmLKtRfkKEA
yRLBZsO3tTvlWNM3zJe8D1CiGomlkQ587/1e2L8CWi4uYa8xGXOs50GXNtv7MqR5
7LTYxOKTj5IcdPYaG8U8M0ON5o7qqhmN1jdAgsbUfn5h9XThABLIAcgPi+oBwFRu
LBdhKllE4A4F8ojZWD1M3PWd/tfZ5Cd9PX0F/9S1Y8LeheLxQnGc68rOi+/uQ/YK
mmobplhmRmPxuFVXWC9uA3S6W3uYecGFmP3mdiDIsrQ1LxxAFm8dvLVkrlEXDVY4
l28gMJvzOxW3obTEFGtRPX+8kSkzZj5ynVB2iS78CGyCrod6HyydWyUi3KsOyC/B
YAsnVRM7YFpj+FRB0Qpq6hH94MB76EB9bo7MCh5vRbis60HDmYh/vNeigGd5tv2e
itIEv3jXrKz4la/IZA1TZ36WGvitYmHyOdl/EqsTILJfdu5NZMNgFDoF2N2bJ5we
P4GcUJoRL5HiAuPBiD6r1m2LGg2WGHNhXNRseuMB7Q49yLyMjbirnk9kTr8e5ViE
pye+KUr9CNSEiLBZRU6wGiR060aYuCIs8pf/eiUsOOVcwTxryzpovbjS7LNKrm3Q
th2m3JXASfmjz4IeWi7owAsg0mRebmjYbpZfor0SYnbBQh2vKD+nmcNK8CXCHW+r
Tb8FQaaYNhZIdNJM4CB8PS2zo4wIDwBarapjQKfwX13fSxgriqhN7/EZvdgOa23F
LdXSBuhmvbUYCsgtkOQe+cbAVBuZNfu8XernaOh17qncg9hIF3ooSUnseTbiUoYq
KAVK2PcXtSi5b+uhcbHDeQRDlc37JM4d4ivzIOi+3TLzORL2vUAHAq1fmSRAQrUv
ToBQD13MurccoWe1jZYI9NgKT2aysilI5re/8T6TV/8BDvZUrjXbD3rwfNWxde0e
zXJtO+noL4UdET4LPfyhIxcVqc4JxoiNE3m0VAz+lcs1i/W/hZORTkx41hSZ23hg
79oJcwKqlsucVqZZdZyCEMkAMBU5KlIkoOTWcrHlyw6ei17Okl/y/BEWBIYN0YeC
fwgwVgWhTlPzfopDzR6YLKVxwYHKMHBvJFtzs6LM1fPyyuIgrqZCz0gPV7/5RspH
9liw6NJLQACskUv75FK8P1sh8L4vXiaH6mnPr4WKmDyHbeyYNkxJeBcVTuvTqxqk
uFHcbxIvWPuXI0US3OBalMWloynhvmbeM3u2BbZ4Fp4hTmQCXO3ParBtIofL6V97
kIqA8PB7ZNUOMXhyoaRQccKiGONEESuI3H60gTnr7A0NB45kaPWcXdwV1vlv/bxj
i13Msx9UKW6VLH5hhrF1CIFVrkQAQMKjJP0PRkh2yovqpG1YVAQdj/atNQqMiw66
RNOQNveGlfqCldqMpLgfokHNkkzeSn0WQidr4ljpQ7Jc5iH05Z8GdqWwJjGeej1j
ie2R0FhgSGS6qLAouGV/gQw2hjKktG+sP/A0ydpmhVxI42Mw8vD3Ps/04AseKIAu
jFyb7NHeEiz5/6EXKqw9Jl7KShRFLualp3pfjnVySmXz66rVj24u7pUuqaFdyR+x
6ZvIVyIsFUGwAvsQbtKA4qgLPU4bO1lIteUPVRaoWwINFNNaEEht2OO92glaAuCq
1HApHVovODVXaT/9o1tkfDXBWo9/lnnCEME34pQ0zocDQhY/lm57hGRpyjTAOquf
Ag51ESA4Q3PT9TZdSay7bWezdtdJkUwnEq1DnnVXe+bqSMsqahvmzxooUdbIfCRl
sLc988oPdhd4zp+k/AsZXDNtzHAnTzrxT9EIYbaDM4tX3BJOgEQE2/u8FszYlvGK
QLt2AVbZmLGe+0eOiN2gLviyBenemq0Zo5y0sIi23S+blMYsKLHus3gg4wyQY6xw
7gt4N5eAZS41axb6ej0RGMxtiZUagPupUTS45zpE4tyLh9cFIP8BtugLQcXls3rd
ygLrSyMpQ81GC4YZscfzmJPgDY1sQ2mnDe0u4lU77FZB6qSLhgjQDM3EDSMC/R9d
Z1O35MKPVa7Xai3xdqp8nOOirFT8Z71oVH3mPnnUO59vADqHzLp1A4SIn0hvp52I
M1QvE7Rkr2tetE+LQs0pjeVBR+0eK1cDXV6X80FHIuxY/MopX3pvxtDXqS2YkdEx
a+qBlzdv60s1XsZytdSroLPk85h8JzE8ERUExd4nIKCqsxWAyjKyClwFAUgl8l+z
Dp6FeE5KR5NwiA5GWBgkSRvvkJmunoCQojZ1nMASwGYGfniYXzkReknF4BmObLpy
XW7utIOw3vxahztTVoSm2IC2rgLMT+3q/8+7HNXcbvaQtHqwcLqWNl3qQ0LbY3j+
fYAH6+uSwHVjz2dqc8JuYEP+9JtlfN+KtKrEGg4yI5cRq5+ugGawp8pW/9+wIrjl
hBZhVfJ1mh8e4EgZAEdKPpkbR5IqxaTUxTZROTBPfskcEinkYfpBNjnsvdPh7vHF
qq+CtVo6DGW5rSSv6Z+GFFgzKfeYMGBPU5KtgM67bWB6KvnseSlnne0AFWexgHQK
P3BNLk4T2fbJOOsr1lbpC4CI8PYb2tHBBOv9eJVyknxNCdzFa99e5kE8nQLKqN17
rLn01yiTo9ErEXqCH9wuBBt1CsW6YgJRLU3YOwGyGinaICFPegmBcklxLuY5+qGY
CoBEtSyZsnyMwPJ6/Zbw9Ytoxvwqj8lHQs41d12S5Q15TgCOqJJ1ZaxpRWDju8JJ
YZ8t/sgKEYSfSYofQ7HPqBCeaM4MsAcOMsLy4mw7NhiFpQ7VA0p29cuRq0e37IaI
MbzxloWwWbh2P8/7nO8nbNKHZN+uJFwUdhbrxDljPd2ZjVLsW0uAyXHnT+dHzeSK
yUhZC246aJ4pcbeivw93xGiYFF0X8nzpup9cNtbbZGgQp23tJmaZTqdhus5E2tOt
ZOWj+8wyLgHTy23Hm7htTvsMK5ybn9THT18owkY3qJEPEkXDiVkJA9c6J9G0rNNK
jRQGb3M+xVABq4h85xaVMx6SU9HH2qlr2SfuJkbdAm9VRIH5aOk0xkrMctk49mBG
xlAR3quAC4ofJiF6Mf254s6mTOTw2bTwyUsSan6f1Sn07Yeca3gnevI2I0YEbWMt
VtqUoOYEs2iPkfeqEBYcKd1ch0qJwsOVpuM9BKeDXH7C//DH/Zxzz0YB7sYznLMl
uat6O9Dl0rfBJUQOQ6bOLarsclKZdSXZYOZlHxqEiiMnBqOHPtOjJ4Y9Cy1iXEHc
B17pi/Yw/tMnxUJfuEP8d5yYJWuu2gbIYbSFLaySdkcf+ot/fbX2Y9+6qBdfZIFf
1XGLSSU303L8RQGltY3Qp1loWHWZ1n3aSOKQWoHgkuivSSegr0SwUjPXDQsaBNs9
LsvImN87UmSxoxRfCbsQruebdopfbWdqvEtVw24VKA/6dhz6ap9Mv1PqJDncyXzf
rs14ZIsSIR2wFQzfCwakv+E82vYW1XM6INzzy92tFGusbnkaR39syDZmGKbZ3URw
es/l8DlMhM8eBec+A4m6XpVTt5gWHyDIGRPuNHmburjXL6g4hTcmLH8apa4qv+AI
ZdMaa5nturEybZQ4VE2sPxz5asrIIs1PyWKyIEujv2c2bZD5gqqeHK40vbz+AQuV
J4MG8IRNKqDKcDGR6JhqzPa2FJA3gisTVSUNCNt4G7ZtgSUs53BOSrE4p7zptqtG
8sDGy9uWuspaFCSIDG1jvj18LNGDXmaIc+LpCbrB8/F70/eeiFWcHVDHCXdCtUN5
ISmUZQYlqc0DY9BYUTSHOs4VBCDPCCDn8Omu8u0hpKFiG4dC11NsxbewVQZkN7M9
8UTUCdNLyyGkTIAp2p0fFJNu6osRiFwaIXku/4z0V7z5b+Y9KEnIpEQIWRIQIk/8
18i7QKj/HVOkeHbMmntt0eQCvS/EdC5p+jns0dzOxFbKh74HUr2cyfrvNfH9xO6p
3Qlpy/WSXBSwt5gTfz9lQIQ2PP2mrGPjEWod3/zAKvWVBBYzg8gIG+Xq1c9XTCXL
35TaW4LeKavqRgJOaFWReXEKHfnYIn7EnK1Cti17l8rPVUZRnvtzw2RcYbKW4DpC
q/MK9tfjcrDQ33VOTdpI+ZSzxETR6sE1nAHF87hweOuwr2sy3fH0PS7cGK/FI8E6
H3Uoc/RLQ2MHo2GzYHpvlw4F2t1X3t7yxZoqLMt8kSQoSUXQktalOTNV+MebGwiV
4OkqWvuJ0GUX3pCHRzDqJz9iEBAcnmm6AH7dQqTUUeivegV3XGgzFIxbZ7z3HSQq
ILYpRy8HToCkhLm6PLKaq8fNqZ+yd81qyCa9GpTLFgFpk8b1MQVUrViOccnyo3p4
Lobrl+PpeXoJjOrR1XM8GIDUZi5gwHiz74GrKqTrLAyLmr3bUCElCPUSQp62PBbG
qXH46UABzQegI7tqRKo2UFDP0wl3iRa1T0jAWP1FlnU5f/JJdiTCCUEP2EO+0k0J
dpvf0gej4h59zOG8UtoeyL3Q9B7SUv8axVipwowmOxIi8Hy0aUobbRCCt+t9ea/q
lacKtmQ+4pgDvSK/OgJIZBLCrlxnpcxSP5eQ0y2riJ3illDWNFun7/k/kYHYyr+e
8eqzbNv4Q1bauK/oYxPKxiZTzioSdGRtydwpBM5HY81DFmZFUEB/zIP66uwbdRD9
aZgY/zJWHyHhVaMRY/TLKdFBf20oL3v3vf3Du+W1PVUF6ao4a6yLN2XFfw7BXqpq
WyOPcDtNoK+qDiIf9ec/06unTCsj778uKW/1SbJVmYEILrMhWFDVYCDKNdRcvIlZ
QlnLkNtAuHiJ8A9LxuwfoWGIo9hn7UfFqlcC4A9FOb9IoUV8XKE/SWWAs0muKbVs
icqm0E5aGXdAsU5jf4SPdYebMjE49/DVaHPFnpb9/pvJwr5Mn9cnNeYnBx3GSSrZ
Q66ppOGC6cm5k7ngLP6DCf+tpF+7q1VMlDT76oXwrqSUqVEx/adnrU3HdPiIJvGK
4QVSndtg/imqgob2Z3lHbNe0VtLqs8Y95ej9D36W0pn8aImHzBTpsIXDGU7iGGtn
UQIaTrb7iPNLzuombISEsrTbR+GvzJj0eJkdgw1K1IwRL9FaLysjYsP9eJ1ZcK26
31vVMfN118p3kmRnT+qOCyMKruB8smImua9F4TgqLBcZcQt0sbsnApv6xambCz6e
QwG9EVcin9amWIRURyy44UVFpXuWnkkoJzEN4x+RMfcuivTiA0mUzUocOlRuiRUO
EvjJfsW1qQ0/ZuGl79nzMVp5QwNyyxysr0eGbBybgWgmmaMDWSQwBzIeLH5BMf2I
6bCAwGPahH59I3gHnnU8JrWEr09ZeHpdT/rHpwfSolf1fSOLTuhBX0L+eGjml3UC
GCJQ3HB1+Ysl8K91n52Eu6G3/nADCJLaqPRMD6cpgLTOJq/Wxn1yec9CDjQFR3xc
fZHDr+KnqDJzSbTvINm6KM4KfcAsmrSABuFVECTZzsT0b3tG8NMs37m5tE8E9756
8sSA/mSfkFK24bSDi6Z8YeUOOLWxfevfRnmwTw2WJWsiiZqA5UVRoduRMXKWxgmN
UQAxti2C02WfTjVqkoBZco2+cMsDdU8Z/sOabvJzuCqRBOmtDHGsu1Fi2ZZODyiH
asJZfG+KLvQDEbArf42RqsQnqVNvBgxTji/JZ7L5taIxgE12a9MLFIKJG+Bdu+0u
kGbwk99C2r06iiX49TA963LMQ8IRH+t9qtytJtkkIHvOHX32yjLO1NO55UZzDpc0
CD3/kcSJTRtpC/kH+GnYhYhp/vSltjF6hSn1KNIMYeje+CKaQCETibG8/zSOza3U
uSxc76HPJyMmRXIXicaCaaJ4rH9XeZsFJMz0njTke+lX/Mzvjh3EHhKZm6nOeeKU
fbwwXplgfJWtA7GaXhUGqrQE3I3R90tEAYC/lSGL59XU91tOSNKP9Iy1QSh4/L8q
odd0HCNVPcVB05v2uv8hGbM0pK3LrZSn+j7oTwidn7bFaJ9IpD23hIUzPUuYx5lK
BvJDcxdM8V5JDnawQDnxtG1zO5c5yTS93AfvzXbeixxHPfGcq7SeBmZj9C8WjgHh
z7obxT1D/qL6DeiXpZ27gKWgc7dbqJw4WHL6fH09fHs+6kXCEF31WVdkfntRAfSS
4IqBOpowYJtvEu0TC0Us96jHRGDPsJcTzqBxFRVx2uaqDci0y/9FDC7uJfOs6jvl
mB2ZLc/VEqzsMdVw+sKeRU9qBuhEvXUnfd3GP3BBjXoeC+jSacGouhVdALE8rDFi
tMyAUdSu+3OSqOA6iRmvBV2cvm0Gu7QUEBIk1E6JGJmFLnxweVhBNdF152+8eoe7
EnLkr1Lqqym/l6g2XoXCaHh2kSOsJNqGnrm/X9gys5QG3RlCUcrMA1Hvqm+gnQ6u
E/BD8Px0LfeQPTDxFfM1lM2EBNjrvJWMyGq16x0hTbz+ITp9D2/0uKPPQkzxG77c
zvQImX24jQqtIfgWdsUDfM7EhsFx/3u2D7iJgEppshd8326D7GNthy686dnuUPli
QgI1dJj77u4Gim3Sh+7ypLJAZNLqXQUF1ZEI6XN1xaeb5hyoiFcgl2napkephlZ1
i94ItXT/lDtJCgCtZ0geIiqeyd2EFRj1x4pbPG/Vo0CM6JeqZLPMQQfcNaeMy+oC
VWg9EwI9NAjvEv9uB+lcMcIbzR6yd1sqE/9Np9lX0bYMHFuxKoSaYv6dn+KgaAua
34vn/kc6yNz92FdGfy/rKNIBd2pv9jSvAWB3gUt7Tr/3H3AVgiRYEmPLejFlW7lD
Xme0jGTXHNk5E3usw0z0pmVsf9nocAtax2bbKkiA04vGC2UfGVg7Kn/EgV8ByGzf
+Fhn/Kiz+gwkpkaOr2WQXkuBScBI9QjgYtDTLuuW6hjsAWcygwqvwNj3EfWAA+lW
0hi+mwwPuxc358fgjVwcBrhWAi8dflZJT+yvA3xJLmdPXW8p3m8//Tl7cJOcGfo7
jGeDJeEZ4/kleC/RMROYOCfqlq+Uta/qxs+n4kC013ZJlxOmRhpRdf4d9ar92fDW
U1onbOgmkltn29UeG0p+wF4OnhebFvJoR8XXgG04IdwSJADjPDWO8Jri4lB2IKJh
ZFwyY87z7cvY+rUyqY0cI341zBXl6qB9AVaYhy/l0mhuFc2R1U1F8uM6VWuBYyC1
c8ohfN/XTP+ljT6dNkha9UW/2DdX5WO+oaRxYy/fgN47Oh28oyKnsBq7fbLjLkoR
amprqZEdJ9z8Gzr4+CMzLwveWQHeuIl1X8q5yLJybGfevlrGENhlaAbNOSRaRK08
SE4kymcL78j4HwmujQWhv1Gqj6cw4kcV6ZdMz1y+6oDz3dRQmWTKDWWQj+RUKAI7
/x+vyJ2bZzjDAvy64EpAsRTFniT+U7G2/bLops5xzOzScYKpIPlYN50/N3aLjxll
zd0L3Q61oYhGlywTJGByyafWFgAcq6Jed7rRsY4H1eUZITNsn7pOD9uydaxrJK4b
C1rRKSroX/qlbGlAXmcnXY1vQriTUeM+aMYkCj97ff8Ze+tGhVVINmdo80HbDXuV
KekmPkV7zNUnsFJAr2WwRloL9h9jWjjIf/8M/GywF3V0awEpybXZ6ol9ctzpwti/
rXqaxv7QY+Iha0UhtkQPzhfT6vh1+hmM5s+KlwhGu0wuA0fgxOpED3Q05YRf0QYF
usRX2/WExWk6dODH0UTzv5QE6AAwvm1n32TsgfhJ5xxYLR9jXWCl9LEFes4I5S9w
SndSEDSq7OolmexCXkb+UHfEKtD6AdqC3CmpZyM84zLiUu+Ig6S9XfOMZxYfpym2
7NqylSj/EJbrd+bkeCmrmePfhHUMnVbUBrtWIEy/EyOSyJucGr0Scto+2aP33vmB
fxsEWeHZBN4e90kKzseOsLoOPGolEmV58U8FbfnSAB9Bzb3A5UNp1Gu4NSGjxK/1
uqUFBxKya13WbRKJfB8mN9xWfBGYMd6P/12ZnigRqULhLBvSR8l4NnyHQY79HITw
FswMNyU2FK50BvsVfSuytiPaV7zsKdJx0sHcfusQCLH5+0tt8f6NQW1mBzKLO8/F
YsBaxt+eEflDeMeooh/DROCGtsPK6HZVwQqFvS731smjQ+kJD/fbYkJuOXrGRfWp
junfpSP44gJY4Xjc5Qe8krhcCMG2fi2m3ZGn3OPX7d4SXs9A1lGoNc4wIYTeyd7P
eaPrIbctSiqnWm18XkUzx37s9MwB5cB1zxX/GZDe7BRk2rtbRGfwR89WFroPKk9a
4SDiyiZC/pcEwNPJEn7drml08X7ZboOgTLMSg9qQeybwIv8MtaXAAHPwWoVCBfxt
/QCwPB0/Lo6l9RYXFkgnbI56NA/jk0gmcK+h+j0KQgbET5sk8pqKvxZVyvUafZlL
pzVbzMKoXAM/gEPiYMWHq7j/lYtI9iVT32SqcwQcHHQhIX92sTWkgQLOQV6d0iwR
gMwX/cQe2Ke1f8Jpq9G7EKpc89gkmI8+ATGCakV9hKesim/Ck14O+Za27S3F92Gr
WdKvAN8GiqcGgp6CYwMP+ne88Bpn5jRjW7qJTPQLthRl1OEuPL0Gqc0XXD09kGc9
UjC1N1lSmSggF922ILYZJxAqoOow/rSGELA5Zsb6Dh1/HmsR9gHK74KUHmLMoBBm
BW+3Qizj6yMeT+6bH9Y38eUhzWvIn39xRxi93jM/8I4Jn0V1l76k09U1NTvDa7p+
s2+1rGsEBSNl2kcprRzN7du7LyGFn9NnhwI1c3ZaNwmMK1zcSgrX/p5LxElh+foR
atlqn2OXqHMUPoaI2O/jCw0Fnnr+nMII+fGp6GbdF1luweFHEVze6r86dWDULWN5
RxRbJipsNrrje/MsYJT4f2ka/5yAleU4ODGEhdE/IdgRC0hOSdgnBznEN42au8vx
LHaFNdXOTfW2n+vOg5Ls17ExwCGrUIiNrCEFIHedIGA4NDCfTFVdtiqJ3shDp6nh
Hm/d1CJlPAHFPX8wZIT0a9xXDm+KAA1BB4HSBbmqp3rx5mQ9LCtJtRuoczNyoqiu
WoaByUtSfmlgj3Unfsf8BItaKkO85+xbUsgEVLYITjbCHBEjg0eBx3poJ75rL+Ex
UVfPhYYcDGXFUTr9L0+eBJvZYszfQaRoNFYwVV6sj7bcC35TpGWgtfJBw+fsOSmD
bWk9+bCX96KwdZMWMtTzCFc7uAaTDuj27fPnkc87T+C25XA6bVubnzHMRVhQIdgK
pC7neOjSwhzO4GfZsK3WXJ63+xesnG8bfeExxk3rEz+JQhRluFq/U02n2tsGGtex
++JluWC8A9dtquB/4OIygRLb0FkwCRb50lohRjaZLn7dE3ltfDw8ogAHC83RmNuT
O/KactkleNpzL4G95qnhexeQrrUHsZa5ksVbDrGh6EOYl8MQ0bDvYnuloMqHBOQX
W4PB3ty4SbC//6An5ad6PARDcrIbI4jTe7KbggAGhvdrR6cCvID+e8LFtmYqO53V
xOw8mA5V5mb2fdgByMHCLwMw00aBjWWkAkvnwyOtcJG0pK3xMeaPgMEsgroLhT34
8NuljRsrao2zSvNCKM0vMrm2J2x5t81zqfJkQWaJjIlX0a4o6aPI0oclfYAq8Fbt
6PfOqIDsYbsauum+1r6cKLkZdGCuybtgYJZx3zNppKSt6ImM5dmb/T1TYlUZx1qy
jnObgVth66RE/Pmf3umx6Wx4ki/5KoHJWYNzUM9TbWOYYhUvxehckVo+etwisC5m
SKuAZUbnxSzIPnLi6YqJEan55sa10nflXNYnWynLY75XLdAQ0ByxVWRlOd5nTWso
IHKBd5loEL6CEM71XJa9FO4D0L3a2FTIbrMyCfTfnPnNx+O+hAUvIPsy1TZA6f7S
Z12zZKXso2ppi8+v6+MKyAedeu5Nr+EUEoua2Kq+IVD1xb3KNl0X8p+Lv2I7NxEI
2aLphU5hFHqJrpbsrYv+3WPgKJEEshPMVjuWzU4KzX+ORSG3E3b1/F0NYuYCLZfM
KWD5AUQPWxC05KFkMo3SYfSgCug883O8tFMd8cUGQYAQxihx8NhZBbYWIZDVfN3R
tSR/AQqQ0AU11KepzICJozIysk6r2gF2zrmmDGA70j8/IRZzI2h12HzRpmuAqhVn
Nq2Ik6Ki7Pww/3nrEAOCAq0jLGobQVZUmh8mtCsrSiijZVdIjBRB7ri9QjRc9L65
TQl13hDSDdkdtQs0Q0O6MShIeHlpENMw7jbtBXpCEVQrZyKTUBhhB5I/CG8dkhSr
+JWjvYG8J4vwxRSA9EAifzQS0s+Y8/+QP0S4ma1O05kvDBil+EZhGVtUzB4VbgK0
omvkhoTnkL3t27pthFSdBs9c0j0NRbHOPvNDzOgPfZn9r/kMLkStR7eBQFbdzmoi
WYHWbTRUeYVXZdcmDoZG/RiCSYAwV3KE9l26/42WqfR6nnTCQEMcCaw1BWBFgx3X
3StuLdGJoQ0eHE9thkmQIPHLEE9EtPMYEqnbcA2Nq9snRAVcgx+zOLhCJoEJMCvj
r6eObSBipTMLRizXxO6kFfoQx7aTXRcrQUnRJLxmOYUO/sMb5s8eL/0mHgcvP4GF
WwB7aEkpTvsgLop0n/OYJaHRk4JYoVLX9Y5G25jQ/XzgDdQ0sZy4anRXLQJzfhhg
0sP8p+3v5QAuprDxPavfeektVQgJzKca28A0DzoZgItodlVqcp73IkODcqMhpg5y
8q0vtDUj2Fhms2kFpQzG4ZvrUoT4/iJJIvbjVLds6tB45zmbSfqaqFoowj81bu1r
duF7mDgEcrd+8Q4znGOa9wMSxSf7ElqcEifbsV7WLjhXnpKdsFr7s+2dDerBE3d8
52HuZ/lYpCxnYEsmS5ZcyhxV6WSK6rDlJY9B2WJsbIyZOvGry/wclXqHQcOIwBa9
NIRla4e4bVPOEreUu2yR733Xys7xVSIXpMwXFfE/FGE1ArjiAUsvnlL0Ec3QQiEC
MdPMZqWP5vYNiayhtFU40QSOzNPmpETSJj4ua5e+NHV8Dbu00/aZbGD92P0B3cYs
i2ZiqJiZz2RHDMiRdjl11vNvIcjxMU50OxEiMLpZqnfeP+KSqN2XSTCBrT82zPHA
e3s0/tsQjrBaHDs4Ep2NY9fSKTi/ZoX140X4aL4B0jpBOiQLODBoYJUe0sIWuz8y
s+YcJ4PQoCQhG2ECUr+9v3UmmGg/4h0/uz/VRuQ+V6ofJ7eJIHopgAJuuD/zQXgx
FhNW6HA1p+XFrBSPnYqUZFTVpq2W9ZMwm1wQmgQlYszMjhnQyu3/1KciOPB1Hy3K
2qFmd1ad2UNe/yNHiHg3WxN22vkTUl3o6lNwk2JlGDxBvfAyh5ZzflKN4OBA1oH6
IlXztg+45SESGyNrfaK9IFNF2bjTegzeeBh7eq7RgswLp7JkigaaMWnGIJQb/477
aUu0G6GCFLBBzUQS3WVsj7NPrR/BRvQ6//qSQKGnop2G9GcAxWtmddksfJxVL7ds
0DsFK4vfNVBthgqR+ZBsoyVecUOY94C6jd9A7KaSLXsV3R7lTGsZv9mwYIQWMjXs
l6VYVzIGxEfS8gf2TBXNuDARgKFVqvfWH3We5HQlh5vuTxtWihLgLQZ8EQGntIyD
kikVLyqdAM/ja74Y+tIgDnByAEgJv+50mPId4Ngu7Xmh2Z0V+922xipOsjsbus75
l6k+GkLDeRwngEwCCz3fhW7Q7RP74eDsitjYroqZLROyI1YNdgCdwhBS1Dg3tcdK
vJuQslasjvIIfSAw2Kvm4VfGBwExV98o1C4Zx5UPX8+XIix/DtiRcAju/5uIY6tZ
ctQtt8YTzQAEKqRpX8zD8Q2kK4DuUJ+xn/6Air0iepbXnTM5Yy/GYq7yn7W0TBCn
2GSgFNeWaQrLc9Hl3CHr9j8gSlNZ9mOwe89L88oaV2e92J1nJG/Jvdh6sZoEUHn/
IvvXJZvYAJvksE7hQ76kb9uQlKm8+YYF+fO7CPK3XJ/uQ7cR9WtDleN4Mu8aDt+9
a1e1q4zCrPYJYkDc8Qo38ZtIz990R3OfsaLJBtCsK0I4TjMH5p6Rh7SxFRwRTKBv
ddjAra3MCAJJ5CGHqYJArSJTzaxfIOLfsjghiQeACmaNybgjVeb3cDGGD06SXx47
/khjhQFuHDAUv2XOjdVrnCrhYt3OYgxwo66i0TF+oPdenK81A3mlZIoinQNj4Jn0
PzKLHzlwYWYZ6SfRbQuxl6mFfDurR7bQtzMBCsgl7QWDa/MwoymboZhiBD8KSE9b
LGolXGiH8ojTQQvgCYwAJFI57GY9AiHfqntNvq62kMe1AagR08eZ2mnUC/XYV7B4
es131baYIjumI/NQQCEn992Xw2JbDzrv+u1r9FGxVFMxDB/J9ChND2EsPXnIO1Qa
G61Zx4qBhahWldCyphSbQXbV8Z0kp4ZOFE21zTtigXuOyPXuj2i3VRnq6bI/7Sfe
5cwEFBkzq14VRmVg3+bpbtDvgQOzj71Ou25a8jmi+DhahnDnApKVeCDPiueCo2Cm
UoHSt1v+ZNBBiRE1TNfU8y/SrqnPUisyRAk7liCZAUKgG8sQFcsoQSlLel34uZi6
fa5nH51fbq83TyIZ3QuAp3PwyQA2/q/MpjgbnJBo8Zb75dxArztQj+WQtzWuuS3X
YRF37yUTXwj7P6ryfSwVpBK08Xu37crXXnxv4lmmC7NcsLp6026sCaOrPJUVzBvi
Q2VPLahHMCXlYjA+TSmtpUWdf3DHi4UMXn1LsE+cL1mJ1uSOah2Bdryb+WLnASX/
/I8j/dbwOibMtpFLoHD/96P91DzGQmGiP5488I+IFBo+TWHWJvl42uM6cDX4iD0J
9coUIwOP6sOwZvO4U28gvYYhcXZ7VI1i7+eGoWcAR2vC8vLABdiALhxoVF+DVsaW
ppUrPoZZKHJsP8vjtu2dVcSyHnyf09zQDnApE/ReosI1OT1K7bjMu3NNnvD7IYM7
jSMmVLfE8u/6ZBi7d1ffSKhrbswjXOD6ttqeScTdf589uw5Z8ugVghUvgCJL6upt
/K/Ch7Kaxd7FwTIlixqmwmRo7oldJ/HxuQQkhjQl74nkzI05zFmgQkanFtJKXC0A
jFZYAAbSEOaA+VuMvhbmDZ1HjJV+iW63oSUDGMgkofYEv0Os8ITZmL4Ie4icDHWf
7tOi2H4f6EZQetCQtl51zuDLihTvF4/5D08JoLvg7uqyp4MdLXF3X1AwhqCb6IFu
kTIszKc6piPlMWhRZWCu2X8Uu3MazzP95wAgORfoF6/llqd3uasjjPHbdHPOv8pj
/YydNg72PdaG9WEjZShqKq3ElB3uNCYyiz8Zn+AnKHqbldm5gR6JAfyJAHdgJxNk
XIZDN+LqNwDMLISXniBcRYCGu6krk9LyL9VCFxPBz3qUlq84LjikVcHXrrFcupez
Wxb4pAzLs7zebXAVzh5IuNtuY+BZvYwm6QH9xMhJ/2zJCMSTHiwMYjiGrgLWyFtR
JlotvbdtysUWDyXlurDVH5MIKef9qS+8iqRbfHbbLGQot5kBfAmEKIUFxBOmbc8H
FvAmj/PVTazENGvjlYhSxBs6KBBFnWT9CU6WG3prUKTF7VpzS3Ml8IY+tSHimXkC
Om/kq4x921j9lGzzLLYQanxBjJzLD8IWvAxNrY9qRQBwqiTDp7B+vJ/J6ZtHEIll
frByTcF+Giz8tG5hCFZMzl1zlwhyzFh5a4nJZvuLAuBvMsv38Wyx2cfvyaxXBEtl
o9pQY0jzY5mVEF55fA0mKhN4vvC5r5hFG/93/dQ+YozY8mncsH9BUJY7E52gfbDH
Cdi5JbD5duHiqocU94/OdLxdcW/ABayBdUzXkg0Mmw8UbXuEYzWIcp3fMcqY1xZg
ORNwEO7DznY8caBZlBeR7Yj9VI60V2K0dyzoGkDWorK78TJqG7YsUspO5kr/SZGQ
MB5C6lsW9PjOA1R5MTJnbRDQG2LMGMIMzw1BSCgaEGQUt7ywrviP7Dfa+ZxaVkQC
Zz+QwcFJgN6r7bZrK4z3oF7fAhsZS2KWmtpnWkAA9NmQfFB1JZevOE3KY1N0rGl4
+uSFRj4Z9TMIV8xsTFPo+rd07T2Ls+ljDQZ7vcQIReyusJdJET07cWck2G+u/BF5
K+FfU9e2X4BVe/flxMOJUQqI5BYhVjoe+Xj58fwUAiwXrVVMYkmKPX5sZgmbBSnz
pNahM7TcmQ6m6dtosP1JhQRokFaUovcPmkXorXljXx+fhI9XDZ/VpfpCWoxUzYT3
4cvrDeTZWBEcIvuiYipFv5t/RM23YBYy+BkGHSYHUgdG7hkSD0urA2CzdW3hU6ab
/q+We7CCYnwcNrsoED+7KRywsthfcvHsIVe1rGtcmin7LJmW2reY43CVCwbPWmqR
6ZqOKxXLlg6HzAf8rGAyP6Whe1Dl9pIYH9jE92dc1vGIdXTazrDEh/LnG9M5Zkff
VTLW7gTSWUGOaUKpxIehsJxoNWuDRdMBq4CMHGYblizeNqbz59D69Jf5PGlks4iq
9zxjxFXjGq9ffrvOdRsqS7Lm9qHQ5jOGNw7+/uVNUFfFMEMH0fur/x1PrPaycPpZ
x3uqk7WJOH1aU1HLXWTLCOA1eeb8GlziMdFB6ezcIloLUXWtxyladfiLNFMpJknr
hnZPCQk9JQBFPrcwoiaFB9biCrVianr1J0izT2jlu+nH+9mMYMBg1NaSkmN0tOEm
IsVfKSesdGOYxNR0ziyPKi+60cJbsq79snsLUiIVV4v6+rfAN1Llc2tNC0FuX+AW
3X6+yfG3yym0eppopHYOnOZYxQ0yrKDpR3K57Yo1Gqok1dV705T8EYNBAR2CKF3p
7rDm4HgIJwBkzqMH9JeHZRgeGybZuKxq0+cgwMf5hzY8RWw1wyoHEwskd5tq4uI9
FkFo0YdVyY/hQX4Xn2ecxxoPPwsZMZH/2uystjB/clxlqtBSUsAAdHWPdUSI97sq
vM+Ec5Vnz54FPl38GxkgWNjJ+FJxq6EsUSL0zi8f0paTsN2jf2jyZXxXQtGHT1UO
B3YSo4NZDonWBEESaC/ziATp+qb76NUkkkv00I56RM3vYdciGPEb2yoqUFkD7vkz
57jmhNn+tcht2PcBiH/YXmzlBqi38wsTVUwapJ2zKyvHCgPyN+AgZFfbame2AwP2
/u0PBJojhc4nmT1iPAXgTNESJl1Hfrol4pBlYWyjNUGdLBeRVpA5/fhAuVN50cZ6
faBHPfewPiwF53+rbA6dsAQQPFS2NXUNwUxmAeLWfANhBksFGFbbYOgWLoVrrqX3
typCM8HrYoEbBenRwh5vPQ6NiVkvlk4IFiqe2+MWTNdhR45ZcZ2WpsDOINOb6YFb
fH6g5iNXgTmDjhbf87D/Xnjc83AN12WQqqZ2czump7/XmE5fw8WdS2gTxpRsWyGl
FKUpo31ia+r4JvhxHn+craTemt8r4Qn2xuWh5GSdlPyMC/vtUcTcuEW4IhxhMA60
FXoBp2XWFxdmL2TzmbFCXGWzEiggvQphzKpuw6sGor597I91CPIhMK7nWB9XIrLl
Y5rzHXBd444K5z2NhB3PHkngFYlJ7OtRIjmmfFsUMEdey9LH3QnqdfwasOTg9fon
xzYXVuG7BNhScoXpbD1SBs6elbwOIuOekMRdz6U6bef4JbbqJ5HNdYB+kjtH0XC7
JVeaJGKOCmYCGLscBVIrvLBKgtXxMVqKIfsW7+RX+Z1CBdQh40Rl2GkpT5le5VfA
3lueumO5E/3Z1KN7y9yoFKR7nkCa0aX49pwWp6VKWEA+tkFccnf9MRMJBrPnGIBw
Nzf0sU/8JzEh7/n+SSV7+LoZl8of6N1S8evuYSLXZMAZiDNmkK+I8KyYd0C4LicH
TpgUHqzu2fh7HwGJjha2708pg+aGuoPvvBgaAdyrsUFs4m5ng9Pm11wGOFnij6hU
JSM9sUSl4TOc/zVtEncgX9+CbKHl1LRzuIDIef/ebxPw5ebNPq7RLgcn0vLqU0OJ
aZQ8PeMJrLWj335lET0skpZcZY/iyMXDG4kRXea2xo0kn1mRqP+dic09GWbv1nvN
14xy/Pp0o3p5P5urU2vS3Cj3rIpbUTdlODInY4NMasBdB/x5VJpu+RbDZOar5d5J
DQH0dnBIfXiLUNwVCxUFdhEa6gl5Z8YKjwFrV5m+tiuwQeFEoASKBd3T8UIGlZa2
gFU8I69OT/OQbG/wqQTU2sAVpZ8KsjTUTziKnCUi4bNfS0pdmx5VrYO9KmhE03zF
CZ+8ofGwl0SZuTCUvdxLaQPwiJ1j2lcDnj9UT3CRlQtB5E8G9b66dJY0HOElitjm
NNqoFAoigtkiaLEE38A8h8dAi/0kZg4NCxT6e5Pkm0CkiW54gy/2S83goXmu0y2S
YCNwghrsNzU6b5hWgNcW2iyd3rddPzEJ0KMHzrLIZxevNk0yh//dq5gfXECx0dvX
0IMczT1uKk8xjMEdk1mE370XcAdC2utb7/17IPGRzgpooUK2BOiecBG/K/EJ4UzR
wuJegJmx6fdi5CN9lAlAH93X/PS+NjMZ4vX6eae7+mGnbGbXoJuhCpfNVhxxT+AQ
jA8H+floePtJu4WnwPdbG5W+537743foDgF8xa/6F/flkwybbx2k4xlxIg11ylSV
sqSSN/2IiOsqocOwDV1SwCnt7hJ01jg3JwhQC6QDyFYHr27CvvMnLcvEv1TNYSQj
vEoC52K/DKgLQeM0Q7Oc1aUQqdrwY/l/C3NwxHx7Uok06sR9sfk1pbGhEoj1qVpR
mfXwjAuOrUviweqdv+7k/qqxNhGf9oeny3Ib6uLPCpP5wwQDSPKeqq07iRW8l6LI
RiLlrI9zTsC0dcvrDA5ZO2k4OL9+D1cWSv1SWkL2UKphZPecHFMJBP1ltUHXZZre
Cj+T3RYAu2ytkFzvQa4van+T9A6Kb7yp2uYWbRiUUHwy4wWP0ZFN0n+XiHZhHYnf
JwRsQUjYY3hqmO7NhMHLHjF9MKwxdKVwY9LF24vSJ5im3EDbrtwtneaNmwiz6aEa
OjATxeW3KnRFIg1Oddp0/rTWtzdCH5+HnNXjPl2NEANbU11HRTohPqzR7v47mWei
+L2qBVjDSc8lATtUs3fw4wZw0yUjE8D82ewah5xebgmaAAhTa/la2E5hTYJ9ZnWF
ILeA+PdCyZc5zU5LhJZwAA0jYFLwgQP1s5Bl/ZjDemKdpPIqZVvM7T+NMNTS26or
0AHskgjV+ztPX+C6q+1qUrx6CED+x2uMXBlfBR3oB+fiqVXH9ie5v0p93ycJ+nEs
hxYhHKbquzNONaYRu6K++DLxL0zRpBfghwAk2rgxBwio+cgVJZI294NIki/w7znS
rapwgHUl/ZuxcSdI9QGfvL6pfk9RclFDtXLItluJ8NUrHcRgypkcZleitd7Aqn4v
mr6KKam/l0yhxu+nI4szGWsN5S4Vx9I2fmJkSgoB+69u9n0e99ix06QNuJ3Tomds
JoniKwtNYG//0PDROM2tSHCPtA/+9j/SZCSR/l0q571nEMj7j2FxzOXe967e3PtL
xb+d/eNE7pdFf7SBeBbbeYyaMnnNb+E8j6cd5SmQ07CIg2t6aGuc1xDNd4Fcm8hu
iyHbl6bpEzNu3fbMgAPfMSfVkDZIy9jdkfDxsIQy5c0eRgljQY3hyG/0a6TnBmVj
g5kHvZjvc1yfcgd5Ap71cwY7HoHBZqpxLVMhtXYoI3KCAw6mv9Mex0d+z+x8h2NR
0SAGR3zYYOjXzkyotw7TW9+xFOdP+4Y4XlmUjt8y3R+DrRmeO8ggTSgavkPXDS98
CwCJcsnK0xcHEvvMOw667bKi/ex1YdHv3vII5IdKl9dF/ZNkwjjmQ2ixjvB5+E8v
+kO4WgjnDmJpVVHOEh5bnDFBLS0KT0oh65DjqBmFdrcrgJEwzqOC0r56yvrCxuUQ
woTtwpRf7bV6Yet/+rbFkyBjd4oDpoPjoeRVB5UX6pN6w+egHuDnbGR3Bi9nTTxI
amCsHOeGdwIElTcPyTdk69NTp7EWANxFd47fynChBb9djfKX5r33X512OsMEb+bT
GswTQ0vBMK+/la6g/xAzYjdgHwN/nqMqYFGwg89DkuljLOcZyCOMX2zePrc8yk7R
Tf0pD+fCfhzKh0qs4mKSBSdGksUCznp4bQSVcF68daFcNiIfr6CtY4JEafFf7dm4
qyvfYv5IDMyLI34b8qfzgSzFJqPGvLR0VBlznooZkEIgCjEwWSPQ2saHo2FKIxld
cH31EZ6bNP4CDlY+WA8dIcaDlh9+WindZY7ML4oO2r4evbqhi5YJDxftTVuoYSl2
2CgE4tyFcc4FOSYGDr3g9Mc885B7vk8ix4M3Knko8uSVxpjqgXHFrUho7w/H2kUJ
fTPHXQE8oXngedpRN8GBd9PDNqnX95uAD8M0rBa+6tAzDmOZU0GzbrU3CeY1y3Jp
ueozlt4ZyHf4qUn+3ADEfQ479pUPtKgZpSaqbOcxRYqK5dvYN3/Qp3gYAzP6NTTZ
JrQPo34sOdW86q3/6ppH/DBu6E28WC7/GCgZuu0Qh8SLcuSB+dMhsjwif7qEBCNs
JoIEW6igdEhT4L7aozZRciKYhLb1DbTrw60lf5fBbJIBP3ePX7gcZ1n23GWr9Hip
g30fM4wWDMbNJJe8dmp8FzH3kY6HGkySjw4aTBd66c5b2E/s6b4Tx7q5hAzO+E1J
5dqxIDEdCnLMVtMeoQwKga3bKiQ3g3j4AomM32yvvi/DQoh+v2ctwo54HIPLytRO
IddgDSwcSnCL6MA25yLz/opjFpSNY9lqxt6HEGIHxZR7cia6lrb25dEIeeR/ykA5
41uAfcCdxc/QsLGR+AeyPIlyRLWMJg/mexH32Wn1GZuQlcKuCwwprtJlxMAwCnoU
MY0R4ico3d4ubMmae2AAvsN4GHsrKtzezN9pjJTP9a95lwCqIkkL3Oe2SZDGgMFE
UWHGYZbht4152Isq5E3xW0rVXvUUcNQm0BIJDeHTphyxhxEGQeT8Ul572BXdpI/b
XpTEJBzNEcWoHCZ0eFG50qriG6UFqjWAMRBQwfE3/dbzzy9RgDY5Laa4n58H3X9E
8Hr/sIA6gHN+YLhjFY1MOsRcOPf00zzjz1J8BsE9SwqowSkLLhXM88xDG8jFWWRl
7QIWeU8CQWq8YAMjrNmcoh+LP7Dg7Smo4qA9Fdz7nd4Kjsvut7Ec32TnoYO0fsrr
8s+n2IHBxodFbpVMRc1IV3uFjQrwjhKZhE8vmTb2xCIEtP6Yq3f5qXFxky7Zzp2A
WzBsoSkg3apUI4w8nFQGlU4SD3ri/21qGxU2SrXCu5OyGWtOf1NZzfZgNKNM6jBR
TKay3JC1nTXclzTzykGQChDMB7CIOPJChI9w2bi9orN0FIIIMenxEflxrgyy79KK
3loY2rzskDo8v6X8ybodNElrXQw1uRn4WwZrfym7YwcQuR/kg2U2lK1amnf5z01m
UyxzrpC9Y2BAGPw2yd5bC4hNp2gsFNWiFslS3MrL2BGBKgSppNDke+BUGzPCO/yP
r+/y92ZdM2C8ZB31v09epK8aw4x98nywDx2Sblbd1scLUiIkjRjavUWJBWZ0rlZ4
q/LSziR/IE2XAjPYHjBJoq1DST9behdEI8SmFw3Ku1sA4hwt9nAuN0hJXDBuGyxa
ugYh034bQvHFTZNWnsrBz9lHp3JJ8x35NzM24c07YIMcCIZRzo4AjSCHHzBV0+6/
avnGJkCEozP6FqgAJPW2lPO7421fZo+ot/ry6Kej1ev8m6JYQxpQ58UhNPxJj9O9
Dg2nJaFDYhqWjkZZCoynxeoE1IvX6CcMRoI+Pvo+wGu8irYJBRVOW6MwG/XLdtN/
6+xM3OCG4aDIwZfmNdMJFkhsKX6rXCkRsjBzGHEWbcAIXP8ZfKXocFyiHlH6ZzSj
NT4tgqtMThfq0UejmAxBs+a9/jtQGZh8PCMJ7QJ8u+JpvmchqCHtla7Nc30uAoFH
mwYuP5RiWM0J99LDP7yJfqL/Ic0KbhmA8qMQKSCPQ+agXPPcHtQ/6QS+UVcAghG/
R1SRR+lXbzqBllhepwXPv2exrL64NOMjdMqUMzsGQuKrxVKvqDukzu1CWptfomlM
zQWXo+Fmz1fzDNx8G4q+e3VFhf5EwT/8XqHcRyvCwOOTw+sMVTp7r2MaU1UJXSU0
UF6uxBnJZt21sqjzhpIqzvMg+YaZrcf3M2hUgu3IEdXpAjAyYbLrCyIO5ykXu49e
wCHBVqKjCK+7qGtRa4+CepdRsT9KsL8VP9ek+TrAiMEmFCkWvz+i89ECLiuD2vJ3
3UCQdkBMSXtue5cApgYKwngUQavWDu1U9hPCnAmSw/MgB52pGp4BU++VRe2Epu8f
3UfAil8TYnQZVMgnkcI7JPoVSiuodJRj1bH94WB6r8JjfNMpcHnnVTGRNC74/ag1
yUfsiAmLvmalUOHF5Ke2vVk+jR5OMZ+SGwUGtJRdqieG6FxFDDWLv/w/neFXhgVJ
pocL6XcsipaA1xD/E5lbasHDnNco/Gi6f/X446fvgU7IQhpJPA8IxEei/kw3nz4X
4GlcxKGJmShlOIujoFUMugLl7ZdLzX5yge3ff2g6fXR9Kcj1yLrcbvJRqyiZZ5ue
liVCrXWvULSZhJ82x8H5FhmWD4rb2o/b1FOBCJemaxVZgsSC9cOcEY6P8eiXzrYo
jvB1NwWAlotDdDWwOmN5gMvM5s1GPDo+zUqvV8xUbhhZPB7Pfu/4F8cPIf2tJkqY
2vcLq+HvSJ9VL26UyoB41aQ1MQsyUIzUkS8tn3NUwADjrpqblZU9CeW9UcBFXQIs
3kVQkM0uXqqGL0cr3h38pCyu5vGgIZcjQ9HnOe8ZtBdfr/ZFaSKxoTGQC34pkGqP
lGX4eXMvFTIEvx3PG4/t9uyteM4a939St4SwJiP6A/sRsQRfvxtTpysSylH1mypA
7eayVELx2LY9wJ10QBMoCLqtPZnx11q8OBH6Iz+YDivD0sdiPp9mHeEpan+xA1gS
bkZvjNdWqtkdrbx5C8tM5zS78EsE1B6FCQUwffFAajeQ6GzP3Q2v+VHx8/w3AOf7
1yIP+CoK8vS6+qrwfvAJ/65D3pSnZJ53LblcI/eVCZiWsry/vTUeYftUe5CRLZz+
KTaPC1SR8YF++wfmB2D4iPudRQiBjYy214Cldudb9lYAitHGFiBPl4G9uG2cMqTt
bZ/GiPiksjH8VPns8PflgwcCEpLWrSE29ibUmqVkcP70YkB69+z/DYL84KVlAFlw
K22s3mFVsvloOb3BGeGI8trcFe7/Mnaer8eVG8Ggr8QPHbeCMZC9yVkuqmvUiGmI
EyemXHQAvSNtSie65DJE+NyWYeNwMkestQ9iVNzsQ52HR//wCtSknGL6amOQI4h7
IwfZHPh7ayLvsQJUTEKlzEyhh+2yHsvxVh3HMlkchP4WeqQmuSRBsNtvmui50zbh
ly0SJtgxaZzjKmOZuUMYOhMKltcGSS9CwfwG8VwAA3BWhXQ9r/z99TDz6TUCyJbr
EItBmaqDnGsRr/tCtfngQueLCqZmXGTe5qQcYFkoqOe6dJJeSdz2Xz7JpSnxuo9N
Pd018Au7o7qXNLJxTpiVp9wW7og1Lc6dN9C5LC51P9hpWpiAgOw9KTXGCTcB2B+0
2zk7j/xnQ1EEtCgXllUD/Ae/YVSjZniadeCWiM+V8FkO79y7o2cSxBsWM5JArI3v
f1bg15cP4D8ieSAOh4Y+l6nmejqGpibGY/Sm8IV0ce1ystqdfU/2G3shONdq73fC
SFuhfdYFqBtd6XjYxtPXJtbDp1Lf7+80m53E3DlaWy5WaG1g48ihsOTSCYbDXTt0
qZdlZup2XMyFDEyQsHC7q3ixd8ueTzR0oCqOH2TB80xEkWGg30npyuXter2vFJZR
ztaOwzBvps8xhUxR8IwrIDdJkKwmiDY/N3s3JBVInw2MRthryleMrbm4s/fy9BAd
D5/hr4keMzUnjvaNVjotXHfi4s68P0o7F0hdN+sQbAHkOJuAPB9uW1tSmbIVTyrO
72X8LekuEANANic/Vy73qeFY7w4RSONqqtmtJ9uHUNjFMLhXuxO+v/Ot27OUCZVN
UU1Hv0KQtX63cwWnMmUXKCdptM8rWf2fuFCTvBNi2SqeCYlBK/t4gJ0wNvk752ya
fXNTgDaRy0oRIOt6zAvoMWgzS1M5XyUw46csKTE4rRkdSuHEHSi3Iu8E9fWvSilk
OhR6U69Ey/B2En1nS8+zHN4wo+vSgLksZdCAhj1gU5CG8efbrNQ8eyZNCLpgmvLY
mbig5858eisYI/c9WnajbPjnA+fzEKtA7pgPblZdxsJvF73snNIfoBOhQdX1w8ci
MUuXXnQjsMRXQIemyyzfwMqt0imgHk+nosiRI66ljTSLH10VJ7xbRa90HX7grmFE
0/MOzpHsqX/Lx2axw4B5jAFcQLNeNUqQ/I/PUwjcwVTeu+8dKl+GDI0umTWsWLT4
fIzcwDqvgbhYnp67agOgnMYghECk06s/l1NPCrSi3EbFT3VLqj8UKe4IsJuAB1EY
Meih+yuwq815q/cJ8yEVtuJFHypy8Jvu4qipGcncDDoAy0IrBzGb12d493cNwG6B
AtF1QRSGCFCDPQxnFHnhhM241LZT1rEaCazXai2ucbfgsBVjEl8bZxJ4Wlq1vt2F
70jtBP67YhtU0tPMzb2m9mI9ZgaNOWgGjBcqXfa87hxxpMntOrIelldiwpqKwHDE
CooKcXe+O3i9f7MfyN2P6xbwy4/JD0Z64t7GI2Dy3gTTTScr/BESDzuSMAku5B+n
AAzVO2jSRVkKHZe4KywTsqX6GrxQEE+1n5hzVadB8Uak4Zz4f5gj633ZrvL81r9r
fpB7CDcEKQxT66D4rzaOUMUFWKpkKZqn/thMH45gsaJ+sXKHjgvZr15KyJq0GvuM
hMIhU6c5pNlUkBvHFFq2muG6TQU8xfrTnbPHgx2i2Mt/1XxVGthL3Xqy2k60+Ftj
1nc+q+MZURmSm65cdeg1ECULX1IvlG2/1PZB8e3+yrigtBNR02hAe3g+7O9LtWQw
5UargdZNMGINHDfwjEFxs1mld46OrcWNc8alLOjhx+b/+BfPxpX9JuvzKdpt1fy2
H2dykve87L9Q6hDIsQKHu9MG3NQonp/9gEsAFYMtpEGmM2Efnax/zFgYH7uVQWrk
+8TDormuZEg5YQIULnIt6fFBqB3djSYQBEahzATzss5Mzzb3+EpN7PR0sxM61+JA
0w0rVnmx68k12I9chn5DnFSPq+L3GRvqK+1RqmfOTc0NuNAc6wsGx18TqI/uNFQ3
+Gmg8mnKeeffN2lHUaKU5MZ0i26Fdye5a5KqBTjOAtGf5skev6MKrafFm51wWuvO
86x5Fh3N3ZXQvYjxfdmQWX4XHnz8PuLbcaMFwrDo2b1NTlMcZxRgubIouVQaP6uP
/C+NEu7ghHHPEVLV/JKxtRiJIfyYQI7/yis1j4NbOYfAcKBU51P2eYcsd+IpRKnA
KYh02YLY+n8Pds2MGpeLKSEfuhh+rDUlvMMcUB7tq/Gg0bGNyCJkr8i0SiUkciQc
JrqHv8plgM6oKwO61+zZ7FLkB8tdHU4e0AvtzresiDMUPvj5robzbLpo1JfxE/TJ
raGqC9nnKDNY+1RBT52TSrt3QG7vyJd4WNYiRhU0Sc/0AYxdGjqTxyYmfjhulo1v
G/i/pJYC4iPVaaH91fs5vWERIWMNPp43OAG/xiYlDcsVacunYiobQQ2ZPBrir9ig
vF2rwRyMncJ7PEA3CW/O8Cb5Hs5T6IVbgN2/tywr+J44rlCTvGCBYd0jcDPGVijR
vMt788Wz22W8q0GRZ+19K7s1GwXOYw+ISuZeYyGfuXdDlsX9grxC1IUO0sh6WESW
0R56zbmIPoOsi6p+2qXppySNgKD0psV0DgYByRR7NITKjcN6SVHkc/CD0g1xMxUP
DtOluPApqC8vJhqAeG2frWPRqNUtqIxscnzTVoo5MkUHfzRrXY5X+6A/Q0AcbmGe
82QZhp4yqZWpWScNRlNJ/LLz1f7Z4+mTqm2uQZfIK8nD9LFauyY2+XON7Ugz+s5B
ue8i752Ion5f81yz9PWhkAeyXBkWyvPU3ZFiVQIK0gAgwMnIdPDEps4SmrnuOo10
51pKHPjMnSdFN1JdE8HRu3xpEAPw3QrQW7UL+fbcw9BiadYNVJcMFnKnvv63DGDT
zS9rIGQoGCbD+JacHIbzLhrIZSDw4bcOyOnI7DB1lRTV2bh5VzmOx1Psl8TETDoX
yI2kBoCukwUx4rpujDFSSIba2oe5fLnUwTyaJII+2jmZ71LsQ0LbstjbQL2tIRdH
Xr59sXi30DAcDJsOcpDDmA6Bh46LRSKNstNFu0p4ahsk8yx3JxUCi/+hfPcCyBB4
51UXKUTUYLP2QWpKKOdiqiyTySENTDxipcNZ5lrNx+jjE4GcYO74xD1UrEF93SnF
O8YH0TQ04LQd7SCzskg/9uVN36WziUETBVXPh6c8K3qr3Zu0U+Q3LOEbirkV9mgz
8iKJOvl6HRZAMnSU7w9R6kEpWaoQN+c0o37SD8TH6qCKKL4AffTQQ5eqcyC34Ek4
NfZVh/Eh8Rn6sZkntJzWRCILYDE6E0CoKtELEYndGKHav2VqHICUsgnVQBdarE/f
rZQgc1OAIzg2HwOOKDgs/9WoYsa+tMiD4YYt0rcBTFi25XPzHu+Vowi9DxbqQbeP
RBwLejRE4kDLD0VBXTxPGPtndsyuJcd8KpJp8OEmadNe9RNuMrJ5hgdixUit99OS
9x2jJdDKgD+o4tNqPdghvCff/UzN/QBPBh5zuz+xdy6+n4yBHRIp9MHsXBvGpun4
4wGFIiiH6m8vE07uzzND6VAwwrC3Z+QmVmvcbODkmplkDjiUvkE1ZbbZl/HZsg+8
jPKuw+v418GOVMAjS9uZd6hk3z4Mzu55gu2tdmrVlw04GblJBxmgjNDybBUrIHn3
VgLemkyt2bztYgFcsFIAUUnr2Lt5W8oyKW8mLxnbP/3D6CDUefzjFcBWMjznuLP4
FTVz09S1oVGIz3M8ON2CqCuMmWeYkYrnX5KvP19qd2wZecD6vjJNXeKHomYiJ/iu
4lP1YVsWXff4yV9RByhs3aSPcq72z6vR3A5Jw4ELCUzhh1epU81k0Nc4NVWu8hKC
CpFBToL3kuYY2Bhudt44iTQ6WhTACDfaeIqmuRCQk7XPQIhWIjw0Xgj9b0y4Zn8u
g3nFPx9aMxNRL3xG7okgmS9sDaUE1uHbIU2LVAuExkWQuq9OlFp9JzgmKfCrinfx
FVTvzgH/YLJeWvdaonfS/luiZsK+zNJbdbWax3FUdjSAwLZc4j2I8a4/KLJZdNh8
MXWOiRIgaEN9vFWzaWdDhB2Y3H52oRosdQb8wZ8GpkiOnD8X4WbdQojQoBX0KbRP
Vo10dUNAGiJmXhqBmqb6iBs1YE8yzK7JgF//MORsxwjlR1r8ujOT0oo8GOfO105w
kEqkIaCx0WX8Zo66u0sM9KgshzU9b0WxpVKXlzeP5QK9oRwSrs+5NCt24g4VAI4N
9l1YjOMKshE6Uebm4SYIn8bV6/5U/Mq8WLw4G9nHdtl52fqhDN1axqhY8l4557cZ
m0pAWveewvUMH+KbQRj2OQMxZe1EC5G7VHqgoBmyb9yxdn4V8I3Z7UmfIaxMKrWb
WvObNhLS/4t06ADu5BvklULlLsvWMyKfivd/n+lBHNRxcd6Zs4LQ72nqUUa6mAT6
Up10mtCGiz4P1xKlffxDpOoa5RQGjEIvx1dS6y5Kr9dz+V0A8K/moR5xCROwvMsk
tL/uWkUI+IRINogmHUpuiVnDboX32CoM8teihEsTjyVVprA6dwmCJ28wV2TN5au0
E3QVjd9Ede4d5grjgfL9xMTH2TkTmVUDXLzsd87ujk9Prectk42Xj8v0rW22NNBS
wWTSLK3VXZ4gx++j/puZQRqUGPtPeolWL9pI6yvQRr+Zro6aC4y/C/9ujTy+Pwv6
Nq0kLa6q4cNzDdAoPdywj/lNSZ17p9rrWXz5LKXRe9tGvC+jDDr+wOX3Y4TgTXum
+vTL1s7im1sHNsaDXM+bqdQ7B5ea8dJrgHf/Nr0nshVxII1FO1ktLsSwMUy8ImL3
QEdNyZQyiVa+Xyd7N1MOpntwgAKI+E3ppK2V8WWUHlG9g20Slmi3ENHj5gA/4c/y
Ve7xEFIE03zqqfmoDv/5RikhbD6TJn6uMzGRnfaCKb047xDLo9HPXFy0Gsgi/9fo
qwRNroJh2DgdsNc8I9NKBBW+t+e4R0ja6TeDD5A8cZHsdUUmou+zhjWCYTiGwh/C
6jrPYQVL7JJa1PCigAEE5s+Mp2sQzyiJW6U1zBv2UwM5naQ/to4mAic5I77gyAgr
WkZe81yfLdsmCDnMLd8NiquPFeha1ZBr0ciivcvaB9UcrMQANmvVrzTDWN1J08d9
vr3IJT6As3Gpi3IQHA81fvB25DdFAhUDZzlNLSDC7OaPXE0CBULg+ZZROofei6SX
9FQ3Sksk/r3LyURVNbZWOearRGXNyH2/RNUJQglCMpd6LenK1CTBpQO0wg2obdX0
EaVtMxBCR0fxduc7iCaDM58UWN/mlOQk9YJvp+i5NSnoEs2KifbrDIWJY0iR2pq6
JDcbMe97HA16v2/qV9k9Yv17O2nfj1+swIY3IWD/933nBR41f/2ryMlhTYIQ8/tr
qoOsZSBT3QBUY0uv3dE4okOJSOMgM4giUzDEWHUVs9mm9CdFIwmWDliYUXC/1nev
rCXk7yx90hs0uuQnk/hzyPeSWs5s4m+N91f9P0naCRWRu+8ZjW5SZFht0kIxOcN1
qyQD+XQSdFli3Q1GmHrFQaRcsds5Df4aVn92ZzWmWcneiuCDMNoDzbbn+4hZzoA5
bDkQyL+Up/awB0Yn+u6Soay79qNrpLZ6SI0VKp9PAtzjM14Rd1kYVb9rP14BjAfY
b73EuLQ29gbIqfRy9VoE5bh22ZCDIDiL3B6YzwJM0GjsftDUB/AV3VaxoCk2hfrg
tYEh1zhwVG7KCdlx9i67cY33noXaWs2WJLO0LeoNGQpTzF5zhgWHlho1zauZAngb
jhkS0uOCi4Qd33WggUV2IHdY6DlSq9u9UGfOEjpQ073iwHiIRp44WgaQ+kq39JVA
W3kpDtAa3OBQkmySn+VVr7L74POJj4ZuFXkGw/jsyG0s/ghQDYGy1B53+Sg/uagK
dJpGdXePN/MydZY8plXHoyIvBcNETZpjGnKvv9V57JLUqMhbAAsyBIJqLcnI9GOs
AKFnJxzxeX4/bicxHC4zb1Cjm8801pW+XAM9GlorIdw2fZ3/oHqSGuHJgqe7SVc7
tB0Qn5VG0mpptjk/iFMwTNb9NNdRUmAgP5itPmNpuIHMf+fdbryeKElzCkdk7bc7
7u17ZJahJvuNdhCTnwCguUCqb2ohR/7pj4gcDwyd274hM00609FP5wEuv1gYFlZJ
8TAZcB3DcdmmGY2K9BaK9be69/C29l4V0mVRw0aPHt4WhbOTlwGWtkjihSf8rJm8
gsfCzgAcWnonH/afom9FKP8p2wqIJac66IUj3I3W8G4xRD8VjBXf0bRBjNN1r4vs
C/o2mjBGfTyIeYelZbT4gxZTx7qivC2MlWh+NElgskzorm7cwdV+soemU4XyhMmB
Jif2wVSUozzvzoaL6sD5FAZdVYgs9p2jj4viHoSjOyryV4WrHqCkt9q3cGF3Be+l
ZqsU45W6HlQcREfHHu4qVdyU6+Y5GdyEcVrRZLFOAw522q1IoTHEvr3KVAcLsQhE
T76LrbgV7ZK9tYMJfV2/2iTWJJWqeh+1vZXiI7sAhxQLh4pCzLRh6sFyDWWnrQea
aJnz/b4OAcUMjF4AArdc4uF7EOhokGTecI3VFdfLtyyORudNODiezfV1pe7O2ZZU
hbWh8Suu0FRSj3hkSjuPxJyHmh9YXm0T07FV7q2GXjo/ZqBQDV0t0hLaVFvHHp3J
ovYmB7eP0BEGRiUQj8DTnEom73YAQDSjQ8lUVL+C5L1kcKL53F0wbL/o5PUGyqzX
AeO/TeYSR/FwFyItUj2Y7OucvWuG/de+szHN7pMwHhzuoR9h7r1F3/WklkP/4CDS
7SsSIZRlOv2RWzvJ8LZmYFTfApgspSyxJPz6Z2RN4YAzpwSDhhwwEzasSgNYqjQ2
Tg4+RB52tpkfQcUV9M4O8Ye8nZM2Wmjc2sS3bYBpoFmTRqXNAhkA3WycY8pwEquS
5IMXF0KMe9QXpVmUwd2Fp4hWnMAgCikUXrfpYF2HFpcGHJjoHDFcZrl9E6+yAR8d
kAFvDF0Nv1hbycOVuIf6nYSoVcNxZacFO1J4sVs6rb6Hlhr8qnVHLePGS40jywbu
gk7fzYxiK5TgImg2N5vwn1jrWCMhvcABwq1Y84/RUogR5L5kUZj3dg8vTN/lfv/R
gkfsCP2lP1PLTjMVbaXBpylhCxvhvGIbEOrf2W3CVk50ODpWVW2m0f8yjQjc13fj
BY3QHGEKCXiDUDUb45bli4T4ZPcXPEvd2BzHxI6H02Xq8dQDVr85Q4MuwLzW2j38
/ZCI0Ror01IE0iS37/o3cP7nm/A0963R38vA5YDXAd6VFdHjge9vjIUpd4ZPndYi
aN328EIS94GHwlfp78mfoNMleQftU+aiHj9v98cZk8jwycQKN0rBZoc7BS7boK1A
lMa/jA2zQk7zfYzD99qB4faCZUrJrn8SbulsLBTpTgF4ITdRSt9I7p0IS3CGJ/Ki
6Ozb3qNaKJHHAa2SF/WbxwRZeh9hCLxDrBMS9VcuU1mY0pwe2CLmK+wF8Uk10XuY
Me6QTUsXPGkGo2dLvVZuU51NoRz/Qyn97NB+r+HSoXqDwap5iq93Yqfz57ju4bbt
nNFekYNxwNtoDR6kn0ae9hQZ5JHcDhsnaHJlScJzvPWS6VwboGSvzJs++wflDx2f
XJ95H/KyL8GtXiRRuGAQisvfHIc4quW+wFJm5klcvvc7vDX+J41hXfKAaFgNWOOG
SYXeijytR68Q6kjjaMm7qx6ud6u7CusEjMOyv6dnXuu/3vaCbzZdjvaLXsYA9kD/
6ewG5hmuvtj8an9aPrdlwjJWyShtyxVhBBKPA9W+goPIVTkF4DhU13AguVcLF7sw
xWxm13Z2nylva2rJ/YwmKiuxS88sBGjfma+1AZq6rIN/Kg4hxZuMSchPNtVpKgjX
vpsOgwqshi1RLfvBNM0NyPrMrS4TTSDsqzWUdhd/7jzXDVgo7Xd5cD1NK31OHq9E
kRF5MGfaDS8PdIXXIY847ZpJ64a2Bxap9zkYEpjJ9/APxuMmfiMNnNS1yowXjJuP
9kTl4u36BpPpKSwrBvwlg/+ctnwfsKqeUedntnTgAjW+8wDgu86wRWQIoa7wVLQr
90bobMhHVbG/K3sGIgdYU9Fq4+9VWQXoOb4CNGaBPuFBU2rpl+a6FVZY17jUgOQ2
/wKxCcrPG5MhiolBBPZR+SWpwFM9obakLXK6o4MN2DHIwDIw6MfiQky8QofXHrhi
s48cIltdBU0YvO7dQOBnbxHR5TnNtYtZ1MxHuTs+Mwek4EizbfIWqanYyUwBg/kM
xgtnfhmhs+HW9+uP1ZzT9HlzQWuV6fllzNLbjpN7wUC+xDFdTgJyRVajupP9tT7p
kLoWgBbwGNi+rO+PmGEZ2o/BIvBx4wSWnEAZl93MCP9UYKQLKwkTUaBy+2yVMWNm
jUZGTnPtLNc5TlixHJZagFo9loiBuFDWZxE8r/7fXSOgIvzboab2qWshQR+Y/f6I
/WT2LcklDiqLpu9BD8CQJ7z3aP5WuAsnYJv1wt/+6FldI717zYtgLrcJWrkPX9iS
HScXg4fTqTJh+SeSb4CefxdzIomHRZ7fT3gFJhE1wJHig7WFu7lwL7t9tsLuDviw
uFECIShR8IX1seV7bplUGga1xS+ueKA2CXxglJOsVkFgOmuq4d4iHXcR52xYROmg
7d1Wf+eWvAiUmp05m38r+OtSBMYTpQl2UIx77vh9T+nD90ls0Gfv7v2894pflktK
6e+CeHUQTljbgfajuIB7TCjb3on/6Kvlln8e7WcAPbYXMCGbkzZqY6WQd/6bEtz5
LzilRGxX091v04NO9X4+pzJkN6sf8MndDgxfa/TRk1lghBrRHoEMNRHF9y18ow0U
6EwEZsC0ZfF8MeUCcJnmYz8Lut1ilvKI4DYrUyT5RbxEy3vZoSiitS/+qyv1n13n
RmdG9S/tuwo4DnsPJkFjBAnFfZOPhQtdPS9WFG8UP04t1E5CTUyAeeFCm3F79kmO
N5ga0crshEnEeUqW/PPLYCNQU5h7tGvJ1ybTLOV//sYXprEp+NR/m8ZbuWg+fxSi
F9moCeWVdQusIRcYpx6L+jRbT7aWn9CfeRGczNCUc59b+4imGoBWCuxHp+nq63AI
aV6Mye283XyTbawhReHegv7hynkNb9JKWR/7pZ2pM3MTRyiYHFH0EhRWtNTAZce2
BnHHevwIHA44qn7bYE7QyBMcWF2gOc2osuGCDoe/i0S7uS4eipv0nKocYeqf4eCu
Fe4xX4pcDNXIun+wB+6PO0WX7zpskxMXEhNZoyIYuLgyo0IoD6+DTX/LoXCvs7KZ
djIS6dfEz827D2jct9I2kGRCV4WVNWKREjzmoVdmhqStsF/FY1TV1skLggcvU724
dCnGXhvfm8K8TFwEfggDQsCJrcyAGfyYw7Gp1nZix9vUft1M4QQblaCo+sDBZfnK
wDV/BVeESp1w63OVfWXiDCvsWECd/kk4tatgBk7O2vsNNL5UkWKB95EMA8Jo+PK2
BJIW7+9dqJQyWVWaQW7ya18RVJaGy9P3CRUrVHCH+ntXRIy/X4BknWbX8nVZlmKl
/r2IxN3jdy2avnytI1Nw78W8giFOSEkruB1KptK5tXkSZu3FtdRnMY4ozmW1bcGZ
MDrS3UbiYL6o9d50RDWn2oM6d+GkkwapvSnedXHnjklHpGngjw0rPXsSm+az/iUf
DhskReCQOiEk7bdfJZRxS26XC2JT8zu0oqz8z8leByVJX8clPL9QwcrdRPGZhwEm
QE1Ri9zj8dIfZMJpB4zKlTZqBuw+WiA/hkgalYE8ziGd7gRKFRSQ+KYuPuxj9t/G
N3ZtFLrN1/P1GakQA00z3ZQQHZF+Fb/1o9RTRlgtfcqLCPvPxhiXNxr7bgGZj483
/IdboCOpcJwlMfHCSDJqxR+8+Oug66P+SUZfCRhaoJeXIf6ZoA7BRUf9JoW2XN+d
BUYO6K0ebj73TKIr1dqkhl0CbyykGLy2a9tSUsBvBrWFUgtqFTMV5ggxF4FJcaxi
kZeQWV2vNr3Q+6RbkHtHqkOwHQiv09+tkuD2nN7veVdCJ64kqQY0f+GHyPjLYfsB
9u6p5w1NfzrMnfivmETYF/MJSH1R6D3+rjRoog1CoIauZd1Dv5HxRwpt7AvDwzHj
OnxgUgDm/ked9RUhMgNb9g+b0FSpfAO0n8N8fPhPEhRXhr4uPXve5X6/RilIYmBs
nU6G49iwrvtdVtpfOF21ZY/maZomNzxVkYeh5FFh+ISvngzUuultd1rLxKUaBds3
Nb8yz9JPEfTVaeoBtZtN9U6VBNmkkzUNAi0RyWIRcaM/aEp398laiPPAthwbE+aZ
vD0V0v5wRNpidvFBQuHE7P5Ta9B0FzakOVNUGQB3TXcMf43pPD2UgUGeTywCLz9j
14vbx9pZi2WhRRAxTpwKvtUdjRZtXnWCCr9rTXAIlbiGJ9fj5NmD4BnpW0kxhuwY
goFls1sc5CuAqOjydrjsAGCkp+W71+5PG0/RCcp/mPWXN8UenOf1BVIbMeP8ctUT
5KNh6BZ0pK8vS2JT3f/5rpOSg+ZcgHEpJtdQfO64dtafRw2Lhz71F6wi371Sf8VI
c960eR9uSQZndM8ozGAJblFsdnluTbxBQDy/tId85+eTnVoBsJ3PBRH1mBhBXHEK
GH2K9mlhyhYuelQqfx+P9Nzhd/TmcvxF+9dz7X1Jyso647cCsCqlJJ53/ERIv2eT
OPXh6PeYghKSwvpWCWLWEfa/bfxqme9B1YEQ6hELj+J6vX56Q3uvtpZFFwu6rh9Z
GHuI/Al9XffbIOoMGsedeAM+y5bD/3I+ny6jjLyGCeeZOAgmJWvgU6T869iyzy57
UV+9QH2CQ3prDCRXUQU6jTe3Icd29YkNqdV3+xk62z9E+DZIuSojPX7dFAC4sze6
F/v7hShzdZ2qpKTVNV6MSUl8bV2+iZd8SfyzUd/a9PBz8WllI6jkrI66iChrNuHl
OWStwDjFnU1mG5Y4lDclgWhsypZzCMr+ZQKQtH1HoQ8dhKEo+ILW71MtehvEVwTA
xsRr4dbh88en/rvEBZp3zg05LPcFE7haxowBor5+e480GnoSdZNaGI8gDg28kYoG
jjrgPDYk76L/aabTCdUFbmflNRMzCDOjvehGAUyYjtQfR9Q3n8R29Nw9nd5ZB/nZ
Y0bifbTRSq4PQmaNIbJZxIFjSlHh7ipjA5wqhSucrLhY+U2oc8OIXwLX83Sgu7QP
qv5YUZm6iFtGBVe0bSx7LlB8YUrZFIaoON2hlZDvkYlWhYiDQ1Z7q9hiBrTlMgPZ
HWMN7i9/EG7HktiivsIU1YcGXM/JAcFSTnlIhK+EYZwnx8oyYz4nuJxGu5GEz/Yk
zetvkyhJVDTo0Z6XQ4DoA8Hd43ZTY4vqvDBOmsvpeTJMBkn5qlzGVSXgeIGasmw1
+wahCFDzvOJBMtUFpE75nR99lDAPXVYGVmNV4lG0BmL4gCJad+/cv/tdDunvnOYM
vMTL106Pe64UkUccmnbX49H0yy3j33kc97Nl132h4RXxfiBTyVNJp2WnSKy9kF6n
U5KzeYD2qN2yQ/irzqhxJJUGCBvZfkUVJcF2oxlm56hJxRMHQVGC6alC5XF0IEop
BmazcYI25ed/S3mfWRiI/FQ6NbN74aLcklZju9m6Ur4b4B3NhOTdWnyblJaq3MKL
2fVFEoeMgLFaYwu2NYCjeYzl0qZjzwwu3u9ZyRskmv1tGeUSq5B//9idP9BRSTxU
5am+iPfOyU7kn0/LhaJzZyMxlDZt4Ed7+9wUhPhGekS99ouUCOuQ3QNIRUZC6oUl
Fr5wnygyQrIsuvFOqvmtP5y8wYbNjBc5GiC8LglcUECy+J9T9KTr6AnapNWOZpCa
MKCsWAbNl/wRIEIga+VNRXaldChjQ88xn1j2tz79zMn7+pxrJRsHrjUa1R1FFwNe
RGswn3PdOS9cPSWBGV+UoZmGzs1b8XpWaH2z+oBTISEiqep1XLtIKqF2fevKWmKn
64FsaF2SFczu1KgrvTSDwrdAqOUlnDYwAbs6EGXDPKOcGc/EHPLRB6DXS8rvBYaK
0dVoZPc33DSWvLWBm8zGcKny1MUOKaYkPh7Cg6VaT28ubtG3mIktRmVISsxpusFX
LTpcA3cxK/g2zCYIcVM4h26fdWvpDNhz7F7rVY4/byJsDNM++GuCkwW2B7NT7G/n
PhTpl5Ymta73wa0rR3KRgVnq62f3oZc/PyF6D6saIztafQ9jFXxvlP4IDipfMJTx
6sKPTL+f15jGWQWeHeyHIakT5ZbmqB+A5RihIgnf5gEdiVXxrwFlqHN24WYKHzAK
pbfSwrct3qEBevcQZ4WpGmVnZj4+TjzzrruFsdSfp7U6nIqVTkYzuZW+HQTU5YHl
Z1xu5grMjQVZKsRI8ZgwDiWcDBVCJbQhQ0+bQh1VXRt3r/CLij4IC59KqSviGBN0
VW7WJk319t/W9+7ElL0vuCFxQgGTSDxv8jlpnCAvorbAb1u6gngEZT3iFj4UyUsK
rZlVc2Ni4tfXMEHmHXTDfjTYyLJqXaLo1nk+bx/0ZU7D2Bij2RfmVQhqYIBOsBxi
u3byXhk2UM9twKKiQrIa2M8KXRYiaF8jVQVJ+GEZ2Ps1MNXdEWCFBBULdIEr+VIA
POMZXbfuucU3+ttbSG89JOOrzfPclsucnL4BuJsq+ZHzz8d3Pw14AcclZobyf7i4
hrOdebpmEeJbD8Ot/EtbAN8IN5X90lDLzRpdoYZ9t9FWbsD5eaOcfsI6zOX+MnDi
izvg0HYjZxoFKl+Im2EdWbxGdTakgW0wOsTJbRDOCZRNcnsNUW1VW1zNthyezsXF
YzHQqRYvUjYSTTpfwMKYs/FnNLY5nSDFV7iEqhqyLNUdrEbwrI7zUSt1xiWTDgCD
MAB/DheNsSgWiyJg9wTSBFhhUFg+CddOzRLC9WSPFEe/qnBQ4tnWL7gqdsBA9yTr
669nmJj/NCsexKO2boRgkV8XCaFE7AI7vuVS5FmkN3hPJ0ppt3NIx0o6AI1jF7s+
Eh/0Uuy73NuXn2wB4Doh7pe4TXpx8H6IgJHG6kUD9LKrEUO2k46XWBdN/6OFMix6
E3gyQVffjycwXyM14pVthNFOr7YbL7qyWVuzKr/Q8Io+MjV71W28qNKlOkCZf+J0
Mn/07gubFOrzcVanG0bSAbpeR16Rrtb1V4OdxnVddM4ada7cBOtF2KfrUGYy+yDX
IgOIVlGE9P+fxfzIjAH8cX+/h/KlpMWjAFDXi5Q51uymbYYpOq1kuVw8nLSuxhPa
GE1/gCeg+mlhYcv5YIsdb+qLcVzgVk0HJVboLGtKUDStE6hukRHuC/8ZCXZFD6/l
A+iOaOGOP7fqcrdDjHKldcm8uyNO0ldaNs2rCj00Ni4ifs+Jy0YLfhn9eGumGyDl
QVzlL3QHJSdmEYfu2UCS4RkQaHZ5e5WHM9vE/eHucNa5BFnyHoW0YmybgOtBQDGF
shbe3u00Nmu4NiiAPpnBkmSElV7sxs4iEv8yxjn336dhDWFiQbsVAsLBmcMkFeKM
3NJeQ0pBGNgrNKkDn9LS9rrLgnKBtXk8OfBtd/InDxDqUgK70NC+OqGU/xtcIBA/
ahCH2dVGpwpxFq9qEJJRvgcjEc88ZQzpTLGW4O0ZlWpQF1+I5PpcT139RarM+xxy
6gPlx1PXMDRpWH+JbRHADuHXYbs2ewgiAQj+T1OZzsg+FtDQMUOj6hZOG+JiP2iu
3OSRMzwM+Xjo8RVVbZDOEG6828DBsApFrD4OwQHgrDe5Vguqd8rs0dv2/DzxzB/Q
nIehp7wSkaVAev+R9IAFwxJXjkYp2ZqLU2YfRJvWpZrWnkCGsudPpQaVJx/PEIbL
C5XmvU7htB4bQCSlsIh0JsoJxjxQeVZC51uz4fYUEbeJWhgms0o67Bz7TOV+U348
7d0C7FjbYTeGnJcGLvlTQBObk1/5oKzayMSzulVE7Nea5SCuJFFSo7fIHvXqItiO
ey+ZC0cnr1RKB1dULbfnIX99k0+OngOl9TtuAb+5ND3Jw2J0JQr4Eqt+ojOzpsUE
MNQSZUbUPM+45j7R2SQePoa4sik0pBmM7zfj0/FrIv5alONiMfMOLfGUg9qNawLV
HCN53Wibu6j8RoP6l4Dv93qOuC+URZeBIFuY9OICrEEhshK4L2n+6r/zDVji3PRc
ZtkTqvaLHxwkuCeOS4ku4GJEP+XSJZbLbwBwrbHas2ZO1crqL75uHVrIdJMwxioU
KUHljqTFWqp8JbWK0bnpsKxztCJW4c3d9/o5AGbJqUyEJFn2W/aG9IeHNHLyJ6kt
NvTp8nHwm6QoWqdHGNBLst8Ld4i3k6GrL7ukvQTiIaj4XgN6pol9FmhRqQ+1PT4J
qQL+tWGh6E1+hJsn+T+PKq6kWqyMIGsjwCrBFZha+3HElXmWqbxNFERge0udeRI9
8eZkQkp8yElFRVboznZAYm37b7PZk+ey98wuDNHIWgAtja/JMcHvRO0VGi5A3piY
t17dStJcW+0srib30ayO5ETQfFPVmOsitYGL580inSEPVdC7YQYR9XnaYHfwF4Bi
sIDrdT9f/0pRMZudwUEjhY7PVnWXln9EtLKj3MA9QsbeFD8Y9YYZ4rtX0OF7q1xm
R5Lp4oi6gXKT0MQdmU0HGA0K2qf2cJY7Z+HAW2cJD2Aa6O8NAR4VZVoGoUcIAmXY
R2/IW712oMN9m0jBVEMFtXtPkCHuEo1nE1EJg5vticLlZMGFHSv+29k3b/UqzZ1Z
WbCVIKGU48vv0YHY1KKDutekUHPbE1GLe0XU2qFwWsM3IuytMExEqLuvXaMQBh/x
svPOxJDYktzoHS70i2wHxsyh+sgQBD0HrRK4M29Z758m3nvdVr7TifINovmYWbUq
l2Py5cqs1E/Xczepch6qIATixwJOiYIC/50+TbZ/wi9gxw+rQ0UYa5A3fgPKmmBh
tP34zEwadoP3uciYlVmEbGSFM68Uf6O/RVPd34taZYi4hRrd8Fd15o82T9QnL098
UpRKtpbsPIcu0axeQxMF/6oDOeF6VAazvS7ziVu3dAh8UE7ShKlBy/OFV0vL+RIu
KonFlNt/GsZnW38qduXJT+NPs/bj9Gveu2KqK1biPC2LBnNni2VCTv/itc8NLWQw
u4KdRRRg64NUKTxVF+XNFW+7RaAkUzrn1KjUu4e5Rc6ZbpQlvnj8fkwQ+1A+IlPO
nl2JOny76f6KwmWScPU2x27g2L8G+4UnzK59L3i/sdj8z10H9mW6axqmtwIIQuy2
/M5kshdkVcnxt/0okjoLw9t14+8a6s2CrMPQ4oHzh6U/sZy3bmOyDkFa1gW3L1aW
ao5wkXmOTx1ZH30l/FxbiS1+DqYABNnrEegRaYHvf8r227GuVNOK7rcYmFjf5YOD
bkKMBIdS1Ry58zKVqbFXWNLLpLuFlhaYJuumCA9TFrtDqBg1jpCdRA2eJL2Stxt3
msJ5n9a7C7YXsBbhGXbbX+8PHjYQOXT5havZvwpuA/0zg397cU+YBadSUFufZ5VB
vkbVaFRDUE1Bd0bq0uLldLnycxAeXw3cWcGKyemnqsrKNvF4tA0NNGmZmIrBdm1i
dWSiBK3AtMKrB7LtOZ3K8aT9U46GKbAVbakk203ab+uDMJzh6G3A64cnAFUzq80s
BTQUFqv5Nyg8s9PXvTYNxKLZzaEL4HG4iPT87yTpRN2lvVrn+QNeGualcGZSv1Oy
xDaOL6mDX+qbOhSVB14/L+pGDWNsXRw8uaeeCt74dd+5msHdloNG4PDHg39mcmLe
KIY9O4SjnoFZ+mbTxNc7r7nfOyIDSt4CoE3Yp0s8PHAgE9hjFLCfRaxjfuSa0CGU
eGRkfndEH+v+xEZzBNDoeRT4F6gsLQwCCS1xdnjI8gdj86Z1mJ/q44zLUAAmnMBZ
SK0cL/6MaSIJs5ONa8cqbJ6PqktCoIlCEhfnmjjf8kfGlwmr/R9zhzI8l4bNYxrj
T5zN4IYYTgVK7pLBn/d617sVVDAcFKbZ3uCvjrEjJd8oA4HpHr2uKqoN2SB7w2wp
NwgeghMStkGBLvWz6gOpcvopPqhnJ8Gs/A+HlUvKsZiiVNp5uOLHcCNGH5upZZ1i
lpl0Xxp7HxOfUti+PfuNREPw4mT+pfeX0sGUTyAnoRvVVsiVA4NuUdXTT3TVeuRA
iArktduQXTAYLvd9GQ4nO0ltoJsvbEZ1TQRhieo95hFUfhLsVZ5nYV4iV2ggu1Qf
vgWmEDeSvdoxr2XjIBljD8Ao9uPhE/yYN7X10xQ/OQvU8y7b06PSG6zYWY3IWFwc
YNgqDvaG8ysW7eBKoQKoE94x8i9H6xDNo2RPUeyWlCc9uzmveWUrcEGKRzEmioPs
4FUsmqdXhWhaelJKoa+lDMePtMDLarUdDorkE8VNcELTP1ueMYiSsx41k4dVCbdJ
25M9yRfpaVYYQ40h58p5LfhyiLfIrFV2IgI2ZswQki5mChY7hm4cwInDXasZaf7w
+Zj+0URdc6ZmTNqc07bwPexS0owT4uQV2FYHQKe3okmLZC1DCSZmQknXZi8pif8l
/7hzZQ3Qal1yPfHTJ29rpXqeb2NqUkeUdtcf/eA+mwlB1WHEh5yoZFFsoPDe1oS9
WY/suYer9QZ8t8+Tkz5MAg8uy6982c/ugo0sYNFQdyOOtO/WpblVT88R9qykSEF+
QDiBmQ2xuwwl7ZTTKD+sscTdnrIX4kjgNaxDKnJ833UU9Exg0iycgk/6FRbO3fRc
SLbd4mXKgl1vfct5PScb4GUpAN3T3eGEnYt7Q2DPrDxOpYKGBSfPPkVu7TJVO8kq
ReLBFdUcBy6vHGqWBWbq2QTx357s0V2QfP6Y4yMz1+txB83q0hB0m8Hp96SHXe0A
Eca3CbobzutlA1mTg73gdaQARfehjxG4rimsm0xExX0ZqpKNuAGsTHdXdk9T/fT5
OT7vkygN+++SwkfneOwAH3OjQbcLUkWCuiXYDoUmgKYjneTikHMe0kVRBthRx0SV
sbCreML8+4UXHkI+Zq0O6aaQJvVV+o0BwfUjEpwtFUhT7CO9oXOaMl29QbsZ8dss
ZVicPq6O2QCg0MFX4ZgM6Igwvbbba8Kaj97jXeyv7KR1KcVCQEAb7hASJon9QetM
P2IaLMTx6nvGIRsJ6sI99Ieen6mZWKIsfGQKqIqlCsklM8Toy1PaKgQAoPsKdHjo
qO7oRyJh6usR5K4QrKNnSyyqgFPU93LsbyIQxnOP/rPCKtjpYL7zBe5OlqDdxQQS
Hm5iPvpvDuJbqVV6ZbR3hkdHdC/c/mv6JjXIGy91H7ZTqD+bG3ImmXExaNK+k51W
8VOTTyN7s2iMOvwZWRmj7uFnqK51TmZDm5uz1LOPIBv6fW5DImMSMMK/jkZwZZ6v
oo4BN2PeyvkFPNbugIXQx/JDSicwNEh27fpANwiUDu93/hvtN0uHiiEat4wvP78j
KF9lm+tt6pILppfzF3YhYptpm8Ob24XHH+h6SrzWkOsqX0zeFIiz2kTdjyyTZqCW
8Ysma363xmmwbpNK1UTleXH6eQboOMplksm/inE2hS6YB8RNiI6GoNXGtE0RZZqm
Gl15eRMamUwfNy1mI3VkKzrzljnBCn/lOBaYBfz8lNt53PQ9Cda2xXjAZ3H5jf2u
tQ3BvGXvIk6d88UEz/cAQbEUGHbH0EanN6R15ypPkCrUB3Mi9qsdEhIZ2+XdHH3e
fGmG0Rxv0jsIXlyC2xsRZ9rHpCWCNwO3mIsqGw2QBUcInuVPQ9KORa5/fihLisuR
OXxOYCju/0D7Aqza0pUFq5+q7dJ1lqeov0xcE/BGkXaaTwD7/9V1dA9v3TRSeXEt
oe0VLLiTWP7I1KE2uLKGCmdZC8ZIpNZyTr/UV1zVls6fC6vhY00iNeNTIP50lIrV
QSHNbHTzvwe9pKflD1VCidZ5acbgWjvwiXiZzfYVLpWvByPLvBZtfTokGkf7KfyZ
nK52DmIlqXCgnYvof1qZ6mwjcGZBaykoAyO6V0PO4xZFsmMbbY9pD1XbDShtiTb5
Q90XT2kDMXZUDw8kxiSsSyTyDrzo/au747A5ne09b1mqwHbFNNiphzRxgZeTWUsN
Qs8yIbUZ1iMuyPp/bpcgg/SocxuLbPIAd3mm7SrG2JaRxtFAUCCU2yzZeCdF1a9Q
4+SyO7R7Bmr2wgJc/vYiH5hNajI3606f8alahamcBKuVYbeT1rQAPNIr7h4KSUrr
HIc8aIcguzlcVrQVrMIE3S+yCBHQ+sfwAQcfFSB0GuhwVGw0RB1URipFnUnCiY+/
3JVIxVF9396CCSlUA2tYpOeyfPBvnFBkiv2lAfxXAGUh1o5ta39Y8ZqqYztl581n
VMwC7o/mAlDf1DCxX0/tu4SFIDVkrgcvhq+ZAqsRUEUgBq4eU0XxXu3aFWIVJiEf
OXXq/Bm7d+I+3sAx7z0b7ALSjQ1gA5IikDgnsw5Yx/IJxTk7QDnQkz0ZUhR1B8YS
WvSJzn+t4czMksvjo4cgloA2tuaHkndtGlGUeEN3myrG9ofDAkqTLRuNY0bPANrZ
kbMdhUUltKpMVEj3dGzLyBC6uk0tSZ/PN2SeHhAwheSoWt5Rtv50jexYo9fobrK4
AKeI7VjqIF+d8bSViFc45MN681AVndclK6PJFv6l0CZrQLTn38oxc1ogDuDAsVzZ
DPJk3lWvxWq/hSpM3JxianNh16Vdi41C3asDFWxcMvNMYvST2j4ClVT8Dautxnew
0arfR0+mzog8VHUKFcr1eJ6MA4GoIuNiw6PsLufcCMQucHwRurk0BsWS/AD3eN6A
A2R6FFeVaORQQFeiADtNpNWA90LuG6ehsUa5M7Ec8PZ3gKa5Tah6KN3m/FcSoG52
LHaBLHLaQfaOFgmNdimNfhD2frdiboE3q7Zd9RNzuuw=
`pragma protect end_protected
