// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bb4vjNd3OgWwnVkYAoA6EuYiVPzx70U6xTpY8Nyn6kY7XbIXqDrwZORMCWCGQBbR
jrtKeErRgM7TKfc2Ff/9YWRS1dMf9id3NqvK/J9Dzuw3/iPI3Z1JQDoP+ENijOW8
AIGMvooquEKSxle2ri+7C52/1jBtGhJfVMT+C8Nnn10=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2704)
32R/0ckMkUsGWD7lG7HhUK1gCVkneogYzxeb4eX6Pf5FUBeNc7eg5RyHLrxmaqSi
KvbWqoExZ+rPk55nL8wCW2GBUcolYZF4Zm2vxTEL/wxg9qArvprZtHXT6/w2WZAF
FLMU/fQeGecU46rqCD0CWuiMUMWy6UTy1arQbb2gKqgkRUM9Qf5wCAsrm885yQN/
MbXaPkmSRohfbLf/DUdg/Donum7UvpaBD1OXJqsocA/3XSRkG+GMAfUDZDRbMDbO
TNpwBh0uFnVPIV0spjg4QHXMwurzZvpCw81G6zOMVU0tO45GNoQuPdufdaA5JfoA
b7u8EUDzoueVLiwJzXw20vECcTAWmNMAtSclHcXXi3ZN2fvoTIlTB47kirODrtVK
BnpsfIqBn4FrDEY8If2Vi/lZ8IwTqELCoI2vx4GB/w5G/HavCVRldqw6kweyJ+dc
FTwctZuZL2TsSi4Es/YwiSBMwh2mauKN6Oa9O0Vpsm2URz93H/VMntcm+wqCzVJI
nwNAQk37v7ZZ9D9pF3EI5Tc0wYMCdkMovMxbEfgU6mI/0C0qEAe7Fnx6BcyfeNTk
WLeYiOb3Inzqvnytb6+Qc8hHt/kt97QL6qXlKxM0tZtxcNGt+CZ49x9r+1dhvGkS
eotP9H3y1jF9M1i/yKogRV5zUVR6ezvz5QDcOuSO34wKdziM7JGSUgLEil7MhEH/
4u9edBCB4YHRtMnTlxl1h+MZSwbvvONOXpzylFgWQfv8FdzOvUPww76d6vsYiy0i
MF+hodM1HE9EIqd5AKLC5C1DMmGN3iGs63kwgvkqC7URkog9HlxTslUaUkwQTsYd
0G/6naWoI06fLFiz3KPn11oQGzo579dr1BItePLphrXc6+E+W7Yl1YGNaajXRgAp
ktQq99D+0AJziZR44IKIfhS8lVi2RSBF/svoE54QS2qnmnDx9ER0WXhxRXvschxO
lmFOB4xR50k3rkTLAd5BItxKUx6cAOJtqASa/FbFQCNh9GrLzdfs2ltZHCpLRKBX
m6F13PpQ4cPyvuYrhJE+0qc/DLUWthiwu+jeKFFoJoqDYWSZtWIvsMvwoV3sJHar
KYRQbbycZOKpBDoyL8rHYiPl1EoeEAJs6PW6KPUHzhVyj91GknWSDsNXrgiUDPNv
Z8E7eg2vBb4K+LOwsMQkMl2c9wGM+k/ALo/ydFXEnzQd5iRXbWSGVOnMbo+zcJXA
VeFJX5ytFb2QneuM/uN4Yx3v7sXVZTKZRmU0KT1Lkivj+mtco09WUR74wiW2JrTo
LvaIU+qeUmGCH/EsFCAfuQlkvZ6HDKgMQdp7NW7EbKWn/XdYfSz6gSyBTgoPu21T
B7fOboRo/GiZhKHd9dXcnb8BWp4TgVPZAID/2bdPzcnMVcOpx/yxRsShJaQtBpIr
HAbJnNWm7S6jrf/hIBIPwO0LDVNNxpQRIFbvOOJS4Z+qcwcs3qy5nmQsFRzEnCYh
EMNdN/9/9C+B0aRgjuAyfmCUcSdTCk6uSb5Zs7A2H53fQwrRPR5t6JCAjIAsYcSk
RK9uCrbWALAwjlx3vvcVO6ZfCgVd15R6CgpU4beqoHx5Zo8hKxlYPVhZbVDjj1Hp
nK9uBJ2OnQ2V170z31/iWDDnUj6LlsCuePJR5BNps8k7eLr1imYpldFjE1L1/Ssb
/C6BNHU4e+tYtFG+JLRsSDUZEhJKgQUoa5vGUmwLX5ErX2moz3FqJp6Ur1A0ZpNC
VTDfM4h7okabVj6UcvjRb1vnohDMA4UuS1wfk540ZrnlvHfkajffKUIaiRxcnloY
cV92OvMs1lyfF/jVLKiEXaXcj55mXUPZqe72NYf63KFI56Ym0PwUYw75ThfREXWX
tXFLnSOx8kVHf1n+JnYGdbgj6AGF6Sui7yqA0XF2NHF6Vv7k4rsKxwbUrBPesoOG
OFaBxwkkr5qrE12TaEOOn2fgDx0VfEfTz477+jSvdQ6R3feeGT/JpQwSp0sMNw96
7nihYAxhePOACfs6k7mQu/dyuyrpKe5olZpM/5301ZlIwyMdNGX2iJpdXi9fUfim
yfLOcd0B2dv7DdmT0oARObhOEFcmiNKJttNzbAhQO/vkJP8zX/gv/iXO3uOYSklO
NEfQjqCCJSd2VnKmCpxMmfaIeuExfBqfcRHcjeNh7wEKCyfR+aQsMKkbjsF8Px4F
HUFBbfbHpCfygTBLdO9FtywtcZyazytP6doSyi2wW71oAmceeUiGAyq9DilT56NR
iqTonJRTjG4cSoXK0dHiRLPak+IB6h1zOeGx57VfvvNng78PAr9KTtYib/CAFBmq
aNuAau/+VlMi3RA6O0+Pd6xcAkmsajaU1oK8k1cE4Les1FBqK+nClLTL0eLcaclb
JXvIq2Um2WdZ5/O21w+eC7JxWEMExnPxUK76mjyITzJWioVxHrdIuauOw25OSBFf
GDdIQMqy2u3HFR91zzA5e9drLbmITbDIVGCTcOT39UzqyK1wna16gcf8Vu1VNknD
ALdKIwfHjaLeWnxZaKD/eSkUwNYxNQzAg/Pjk5BXyLuzfNKGdgw4d6qPRlZ0ACZt
8YLzhUWrZ0m+WEQF8AinK2QwX8/f1eiUOAfoBReRf8ayfClusNAQS4yjr8WFTwaq
TYCg9zs3MaVtFyyi2hRnn5UOKu8Zd6TMPKJUrX5K0QMAV79UgJ2VrVcCrmZWIzT3
fmnMN3jdVq7kUNTujTYmHnBaUN3PZkQXTu75Xsfsij5gjf3GOgnXoTQjtIz9Ecsw
7K9pBu3gnH1E5c/TR8dODCfJitWOY7aTomP5b8dmNBgJrVHthf6vIKuy3d7iSvkt
ljrNEBLvx8WKFsg8n/9qWp58WYbkE0SMLEm4f9BuDrZw9e4PkprqfnyXGaiBnBmb
OgpoM2gVjOeIoervPAe9IhHwDR83JA6s3giEFKGLhN/2tcKsVM56wAtSVX7kPdft
grxl8iRhC1vNkivpfsApzh8zaql1hgNFiADAKC8yYX5V1C3ZHlUyIEmntB/GM3rA
Y24+wbkqIY4MRPFbXY/rmSTEOgGhWaNvXTk4Z4KLPh+3bQ0F3v8v1LlrE85YZoNe
Jk5uUJe8/poeuz3pUkspYodAfdUL9PXNGNdPWQvwJRaOi/gB4WFercjrfok2JRON
TH4aMVqqTHp+ctpWqo+gpN434fX4SVMf6Y48HDsYkstJ/ehvmht+9xLFzA7qLZgA
98lS4dfU23VzUsUUzhjeBw2dMsnCxrNnHGsEapCBurMW3KshMQaHjnfFtke8sgea
dCFnfJvzm3Fk9GtR2aGaCQRsBnF3knFe7M+hnHfNNoHz+tQpjoxgQFxv86lZzl30
p2rrC1GV9NXWaPJiMq5Paza3cI7RaLMdqT7ImZRGf+Sk2A7o8CcChbpC8dC4q6KF
qkmA5JrdD8N/LW4HpxYTFaUm60FSdBb5C1B+B6yPgODZizSWPGdSyIvWps9Hywfr
cNhnY2WV1Xo3FLMgZNU1+95Q1GRhzAadziuXNk1ndJ3h0UXBJrw8dboYTIvyW9xo
q8FLlUMRw8ij5bPKvTKNbD2RGcaz1lT+2J7s2VOjmaCu3NWB3rKOsBD3Lhoxs4Ie
AZKskZ2x93ADHg4aCPSNnA==
`pragma protect end_protected
