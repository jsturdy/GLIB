// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XiMZdFOhVQv4I0LQBmvqH7d4FNqBtVNwYUFrhaGkBk2Q796yqSm1UfKddL4aeye3
z6/RGrcVBO/4C6l+CzJjSS+VlgdA8MRXOwkvCKM00+ZNsnSWNeDJPYeCn6S0vbox
rijqVLhRoW+Wgi9OuPzwdMvSFLIhf/GVJuUboJjfTAQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1952)
EPrrJYgldeqy1bjr5wM9I0nEAn4oXjHYhoXCxR1Hf6Su2aJObSz++e6YQQbjBGRn
dLOtmgFG2PVidZ3DZ3O5SsejRcmPZumcnEHG7t1kxDfaKLye4wk9wuqChtcW4xdp
Bgh112I7k/+FbHBR8yT1Al5VDPCmh4qe/s4XQtFk0zspOswQGgH23TZfM6rPFb0s
s/o2aywNjfXOvfMBaxKhgKv4gVOqigvq6sflZs2IWkPFSrgggvJA3oQXVRMwJHuG
CasUCszUbWFI76uBiVvU2Al3viLWYnFWGh9jClht7qfFexdmwhS2qN5g57am72/j
0W4ATeVfGwiVYR79Eunp3K7rnWmxQqLtgLbEhxjmdZ4JW5dw/ca8DQbipCSNXKpz
gNC0Z+VNU0VUrvtJSZRc3LUsT11uIep0sIRKszr6HNv4gZYZ8A/7RcLOvzqU48tx
307jUxIYfbjQZesBXASFeCc9AcEhC6LJDCQ9xUgIovJ4TTqDESWze98FKg5RGr95
fsuRFAXaH+za2pN5yf8hG56iW5ZF/Si0b3JQqVgPpz5PuBTwvu8z1mxZ/YdNMrDL
QeU6EBbdmTF+/ku18augE6SO9+Ah6s9x95nbGkpCcWV3DHwzh2TT+ddojwvTY6KP
96PEA5+H5ZliH0kWW/h8oEWODlfhTxawGd7S+1T9PaXZRZ8gKKuY1e+vgogAN2od
iV2DSzZSqVrjV8YExpfVewiTWm8yjUyM2nHiS0yMfg93z9Nd+kQ+Epxs5a68EBzj
iIW6ZYX9bZLt+7cWp4dypL7p5sEeEgH57nZ5nijVaOarvJXkSz+0skIpGR39rgAS
ROkq0NeZnnOLzN9e448e1eBPvDvE7hpOFxk+YzobbK65ESU0pXeEDi4ZJZDaQW8N
JMQ/4ZJ+aKFjEbLakgmqPmIzOrxfzOWGuYSzrRifBnj+Pi5p03en9ceEWp1QQEtS
Ev4dl2OFFrdz1XROVlJiEU4wz0pLN5gK+2ZK0F5yCaC0ZzTgRaJ7RA2kM20sats2
eoQntNrVpn3RFzAMXQUzMdgoeSSBQL7kLeN6h7aGSEAkBIyc9Txe5E4D6XEk08M3
b0/CGCd25We7pvDBRf+3xuAtvJTsQ0iac/muBn6+XfymXCQMG04+nzMJHqsLiJ3z
JGJczVgAe6uS+DvG3nfvqe9zfkHD2iWncTa0HW/1wqOKgzdLURkYEBf2T7nHYjSB
AlTZL7kapNDjCVwE9Y+ZQTQ64ziQdrnGt0HoaSrjsxij13gCjvyzpyO9nYz/obip
sCj007efZxnesBMbyxcfwkxBETvoLJiDoa6wKEheLEBnShBLF++q+QZ6xQXm+oSb
4fuyMEOk3j2aDucCHCLdaGSUSq7WGJJcs+3xWsItb0PHeirzZ4JJM9IEf79hGgxG
Kk+c2ZSyEEycpsppKW5vueRsGYQrg54WuOr1UyREtpS8xa7SNMSs7LAMA+uGwzV5
sQl3YUokEAEJSrtf67XdNJHpoEQlh8pfW5POKMxdDw6jHaQU0SH2NoH5Msr6nwTT
d+Bcn6r9wJ8aV9TKrp5xvoYXF/4qy+rN78K5C6/Pm+8fcnEulLhEQCbfsIa6StvM
GC6op/3sxo6+kbEX6OQ+tTC/lQPly/h8jfTFSLKs6Q3lbzMOuVEtbciScfG4Hzkp
vPOR074I150ho4qkbptD0QcE2fuAToLqfOOJsUrnaqO3ir0NpYxb63OvSmUuv1+A
xw/eZXMMxj9df5uKKNZZeqgik7k9UEWqX0jM9Px7TXd+QtEZ6S9NU54I9pbbvw+Y
ePfWDyxWFOFcEKl9YCabf/zHfdMd5dWfkcoxgO8gSrXmU6MLVJjSNLACrwsRGBAO
hxW00FY8BMZZmJ5bZBi0S2mrzxsPai4f/nRZ80iuuKoXqS84ofeXAZtbNZFvr20x
0FthIsIXO7WwLgpw95z+VtWbYLnRTGmpojGrdDnpYVHBMQkYTJJOW8lKdNZNkqXZ
XQOot48DkrlDbWeurhfIgt8u+AyuT3E7GdQE18b9KyXw94lACmeLMjsXo4K1teW7
YbanElk7oTrXN9B4V8QVhicE3FapCzfM4SCaAZYArK/js5BzcPsx9mv9knmmDpU2
bsvOmb47Z5nER0Whox8P3Kt2XyCHHFqEMpgUSggSWIFC8nIhiSNR4jqQBWk9WDPM
XDoSkNkfGTfaDzdAbS5+YoDBfmGhisJIyf3IkmeJRC6//ojWzo+6EtPWpfsRGn8h
UnCBdi15XQnspNQ+v5KqJAQLx0bgkjQtnX35+Wr6VHdYdDD52f5PSk1FzjejZedt
pg2OWHdFoIUDot66pU3KejD4C9xEMotPZ8q/up6WLl7H7AIQuLwGFmGVDiGdUnqi
v5DV5SHVFLhtE6jNgZ0uFV7ltFCNURKRAZgphllmV/yrzUKTladO5whDx9vh4oBl
NrVho07gBwx7Lr4jmVhG/R88Cr8X5ucuPDxHzY+uOby5P4sPRokHdkyMPGqJs7+B
JE30efjnl8slWCVnI15ewt5LKh+qzSI6pwqc+xsVw4jwrd1FFroDTZBl02e6qw6V
hd4kOjyhV6mDfOA2fPN28nXVzUOjSBR8Vvot5r/GmfI=
`pragma protect end_protected
