// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:09 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jUybG69EuUiIXd5a983Dws/Nfn+abivpZr8qscTZB/6F+lFDolZMfra19/5q6szh
hDSUwA+gYcO+dtwlxSeNvkHNHHbay2axPIMY/6nt9mqnGYJ8nXvbTZh8CXhw9LKn
i8YOD4hZ05u5GDdQZPRn0kgLKupcH6TYCz5IpYSc5z4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6336)
nwtu/3o9LW7y2TXBsZap0AcCh2nfUNHbYWEstSD0NmwqzPv97TSCcIbpr498DAUK
+hyo3GAKDOBa/mZIJwgnqxBZjXobDaLK9xmWmKDOaL2Cw+YkTS7Lz/WjuxpADkWQ
y/9TasQv+I0qBrEZghdiJ0de+ShjWKcR/luWDJ4Wc0dL3NAkONq7lFVLepbVb+n3
4PudJ+ociquyMOl+aYhDHGc6lF+vQBPoUOhNizwDBYaVttg1GsFDoF1cDKxL45Cq
dGuFmngb8wcuLGTQJSI6K3eIcijRlg7fr0wFkvh2Fp9waywBVwrOf3AaMBqxcGGp
5G67qTJ8Q4MSKWHN3577yEiVJDotXqxVQP/niU8vd4c+Jz7Fq2x0wbnBGoK32aQ/
0Pq5OF8b6qXsXRhkjmuJWypoxPW3pXOsiMR/cDShGqdzYy7b3HKqQFoP+Hfg8bA3
gcx7gi/msz5A24LymWFwTm9xKoetVhetHmHgbMmQrugiiSOJUbeAhCm/TjN1v5Eq
wRwnjfLiwV+yu2bSW0tqxEu1BupNFk2faMfYCBbpZtHZUpWOiLxBWpmqwSl/WaQK
dYqMfLLlfmDaEX2181UHz0Vbo2LPeiut2nDlw3VmVAVkwuWyknED/Q0APTD+3nxB
g6IayaSaX2qfxc5kEvha+/zlYm9J8pmW81qBiRgvzUjJTil9Im/6M/zORuyo3KjY
S8bcbuJp2VVUFxOoYyfWzGqwWfplEQiXNpIq3laNQDnqFeMWB01OD2M0chEML3Gf
RROPGtTemH02TL4npdlp9zbulkd2kkHnjaT2d9WC56rSkZebCnQuqS/hVEEWzKMV
Ex9cWMEfGZRMBSohi4kIzYGvLV8wcPiXRMOA1bjRLSChI4/FpbHlIbdPVdYwVbS3
kXGLpWzBH12blg3ygkkZQTXAssB1GW70LnsYSbehyNh6XD9wKq8B4QebCYOa20RE
Ze7GqvQ8XWHUhDwutwWofMOuNT46RAXQiEgyxbCJNNPPuxpMkYWpQBpviO/rxpSI
3DUclE++LiB6GKQEv1qZ/vu3/mqg/gjCYlf+f3hernGYX3Sz+Kt2Q2k2T4NNCuSs
kzART9SD5G3zRQzcyC0xx073Lrn7JPU6evGgAL/wBUqGh+fUqphSr9ZYCndz6/LM
eKTARIDyHe8ZvMdRfJH36s2m+fLu2U22bfWYNZeQdO+Cb7mAkwemDrKtOnqJlWQV
y/g21iLp6Va5btpc7dwF0ti7dl1FeBg3/lGXr+CLSOcXb1vFnVI6ZatjuBS0Bgzd
h2tmADx/0ervSIeQJpj5IPJlWSuh3gIVO1WknnxqcQ7PQDSF4ECa//AlVm+VDxUq
M7qBX4yfQglRSp6LZ/6eJyLV6asKFCJ5+xkCJ7Rs1HlyUskUQ/Vbdlk2WXHDGnOH
oBRI7j3WJy2HdfP5Jjmfa54g6HENGrM+Z7/7meXIHRcBhCWfZG3pqSkF2tnkCVPu
hd9JCarl6p2smGng/sMmTIpzpkLDWjtniv/mLbiYMrk9iskOI3byLE88A6oDX4QU
FirpI61OiL8xhjzzXkToRjOl/IgZO+KTGam7vhzUmgdtwGLhJmnH8PJjs4FRk+wb
LIf+2h2FXH2G0VJyr+RRJBOtyBj1ncT1uub4C7lkF/U63HAgrPJDlVtNLf3/9snN
90KpsYlW/qmSfJMlk/W5X2S5RLe5ad5hZ8pNvI06hFzafY6queHuoku8NYcEXED2
wUob/YTvYyUanTk6vlBhBpV1zEi6KHMN2vQ7e5IrmCEBtuSx59XrEChxApuXqw6n
bLnj1OkFQWsZ7dFCY0SxWaxfgzEAN2w+W69ABmcHsIc9LJ5ZNIXdQn0FFfPaFy7/
l7TXjpUU7XQLWxSnxGQhEkUsCi6Tg1g48u3w9NNoE1fSziPN7kmaGBHaXBCMlnn+
E0VLADpXRoT9ChDHad23W40BawWECAjLLBIKQzmoMmBwGdXBfhwO6F8XohXVkYaD
8jEbnrXs2CgLJlbaEum3ZMuw1po9G1enOWnDrwFByxGglRBu6C7ShjC0YYf/PEMK
Ef/tx/MHsHeLWMxKYiN8PlSJF8Ihzr1qLrzMSy+uEpOOzcQyCEacyvdD+P9z/xbx
D9ZgTgJ+itx4s3e1IEuP5FtNwxjJSQN+Pflhqh6dS1MkMlC7ADE1eI7Xr/N8FzD8
Z3dh6OvhOHLDEUPb1HbxMvatxjt8vUd9uR2AYJrXxdx5+5Dt+p52zE1u0RP+Sg0X
8m0iZLoH48aVN0BnjpcyN5DVTA4GiAiunn8TtVUnL47skneF7EmX+EJPXWFMNU8S
0oERLY42q4kJR5+6EWkBgXvXJ/NvU+5eOxEsfZY0Q0Uiq4t87+5AiBiWVt/Ky0Mn
wNtWsJuXa6hdhKfafVSXjYOno91gdRLQKn92ncVkNRIm5m9uXvtAyc53a5znHxNH
cC6OzarzjawXlk1Tx5ZAsAEhS8t0UmOzOB+97eqRLvC6Q/+CQ406j1YEPCyYvxJg
EPrvJRkIy9wNnSgK6YERsN+alpP5pBC1TgRFrNJ4oDWFDCaQAQxMCpiU7Kd8v0a0
+72HWv5eXQL56axsoMEd7J+o+nGHyieKicxniFJKgRnRoNXDxGa6ChgGaaaZ0tGh
fiHAUiZTOD4N7+Niy5GhNgNfZ1IMkgAC6AESNjaowFjnroybpBDo0r/MsrQ4XU5m
ZnIrrsY2z4qPVS+9MxpW+f6M1f9wFbjqeMR5kh/gEq9X75LVO7/Rf7/J58LLZJDR
Wsdaw3Av+bfYu8vy7tkaNIkN5iSyn6RGF+6cdomfp/CITZuSzr9KmkThuEx84hqu
fCAb7IHzG5GxdekOGdhnTFKr6p9LqOsbcOfUMRfaEb/EY1+jzDRns6HgKWMRLOXT
/1t32oY+cs7jjN4eRj3xiJNheiq7+00oQ0Z6OghcgVgdbdQBctxBXsuPFxbSivDy
gltp0X2FbellzGH7eBpH6AnZ4PBSjzxTF/9bZKFWkdc8/vjNlmWAn/+phvasm8AS
ISAknVlg4i8FWJwRCzKwnj2jh0HveiXzG6dpc8HffpHXrQI/eZ8BqKBnLCdlDmAW
2aHvAmGRZl47asN1QRKfmnD+Q5R9XWwDjbvnraHfIYo7RgY80V1qERr3ZFPRKz1f
JRUdUuXn4tllG39hrd6Vhr4hDFWBBFtFGgAJU7v70QBn0vbTT6ERYJZgeW0eTVcy
T4BHkX2fcQ+b4oXCRGVdN6Q4KjD4G1BiZIf2Nbcgzi1ct+IDSvv2H8lNelagVyrB
tAInwikLAJTr0ZtFMq+Pyv1frtgHsgAyziUAaRiJzt/6+irMEbLlk8/hha3vOWhm
1FKmYO2bohjpbcIsnAAUdqQvfX9fd/Y92tbHL/gE3/P6fNTjrhfaU9DZ51NN+vqo
6rxTOXIzZy7q9EJBOFZCz0ibTP1R2OQ9Edb6/9L3M9/P9gEbogreNhcx32srl8dv
RoA7/QdLZcrLht8DWnhDpjjMhdQ26m5yPYq7uQ8MpyWWuR5ah1//YWhKWvy4w8TR
/vudnrqtxQRFLRemE5g3dllyL43wkHXLB/jOjUx67RMMFFGdYoMlxih1dxtrAN0U
zpBOC/weHv3qj7NDyPkrtif0+vJUz5kE5AXE8mUOq0HS6blEkUbj/PRfMOk6oD19
z3knass3n/AgXvXBRbm5vYTewhiYA28Zk68TdLj3CCXNrS66HPwef/9/KTdMGKue
rqGV6W9Q+kPfFVNVki19Z4RNZmXyn2SI9u/miWZtLaoUN57A4dKRDV6AlkRJ6q51
QFRlrZXOh9T+idBA70GjFrjEokWW1Wq4bR5iCB223DzeHMHCQDQignObRIhtj9nc
KL87nST0jIdi95fvtBnS1Lpc2umxMB4n8fUOMYv2a2ok1rkbLqPOOMr8PvAYfsJ7
Ug5LFnuAjOY41HAmXYwS416bKlv8vv77/bjniuPgAuCH3KUVenL9qYgKCJM8juD4
aqqGNlMTYsPyvuPLmHgdoWsjOyaRSxfRi3pKcRKmIYy/kJpPjQ8pWa8ZzOBy7NIm
chJduJOPGSKW34bJL4Af313Kag2ZqJyYepic0bV3zN1Qh7sqDKaxvTukfurIBTu1
vpObqP3GAmdbazfGYZq5DKbJsRlMafknfGc3wp1tao/blRA6E0Y4yKWcWm5DPsiE
keNyHARM4lFXDtOP1gGDs0Udn8fGkSeDmtci+cpFS1xAH81TI4eUoELDI8B7FuEx
qblRNDPyCBWPqpS/yv+Qc6SMP83YfxWGuoqbli7IeX6eswgpOEdimQxYKBhQEZnQ
VlW/wS/29eXbWepFiDkbyvt5EMwnKbeqaWrJCtJoSMg026eijLrKJrreAsYZrvM9
89DA3fFq/PKO3huX0va4H6rMMBXZJdmO4yRvFVj78wK00RuGZyWtXiRmf0U0W7yy
ETymgVzlWEZo8KgMBGvCo09uzsbBun1KFR+eIgUoFHIWUPGvcLQ6YCQwtO3+EY8n
umTohkDTa9CunVBN3Cfuz8Tz6WZSUsKtukNwxLpEdmzqi2wnoE650Pmw6a68HN/H
aryDfowhhg2L9BklGGMy9R0eU8DftZlShoLfp8a287ohAHOhYS6OprxGh7YPzwMu
gJBzMOSyamBOhO1xHYiwvbdDWQS9q7ch4INblrkiUyLr6mNjTBKVrJg+ifySAKjT
TcjZzebbPovC0yO2BiefNGbXPVXRaBsmQg6SCkRFFJxQ4EQI5WMiBHDv7ikQpeQi
rTyjM9DoOlaB5O0DBfMMOIJZ9QRiabz03Q+VkgEJO6IuITQPEJ1igBsfvFHcOFWq
bWD0piyVAd2yXQITg4gRG/PRv1JxrdxWGajyLyFJkVHv9dQfb3iP68fv5TfBZidT
VFGaoZn56vrVWC9TSsN1o2EFn46dtBtGpp4tDSwPAbC4z9KNcQlZDIteTriXJb0D
/RL0izqE2+JKIhYHjU2t+edQTU73w3WK6eQdLz/+3/2Egc5xpa0qNeAbuU2Jqm68
pUCa+9yxdNq4iqJ0LezTF5ZwrsMLy2L4N4h7dWfz8ORRcK6f8GW+QF2YdXAyBTAV
YlUmey5trRqgZ40XQiW/lyfldlih4i5fHcGqZMWLKu7anSk2QFVYZlz/ZpmDBbau
O0jvOSQSh4JObSRNJldGUCgijDfydpmiSlG8QSDVhwoIRyVBKR90GvOgQQTIR5SH
LgHxmwrZhFj6zptKw1OOCb4iJFVyagQH5TC7h5cg3E8p++UJmLmpZLwqSWr0yoZ6
YwmvMcLzXcn3NQcMMLfku5JLTesb1mD6p/p29EUZO4V+UyrCVkZ0eyobCm7aE/EM
LieKQ/eQEYLGRRdlR49JEDUpz/3HdpBzUtYBv2YPVxwOHMfvjlYtMai5Gab0J+ic
7HPkE9a31M3G/bCm2X5h4vFBTrSjCAXpEExS7qYnCkz4KPQ663XulIDfVkjrskjs
KpFGpOdLYTGeuQIKGMtMu5nozykCmRVlVm5IFlJRUlNgPK/zAnj5tiTv7+XZV3dL
sBFTU3gfcsWOPZw3ZYGeTugKkhjhBY+2c/rXK3T/D0+CaUY1wZWyEOI0KmhTfGHK
Ex3mHkWWh/A0EVpWOewcGPuRi6Vp8+7KDoqdvZ/moVsPrg0gGrFjyV/jTdPBem6G
ibwnFxgZXi5YFSS8nta4QXTqfG9RTdtSiInkxrj7zhKnk8gqVccz+aaBN+8ZQMbx
fCJSHaz797f25eAVfqTIuBesD6OYt7Cb4UM0J6z1i1IHl1QAJdwHE8gXdijdr//m
D8AADCz/rHMaiiIy64fJDetNEPEs58kuPZF24LLZrx3OUEg3Bj4dyQtKMBFoHeDe
mkOpbm7s12cDN+jReIoCT4FGN9OBjAvch9Wh15pObD46p4Myr9fkiBCQbjLU27bC
zzqE6/d0W+5D/ATQmZPdIRsmpevY+HI/teEeGzyNfnO/G/Db/GvJQoRNPQ1UanNn
RGd9OkYZgm5r7d3KzNkiizqNFfnj05pla1BEbnVzwVr962GEvthHOtVXHIBAfCAM
CwEz4y4EYkB+eJB7kzP7hjwd4KR/XzkM7ko/A2GNpffJ5Yg6eDBwu+YZbQObip/9
DA9BTGWpIE+Z2p8/SKMV3DYDM6/93d4WtYIGeVPFsisZ+aqC6gtIi0Emk7C2fSuj
4vNHPnzNfvhva7ZOX8+vV39tEMvA9mPInmiS/ITm1xQVE7hLdP5aeBdwa0ddxbbA
I5+wRttq1b33u2I89/z4Zm2JmUKijpiOFrCiDSsqtzLndiUN8VCMU3h8rymaKFq/
miIsWrWrsoC1ePX31IrkzYEopUQrHK0g3kH6vBJrfGOWDMWOsTVZsfbYBzogbKJk
GoEooDFDhrzzNqzu19c2bLP4dCDO5BoL9GJh1n4rLmAjO0dmegG0jTl/caQLvpjD
O7L0zZdzY8rZRPJEltzEdz8lptP3muRWk+wpzj4YGFNRiIq9vmMVvovzk6fcNGzb
p4k8+ofwXGy5nICS5gmbhVROdBRGwQBjI5YNNrPPKQnI6jfUYTtB/t5lTcyb/mln
f/JpI6TkQAggj2XiMU/yn+O3Y4Jo99J1bWbWgJJirt8swDHihXrDZ91ELXhB7cUK
PXMzEWnZRbl2NmG9mb4MICygEW+EuvTndBNjqFfQ4imd0rmJ+JoPjvrSxOvEsIFn
Ve9BST7Xul1Mr8IObEHfZXf3XoKsT/QrhVMFLjgZCoFiN2Yj3S+s2CZPkEMwhEng
7XD8sfbR4+CzI5hmIpJWOpuU504o+t04wMBEW2oWoHMq4LY6ZXZ48zcRghcexDXz
8mGZatO9fg8MqFfUAotCKuenASCXPQYdRElnZGYOP98HD/OOV2SyEHFu6KOaj7JU
SS0dfu0LYF/uPJZlP7dJ/+iDBmoswud0RjXTUuaRk4q5hvfswu6va2PRBxvHFdYC
uYwLGr+4EURDxdPJvItj9aFnEqUn2VpjEpIIEIHw/PA2d/FXzy9EcpSuGGslNy99
wOxGXDuCk8vfPW3Br5ztbFJu5exTMaRb97CqfD/T1cmxNKZxaSL4kthWwziEBBGQ
EWDAnHWyQb4DIyBIrPCAMoZusOOdFLgJtFvAPM8E5aHiRcKi6qDCKvtad2bUofa+
lz5qt9fdzf3ZJEMQMBe9P0nj9HeNqajgvTOwJQ72Tp6u0ahXrGDnbYt5n6GQHapT
RyzWmW/4DMv+S34UcZAL5RFcw/fH6EGsNvbU0Q/oO/1GvHBEBfAHCV/wQ6M/5vyr
9vtqNSt7fdJognTKTdBrYLP6V9GQPA6l6EQbkVQm6kN0x8IU9ELoC0RbU8uc1QjC
fTJuwo/6SycT88YgSJ0DeVRpxnQbzwtX2cv5WuvZxIkogqAPIFWLPdZWXmE6l4NT
95QzvCTkTmjpqCs0Jf5q8XpzU3fKNbndX+lEMicWknxDstfJSRfnelDKJjx8hCDq
O32jlZmoxnpBtxbQJrG/4rhCxYMrrbiANvuMk8nCJWdnwhYsX1bXZSPnOOqL6FBa
YHLX7CqQIlCgb6MYh5ep3MknHKBogKgn+3HYQFommSbWYKVLd/Y3mTAFsdChmlOI
3HTP2F7o53Xdh/5WWr1sTS3PO8KxdJSK+23rLdtOWt6+QQzFuKvj6Hf7k/tl+QmS
a6Yp9edI7/uGscSSbzFIfqBZ7O85RS3Dp+mNwjhWcEhG1Twg1bxZhSLl+ftOz4D+
aw7WoNnbuz4jOPUkEydLLH0xqt7hBzvEF6gBGWpkRm/4Iid26m8ing4VY2/ZT3Y7
GtjY1I/K96Wl522L+zTCCG17qTdb2WERkjDpxaX/kEmi38dBFG/cxs1l/Pd6lzxw
LuH2L3kA6QFelsNPymnkEqSAXbc2CBonv547J6ftm2dbAE2rJE5VxV90czwKQ0Iy
r/a0YyyCKz3Td71yxtwlQ2zcJFN+YAtFOdNI75GE9juTMa1nScVJz8ojq+z9NE5o
xjIoRjR94FpKsr1QvhI/uzlcblIzdGzrbCvWEEGwIalhH4Q9M1yngd8kBzKwDeO1
v2R7Dx+VA0hIYcDTtqsEvZ+SNWoHPtw+nbJqnCF7h4g6c/sozskiQTpOdVCuBUOT
5zws4kEu0pR403UqAkSPrC3C34ezcaS/GuVNCPDOtz/PZziPnlAsQeQLQVvX6wyG
28ZwVUsJy2ci4a4T1FayC7h99WblSzFVag6Fehm0h53BcGPfiIPKE6yu7fe9sP/K
IbPS45FJf2D0NSD1cMbvhWjjKxLdZiOVPWfWDdzTxuK5pP+Zto8m33JfbfLfKchS
Z6qQ1Td8x0M/5HEQ10cexYYXeVwWsnRoV74mN4QnvJL+k7xHSQyMcqrGdoV6xyVG
QWbbcIPRxjP+9idRBVCaSjglaFboQuDbwdLx0Zbm/GeupV9OKQrULQGL9ob8TFkR
+0Eo/HA7jDtqpaM/qaqqUdq04lCweQEBR0I/EQxi06gAKi/wyEpJZbfgyPQsLejA
`pragma protect end_protected
