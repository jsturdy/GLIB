// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jd829/zhjE31ONX13oBgOGezD7gb+hVNMPx0NTG23KkrJ+i4wGF77ggo9qbT9d8X
gObycuA4rqQRZT3xdYgOWxKrixVXSJjp/qIlLyCAWtAtEZuEFkO9GE6PPmbd9pw4
dbgATxKCq+V3sJD0pHcMWPxaTbM+QHOD6iFvUzCXiGc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58176)
RfmXmC2TpkqP058HMH7Me3TRekQ1H223+ywOcjp0NuBWZmhCT8qegtSYHEOUv6LJ
zC1eLACFGaSugYKu90YF7tme3oU3VW5IDpFmArPEi+fPQilMyvsQJCMN72LiT2Lk
6oUxZBgTmuClme6c3Wn4ubS42XYXrPieYTJ3CcfFY7BIUbvroLU3EEvRvjpzYONE
q33qfh+TeRheHBbau5Fbm9QoSTxvT8EFZ89voxynZkVLBzggww2ux9MnBNp8LR0q
wJfLtWsmJ880UlCLu5Q3s1ozR5ahkTW+AZVoDlvLucRw/oPnfBSAFsl3npjNlSqR
QY5mD9SbRM9Xle8FghmpIUkyBAjVGgGvAJx57YXi5WngUtPyuEMoF3vy1ih58SOI
9YlIimGcfh079eOkkBrdO17V4KGw/EaPYPb68g5FKXpr//Sl21ptKncSULqp3z6F
p48C7dBOQMsuhqUUHQYMOeFQNdz853kDJXt1ev7bt/ikoIOId2n+Obfl9fCdBXUb
s2ZhrszYVKb/KgCZNfQ0agxt/52oOnC2HZiKvxDZ8CJboL4lEmMNTWOUkfFMJGGE
OD2iDp+m2fQ8Nmnej30EjOyocK8OL+xOLH8M46fq5VM6r/oKyZiFMKetP6pGqPWZ
eOYAhNx/UZTeQreAq6+WyPci7TwUAyAswBuFuYDcsPOoQ0q0l8Ye5HabIZaCVrz1
oeQW/eKgaCmNlJwUzh/2zIpQeurkZadiIc3fVORpHv3XKooRp39H7avXFNAlaWET
oaTkygnL7f7xKq1eEDU0d5Gso7jxm4VBa42hy7Aj3CVRmeAeO4L4+OAXRVfp9Pdu
j8epe0BFLpsc9ZvkxQsYQ3vEItN8IIsIIpmSLyfAJJ5CpIJvs09T+pN37Nrl7+xc
yvOm5dT1KcUU65FZglpYW0QWeg+id3Sn4PLeVlKzPkG9cQS2xg+F73V2xTd4vgkg
lhiBsaokG5Lsxmb4+iV2e2B8KiqUD8Vxy+5ujhRuIs78rJcj5s6mzUC+jdziaq6u
dM+iL1DShpMXRf7JR6MW/neYLbv+pKHCMkgExq8IHGSStWjJu9KfHTv3HgJfiIgD
By+NFCiQMprn/0ivJ3Yb74s/PxZc43pw66fU0D0FEwvxAgmps963kDTIA5jRn77q
jvuDxIMMGaoLM5W++/xk8wW4+1vw+zSHnHH1+dLpPxqTgBwgkyjERQtJ0Y7YA2AQ
qyLbGjD8I4YYuj7++y2VVApzBsIFd5uUeGFs2Z+KsApxRZ+24Ac1J8cJf/X8BgJj
/aXTeD9uVDCI7Bw4ZLHsVxC2BkhvtL2Xf29+Vp08QXOixMOdTXfEq6YLqn/4FZQ7
/n2m8uGG+SMuacIqmzj2uqQyfPvARKbU+unaB8LXXDvRpLq7BWBj3uZJ+uON+6Xo
I6N+cVaaaRZYDC+s5XQqbe33ru9LYkvcuQOo030FVd7ghlFBfKpJvhm31B+uxyvB
y5qNZn3xJjZelOahZ48voAdc/0PU0/hedZyjJjdPznf5j9Mgi3HY5afxcGIqwOV5
Z+qIQ6zbFxfslxzRm3fV4Gga4Mf3vOCdzf86LWSvuc0qwqTREe3WIhV9TLL0tR/7
++Ti50EW6mwpFqJMqEzH+f6c5LGnXFvXcTnH34P3xVy2XP1+l0y3LLgV2QmR22hd
u29ZeHwTYfWwS09qRshckCOcmyB49aJ7/xt2bF9d2tz/TPOK27Zwo7y5atWZ3xgl
DuvCGpOQZ1YjAiEjljNAtGUBAKT69YrRCT36qhhomKhGTwD1gg+AaTR28fWRNGU4
z+StlpmLp8v/AqzCiJfKub2uoahGam+wio5gulDZdyMPob3x48FCTaPzcWG79MPM
jkAyHYnjKoR6RiDFNVZhlMA7qaH9MPr9vT19BiJ6xk7rAgf8ZB2HKjexUOsdcYnu
pXoSehHjL8COjBD8ryGt3MjwSQIvlPvLjgbtZ3DXWj7xLDEupyhfTCFkggvAliSn
LsMqY8Ofl9x12kL+GYYHv4SHP+5VvFiwwPbrM7BJS8nN1f7EBICQ3d6FljS1GPkt
z8eG+DCaQOELIcHNqKF+9rNDmxxW7rF/D69vUYmt2Dje37R3I2UNQw+iNcutqXiC
B69x0Wcr3oHCxilYP4JY/XtAp7Oyvfc8oBhqdYU6bKmGOGT07rabkyOSnqP2ysqP
XUGZLw4VcC/92HuJOMGU0I2LEwTcaeo3PKu36T5rH4GxzK/J7EMNf0v4b3Pdn14n
WRhqvV8wezciSv53N/neH2m06LoPq4sq50GEb5shpw8aMJfqo7wBVFrBpS/nhrBE
EWEUEcM+OgUj0KMNtlpWqvKnLsoIFI6HAPvNbI6mBZp9NEraqP3GUm1REv7BzeIm
lOH3IIOoMiLxAJJ//yRDK51sCLL7DAmINL5NqOHf0Eo+Q6vpZ+mLpsXtRD9vADKR
HkfN0Bl2B6M4hmVHKNyZfJr6MM9arA/clj0xBOh7LMZ19kvCwTVdm+1bfhKAIFqC
lVyt7A0uf+lftTetPIsMrZGtwNhmffxIHH6V+l5cGY4WHvufZGNdbBxaHRhEWwhn
selFSF51dDXKdDvczGWKtI+6yPhVxkXQBEilKJEmufkzwdvr3SdKEBLk0ulPEnPQ
Zj8qQhk4Nw3zmX0j7KS5xRPNwerdpbM1lSpOWkz3APgg9qhSgpHq0rjvyWj+fikH
o9zdXqJ2+3LkDwEigeswypIq63MvGgvi/aw+KoUi2qzEv95EohG8WQeRzCZvvna8
iT14jJO3Pzf24wNGu9wb/Uzk1n3RTrA0vlFgoIocfGPucj9FVyJsmdrVZI43Fh4g
7pSzhVx4L8NSoBrP74h12zRxi8NpRYGTVNM9g33aXfgwYUH9idADfpxEz7uiXnsf
5T8BskJjYVhD5eOwHYAmH/mgnOCq2AJ34up96wEX9p7JZaqZTD2JodlKUNrmWRIN
iiNUW6J4aroVDAFI5uYnNjApbnGcNoeiVS3Xizy9syeYHP5RglZ3SbKhVhpB19LQ
wPEdoQ1/anvZx3zzPr6OrbG6AFJtEQkNiTYLKNyUSZ4WQ2/59aiEk4bd+DVFhJ8l
jiiO9ElMS8Zj0Zizq7IfdeLIgOFEuH2/FoxwnpxtRrEiaw2PBKhiRy7K2vjPkMqI
blQB5Vj6CuqDOUlYAT20BlZ/NyO7QQW1p6F4KXEJe8afLlHnhMkoXufbt9IGBxbR
rywOPM2YFP0a9iHDQzSVgyiJAVptDN0QKC/UyQ9YcZgAdWNGZJSdPuL81L7SLVoT
1QvieZyMDtcoriSEJDmmqYWHflkho3l7qTaxFG53/DhEeCN0QBkS6adX6rsz1V7K
2V5OP8K0ZdeziHIpPlJjrlADczPgMAYvyEpBfrGP/9y+sSFKQs3onCiWeaHDYitV
HUMpWO0nFg6iPocC+3WcEVBGxkLdnw0+vzGwxaYXL5MYKL8+FKGqpN7SC4J0JCjc
KyB4JF026Exa66arMD8DsWGmkavmF1NCZhqsXxt7hP7y5aby3y8gx+zpbTG+lA8e
rk0mao10iumzCVK/kKJUwIby9GF+Mw3VPaPsaDPhrYFcZLD3BZ/0H1H/+nkhHfEk
GUJkKMipI1WFK13nFcor7mKoIQghp/zPf38sMtYPLbgF5WAvzYZdOjP88qTr7SEy
FLDW3vn91xrLL10MJma9xGijqTxR1NEGPJqfJgt9YFCHmhXwmNoU3ik799vw64Ii
bHUWm9b1w0e4sBxY7F7nSt4qgV0dHi5jsHbuxqAyWoGjHYLKIOQBZMkRgoqX3SO8
lN7oDcdYCYyveAt53prnJG7FmGVgE2qbCdcloeMqZE5zWSqbSn7lZQ9YcYwPE9Gz
uA2LZZE071pQ8hDnHI0q86trk+dzzYwZ14U87pDCCnR1grRmwmciDVjAc7rsxMRP
fGN/UYisVQOwXbf5HMudSAUTuz+ZEnIMoFfzYe8/rAp2pZ5OLTYIxdyJU60z2/8G
QvU1uGtwY4S8KAwvyf7bqvq0PzC6HXh6yTLtGxW1mfnLdidkZVK9jFak1jwOBAb+
nEPaEGSsoc5OxlfKqzv4+q5zUQbuydl/JEpzd7Eazq4cBD8vE0pL7/O3oLuURgs/
eAi4G5bLmtT4SD1c3WTvB8eGm5iyjZqnWShSMHRotDLcZHAbMdHzbDHAkJxKea1p
zkKhBOwdPfALlytilhUG8hF4eogjaiO54LSFucISoQKzxK56iPPtUsICXaO2XgQJ
hqP0ftGYVFzRNFixd9jeaoaoN9v+gOZbWxLBWvs+h8au2Y91kC0MMiMuMT441EJ8
PIHZWccm88zTfpPiTdvb1YetdlgfOyNK6FOAZE31wK0f+baT7uMYHYG904U3bOtM
F0kWVB67LwU63Ia2h4QGM0iY/7zXXzX7r9jG+qst50IRZDtVRxFFZUNnkYSibkQy
wf9NVXfmVz01IbJPFZMFhBfL4ani41x/nPTfeq9NjmOZA0rhSizxl9lLKFBZhvuK
vN5i7LTWB266caoqjLpn/fooybLxTh/CBmw2tloYY/uxFw0LABZRecYeUN66YSLw
1QIb5xECtA/Qhe+F8zrVoecwYb5w8MsfVDMI+GcohF8jPuIM7ZDqhWdFPjYsqK9Y
WBVSugFSpsqRa7v85D3U8kGlWWW29SSkvFUKrWgj3E2/HG11SuvAD9GO6WNs0bIS
xq2Q/0qyitlZ7fRGoLMeusoKT4vU8ShhMvdBffmRyy2BnWQpH5Ud+058MtpM/Vke
oW8Tq1VIXok/D5ZN9LBsgj/J7CGOU+uHmyaruV8lDcDtDyzmPUQAoN7Ffdn/18Fx
ZGlXn47OMF7hzTrR4jxzuN3iZDFJxZknbxbRHTEXlHeZe1bg8pTEEGJAoVA8qfH+
s2/DzdgkRXd555bo1Nz9E/pWczGVbbN03ypEU5CE62zpgxg9RxdKMbQJRAsTV7Uw
BL78jKyq+1Zrmd1pO1nciFXjRe8X6ADr+jGhIGrhTJC9XgcFgRgXLqs9MYG/X12y
oReg5KTq1pAzNWDYgpGq5wmjjJD0m31hZH4RldYCM28pCmuCTGfqLcfDsXWmJPW0
7G5VcqmcM90fJlJRWKMg8WyfhH2keFowfb0kdRvIZcxqGlrQUbQFcfHVJfpSKV3J
63UO9HL7+GGN5IvVp7zEMKmTo4Ebw3Cl8khBSeLuSSqmk/hn+K61iCw8JyJp8iiL
Ms8P0CY5qZX748iSmTCl+hFyLWcEPyvyx+oRmhstfW3BfnUfc5Oy4iUD37+hWsu2
L7XHvD/SSH3wHlFpKWjVNa92hT6mcY296KJJOt6DNImpQzqML6HEZUkgB0aptB3y
YjpdeAZctBM0XJdiDDP8cUYtequSpZ/uXc4Q2uAuq2x6BDNC+HCEMWrQpQqv8a5a
/ft8m20NIdYHZn9UUMfXioz6y+e5kl28nktYBMWqjH/OXabwJS6+Ty93pOuUZa49
RyfUnN8dbczlZo7bQi55G0ymSzTWpLdmaF4BLWpkCfc4FxX6yxVu2gs5ot6ty7EF
A0pcuF/fUeBghbolPPQp1zYnbsi4/i0srStEOK0rhRhAbNsvCTmsZj8ojSR4HSR+
GeuND8YjG3SAbWJpiF1DxePtZ98MU1wQtIPw4rR+lGfAL7/3nZjhiAp++KoNlMNm
eeg4qcgdQkkYkejOnfEjJa7ist3aQXvYV088D4xNk084b+6qkW1TTvc0+Z51Y5wQ
Vil9333TsXOdbDBmY5Pr2c3UbIyZ7uD8WcwyrD/x/xy24fYPR4BpmrD1LLYCDqrl
S1fRTfIyKQwId+6WdBgmWSOX3DyX+MsYWnIitfU+AaJatoWxl08PWP8u3f3G4AxM
dWB40LsblLN2VZ83nMY/EnbdTGg3R4YBKdulHhjtnJXgbQrINOOAUJnCptYCGGqU
5oy2gwY/wep/s1B+pMON6C+dbJW0dJknMj/y+JNfpr0/Mc/z05YgE5ZQQPhE0Idh
rbbhQ/2aozX0pfaLgCcYn4C6WQTZ/xEFG2+jlFE/vwkLQ7IdYIn1CcNtn59EcyIG
thHxTRKPrwHYSKdsaqM16ZacRQWzc8cZ39zoti55JQpMy8xIK9IQnSOvX4UfslRT
k1c2Js3xWqv4Z62JDufxWulc5EpRP//56MD/N1k2i8L4DFO/xzGP60HKNDW2IcZu
fGOmtlEvDTnjYKa/M9U1Ete3mdY5yAALU+496JcAIaAWN2FH5sMpGpow7ZAGpz+a
7WZmkOmBO8l8YMgNcY3uSd0wDP6KHyuLzS1RphfdZb7OtzvkBsVFOILw1qLsU0vr
b9jGPcU44QplupLtFkzt+Dw/TXzdaNfNu/VRKn2RVqCSYVzXojq+ttZrvSJrEiSE
vk/D9upll/OJtyBT+5okinzocTLFSAqp5mMj6tjAYkGYBvKRwRmkXbSfd4ca5aVr
JYLRCg4zs135ngngCn0WozD0nMBWPg7gX05rmBQdJqEWSfVAUonPJ8pRCLxOkiIF
8Iz4U5TQ31PQ3DjoBWJV4I+3AILvNzUf0ieh57j0GFS4TivHlPFzL8zyqXBTGFf4
uuXy/ptgqtrboSg8nZxZmv829ogpZc66t40FH1VriR71ylpBFe8fVyNZb0PepPuk
pQoKYkhzl0MUwxzQabfNMuW4vxgThab7t7IXNyuGizp85kK0jlcuELl9D4bL3v7k
5WIeDK2LoN8tA0yoS5E7FY6XHj9c0GDiUSpnvYbLIHRbMvhfBHK9LPPD3RzJ2cYz
0WlWtSHaFiObg86s1k8rE3habBRbrsuUYJkUY3vP7Gc0Cep/bLotjCmdhgnXmcA+
T9q4q3jkH8s6+xvzMGNnkS31SlG3q3eRFoQB082Fg3l6WEj7nOWo5o23tiwJgJo3
2CmSnEvrhlQ+q/HF5VeN+764FWbCoZdWr7jxAUl/R6kmotO9Nbwtra9fRixOjLwR
jDHKOsHMd2nv7BL/6ttXorIeR9Ohe5ekekxIB8XHMd6ATrlTmorkycY73Dk4kLVL
+25J8p9RDjLhrmyoqRUGMOR6uTCuzVseXgTtpqn9cL5tEPs3n1A4pVy8mbdTJB7u
42l++zGoPHUg6PNrlR/r3Syvec10ln5X/Q2Fcbnhk0FsTQ+Hb7oa0CA0gXE4gHF+
8Jqjtah7QTW3ayly3rJXsQLdvh+qzTJ7FGRK0X/dcs9Leh9VQXKPnCxwYIj7/uMq
3YEcAGQif1RLYKQrCFzWnJI+4Fw+tVsiDHa/JkNYRJELpEr+wGoOeIoB1fpSgE+m
YXpLTy83/ehnAmsRXtJYCTy46e3cjgyG9YZKBUzkcyFWPq1Izc9/TczkSEQ1245K
sIc1D/A4KZkTDRXx9pjCXgJgNtJzmC0nUKPMVcET+O46YdoRZAyadkX41zD+yVf1
AjzCon6P4YNyw7IcAT1PGEk2OKukeEnmEsop/ojtfUYi6pCGkBiGI8RpPtdnXn8w
6kUVVRqo/swMK7eWpMIp7MX9ReBVvMovIKEl6cw4LOpfL8JPHrGDN99W6ca/ff9w
JNXa9hSmYh6ao6nEYBoZkei1au14jKANwJtAzP+rX9yHvFd80rSMKLLryFde44yH
PdpU34r+nMnZklc+X8euJVar85PHQBHZbMlfw7Iku13I1+HZR1+EKeUDkunfUhv5
Vkfx7C5wKczHgdmvTyK6jidQDXmGvx9HvOrGapXkSgOFr54c+5BKJKAdTRjTqMjX
U5ly0xhjHRpaXVpnj2k8XbHvhi5LO8VTmE65j5DYTsUKbzOaIVYxbBS/5jXU3VlW
ZGQJP3XIrj0GEfD95eJ58zVYaOZkKpQ4WBaOO6JTyVlK7Rd5lCXrGVG6d6vpx5q7
OFoMA5/KG8y4NO4yQj21xrRoXOTTNxPOYUDTBWH5XPv9NpAbeoHQXIHbtSqnvj/a
wCVUgnQwd/Z1JsTpRhQXNhj6NtFlCZnUQ0DVKj7v/JHzMg84YMXLcm9DO6arOkgo
SkJu3pTVI14ebbDFP+24wNzuLWwfUN/Hdwsw3+e9ddwofbbdrMvPPn9XxJ+6TKUc
zL2DTZG52apiXIdr4h4qen3rRToLD+bpOgFHX1Z2T8HgEuckTgiksJXjLXh63B80
WCGiHY+Jv6xUVYABC+D3UaTHLzVT+C1wkbWRmbi26xxoN/6q8N+GIi1LK/+xsn5s
b+y1vPmneknVgh8qpqd5qj99eTlCQTFsku/KXwhniwoOReBQIaGrIZA2LuS+1mlE
hUEZheHBvb8UaJr2mP8a9vlc3LkvwxeUhLDcldis0vnfHRuLf/l+U3b5Bi/vEh8G
6MSq6D/o/8MuilAQx41VYRi2KyZtjzRUC8urfh4CIR3eWMcKc1FdxaHGmCx+QCOn
CeHxw5ybgNanm1ZMZilUviA3Qy/6xBdgCMfDv54afkYYoaHyL18gcN4J9NvymYB1
GKuwBcsq7pp3ztn/etIH3g0bmc/MVNjKcV9gIRqNAYOszDOtbRoEn050IxzWMrE9
iz8FlYx8NxcN34+A6MSyJeLgN+RtvtWtBhldQbGc8MiPYmgOTGyqQFQfyhRDg/QM
SP07h9lzwu1dqg3BmIwuhwTPmPmPFHI30E0+YvSKWnsCjP8P3ObxAmxijnyzKUfF
p6hL3Gb5lGzElwi277LqqitSFoxhDK9hvIpgMJpa+W4lV5S9Yro9P4NdtfCdgj8L
DzA/+lHhDY8NSsIX2b0hh6IJQgoW1/tyffHwqjZdc7fzTcXO2tKXNgo6MUVYbbQq
KIH+5o0Ck5yoP7xE+wZ96qFz5hRaYKdMWBdTcLIY00OkyK8w/WnWT8o1r4Vch6gu
SMfWTnO+D2jWQ/B5FSgi9YOgciLlahcx73AdauXoqU9ehtT2vShsjVMetLE2pUsw
edc7gOlU9HgWlTwOSuCZNDe9itaFGxNP5Cd5tlhIO/2cmMSPKlMeqih9bJrTSqPa
eV9jkxD/gBTWIUI03EtiHD30YtyBPqDSJcQlWBh/kyTVrST5k7Iy1uEaO8Hj7Mnf
Jfh86TjdQHGX2ZuRWIeB4lKBagagFovtK4G36L0b/mP+hZBuxYjtiOjoFKvuKmd4
UYoao6E8pvQExpehk7NkKCM193fjKJWrzocyLD2fmjraAGDsmnzJU6GQkiIFVvVn
ZPOX/OpfQIWl8hPxnEy623cUq6+FJ1BjBNwKj+mtTrrJAGRvhDo1fIJIM+eQfDUD
L7QhRYGoJNVg+AV3Bh2AlDZGb6zpDTeZ2rGmDxUWEhFVxq+w3X9uP8XiJXgW5jQA
JBfD1hrEkuk3hLDGAR5jf3vHs4XOGwmTXO6a2M8MPoykCKqKnFYq7qHlZ3RkX1rI
6HVgHKQ0vlwMArU3aOkshHxJorWjuZC4JB89GF13j6eEe2zVe8wY08fITmhQfpHm
DUe7nbJurzq3O8KzyuL5LdlqVogH6pUlPJnf+Dw9h3yv4P/V/lay2pvrS87ryyNd
zmbiBVJxcd/OJ8wKFx6xd7RSl63OPyKOyq9j+taXbpLi2kocvhkxQ9tcpOFyiRDV
dDDRS5Vg0Bhh1M9cjY2Gv7s+aR1FZoDOyG2jqOg7GhXOfAtMh1nOc13zXDCQWmUo
piv+AkIYKBDTav0gOLR8n8WfKGq0/tWHi8TbTDYmCo7hXe8xj5MpqIhDQCqXBC0W
dJrGDXM8oNAPzEj5YowZxGN9m6Y7TsZS6bkHAl9OLwoSMtNPTJ7cb2munibMXZe9
Vi+qqYbJplCWBalV7hn9krsa6p4wRJLg0MewT+BoaRCK8lc5JNMeGx73xClmw04n
azv7+vzJrwtbi877f8u36yD1ZV6Bqnk+StAz68N7udwkifAA13uR73ex7sPqRDUe
f2kXn3drjlX15sXbiqwIKfm9oSBcTQ/ufrvh0Bra+dl1vUYd0045ijnHUBz0/AD1
QyhfAYI1/qWBJ8mRnk4I6Mbf3W5pUmiShlxvSe1jomhiN0XgCyH4lcXCYApLFxJF
fzqUD7WJpDsU06RA+nvhf08bkVYfK60gWN/IUn9C4gh29j0KGECm16PPiumjF4/E
GgB24gZW2Gu5hTIp+dVco6Ci15ClaksmFFSpA7QYIJdcZsS3OS7015TBGX4J8ujl
DnvX84DzUYek6Td2jgozGJR6EnqIxcs1yNC0iEzSk3trXtcWG/nArJaovPiHm7MR
PkgrqqXSEDOYjw66FhFrIbPLY8+u44iVUHd0PhUW1FjpypnTb87Oj5s7ucPE8lxF
kW3RXKvx1oJyxhLNPt1r3h1itPQiEZX0SZ2vf/R35ziBNT8dYblhwnNhCi73X8Mu
YXWZ2scF3fg4naNkvI6f+TaJuROl1dmEks8xHndK1Ym4jexUoFkru3Z69hXC11rp
mMMLn1SPOjBAVGAkHbqjg10GPZs3D7Z3AZAOCj1DjkSkEcA98zWJUIvuQ75PgLK8
JM0Qrnr0FuGVzDnsJLTqHmKwcNLx7PTtXQc85+LvWAOSdB76v+RUXZiijsZIseq7
BKvZg07/+Z4iFEPDOh9r7uJupgwcXmtjpCVtgtdKbq3RfFUCbDJI/HTzNqGpEzCY
Zi7/VDTWXVezVxAIDdrcBKvWUIRZVqRgZi+kZiQIq3MFdU8DDlnZXuAiWHReDDHl
CCN363/EhKcm2UPN5ngHx2JEGN7ld5SHLJD6RKqjsIK1SL6DoVYhWTfPRnoZWNlz
b/ACfesboPJcBLMZiWjghwBtlfT/Jhq+O7+lI5QYrZdz4rMsZ5jm8CAJ85uh2CfP
NJ6YENON0D0lr2ZWoiFvEGBbbT6CMC2LZSg6stheiTq2HfqxFnLM6aBeXRrjUTt/
lwIvnBt56HeBfJA0kqOdZDWtgO3k+JodRo9L8SYBL8C6YnpgXnmDJqRUqcAj0fBn
VhZrBmYkgBtWvDULgHYrYzM3k5rJIEU9L5AnbrAxCoqdngcstzcf8FnRd3jYNvZW
Iwd5mtAdmCwDrSbi37JAotTxe4aoiZRpcU7Ciet7Jw0FkzPzFAXo3NW6mIbs486S
GQZmihP/ZkDOggAnVlgttuJL9SNgn8CyjrG4uk5THLnyL8sjQA0cJSoHvfPiRk61
oz9Mf+fAbheytENy+syYjqFbiF3fNHuyaKk8Z68YyyXdaYJF2b/dil6qpEAK8UjL
7LHJxuTG75OZw7PU15wA+mAmv8VQmv+e4XXZasEPF/yUpG7O3dXc2VlD6Ejx9vd0
ugmOhnviTN1VLm+bNS4CoDY7WWSmJT2JGzyIurTDAyzhKAOYGHVJY6256ly82M0T
oXEFfXjmjhI017yE1SPuOn9ajvNUOJ3ztoTPjeRVKF6ioq6STE8rjGpYDsrwtPcq
cWnKkGqBEseTUuQlALTMnhk2dIOKxLek1rzz4IRKi6muEIRGezi2l/n+S1K09dD4
07UB6WgeuOHfAaCOJtrJuEC58opTJVh1FLY5IcBeDhyO1iu/Zxd/JjK21GUZ8cld
qk6YoO+QXStI6cS7ufwNQ7PzGXQGzSyQvU4ZyjRZW/vZf09Jo1mV/DViaOu7XjaT
LC/dwsqClrtpJbQF8v8oR/5b3URYKynnuYrz8j5D1Xb/g2OD5P/MHqPOZpaC57Yb
CjV9Pt7pG9QLtFe73qWtHcJWgIfqeDZLDrX7ev458Mm0VQ0Igu9WerctjiYMlK3h
MJRzoE5FgJxB45E2PAeGAC9hVI11zijfu3LoS8zH4FINCSfJTqhMfpwzr0Mf8fmn
4ouf00XRURSptgooRsApJ5toj5oiKc7JHLv//IxPWnULDL9JZGkrMqMMQz9ciOKr
IX5Rd/Kc9W4Q/Lk7AjeoP0tHvLJkcYNlCBp+TM/1Kt/VDgaqeQ4jaDTtZaOwObac
oDb0RTWecOoDkcdUcwH7uSZGcCy6jZFyXBs0duyoqBgHgM1Zt2S33NHpeH2xFoj0
jc3MjL8t1VWLjJh9C00dswZBRlPaznUAnwSt+BeQlTioAKW3ozjbO8D02TKhb2Rp
jO6J3HmoGxGtu1oyvwDFH7HWcv9C0pvbxfqk8Qew1+0VlCvcM/6aXncMIs7uTFtm
1vvHeRFkf8L5+I1g1TXv2sAxY3vicRU2SWCuXpClXU2YQM0fHqN1zkWrw1LsaECA
vweD5f8IK8W+ohTST8xYYXtAbSYzBFs1OPdbQvRYnO4+X0/LrkaB1RAo7nsYYwYy
tCGYzQoWWMP79dAw1O0nilUUFMl6yx1v9FrE4J+E1HKVr3rzouQjqelxWq9zXeRq
QpMjOiXi8AUgSFEQ1MZ4C0GqxNeJ4PwasNh60IfcibQNOpzoUeVEYEwp7eGOUA98
KDl2e1nbNrPIJfU3BJ5/yjHEaT0Fy1dC97CqJ4x2Xo6BChYyjlGt+/62YILmPTgL
boPG4f5oErSEbqR5Q5+HZ4dkYP2q979PfDeiP3JYiLqQDQyMxnqaxxGO5WVEyzyK
oXFrX+tGn19NMQL9c7gS449PU0m+yRybSwe4Sh0qhYN4H3JTDj4grIX/uMmaP73G
LoyUilfoRYrGXRaOCLNjchuHOoVwpNluiFhemxD08rFaReRwojDZL/tL7SgHZoP7
gSTzTtdea36L7X/PjUdqLRfSl8Cel2Pds/qKjGgvW6jFf+8WAVXraWxQ+cDcZrLx
tPShkg7dj7cnN9+RCBhPL9u0hIKE39a/S+U+NFKjIfJgiQ+NcYe0wSB5bBgZAbrv
g3h7Ob4j6IjWxDn8ug1aX3T0WtUO8OhrwlS1oRz+PKF+sDpDGnEcEenjVejDTRaK
62K70LNVBSqKd7Jq3EJxeRJmhtDbzb00DxXyp3UB1diKB4rYiQbe23IhjZ2gv7UR
OEhPxbY5inHBae9biEK6BPe8T1gq8/lAHi7hwpRFzOE1kWHz4jxEnatRmBPyR9rK
7S7RMsUcy+wAuAoreqFw1msSDlcE/8Q40hl9JXXK9bAVPPSmGjTETYa3yw/4LabW
MrpzfUweCd8jsXsYdDgSj6BL8ZcVsCNQ5fmG09mrM4k/9n8BJzILePHuoQGMFI3a
Hx5IRReeUvvyRJgYvLT5sisZ9d2YoqGcOfkdM3tpFOFXeid3FeJGWvX/K2QcAxdr
IG0tKbehaLByRX80S4oQoUAcqs8gMzgZtT8SWTEpyWO/35v8+6kdghX5KlFKQL0Z
wkZyGAPey/2TFyyJWGCtzzRv0XCG9upD8AiFUswAgluBdLnWNJP89UdjFB21k0bw
P38VpCew/KDjcZQLryEobBEzi0RR57se0gooZ7ubaEvTuXDjBELsk4pofwUIA7Qw
krxf8wHTOC9a2giezjfPBAPw1bQMPT3TzuWgTNg2UowAwJ4/V8+2WqjKURTYJpVX
LAQX22sq8czU/87EqxCzwCg/OvvHAyD+v2KIq0suZUDQIMFzjdzcvwM5wIIFsi/w
4ytWWZCagOSKdQKG7fgLT1PSu2HKQ4ZXvvmzjoOStgyW/FdwHx6RL4FXGm4uOzsW
YfU/nyK0xqny1WvFtiN/Y7xyh1vuqaHqcJWhKY5sXHnMH7EKyY0JVvjR2A9xRo/O
V3I8JvFVDcwbW/lHodEDk5Vuf9XbbINrnSU3lUPQ/U46llA1WMPKuTsk1TFQqRiP
kDQC8SgaDgH3WHcAAs5PnUIRGJlqnOtQz8rRfAYxFp6wXUYNo8IHx/rOLH6qr39K
Lt3e35WCiQJuznft4Y/z2DKdWDt6NgcvNNW+6Q893JCFB+D4XZeNblEJY48Bn/zB
Zi1q+rSk0UxIvuuRIKf8XNI21Ft9i1WH5EwvLeyHVbIBStjcUWUUFTQz02tqCBKC
ptgTT/Ur6pApDQmx/wg/o2kZV4yzKU4P0m8imeQgyHFTJXFhjji1mANfIby+9mZh
scmRctCNbig86W/nTJKg+NbIHartVtYDqFc0pY0GmEkK3h+dZ/mrh+P7NQ2pw/Al
7f9edQBBJmZ7hSXbpqaFA/Duyyqnm4tqAUBCXDaaRkG3gGRudGpJQcWkZuOuv1nQ
ov0DEov3G+CcDesMF1KFxJHnFFP2Vm7kWcyYexftjTSi3s2WdNBMah+iR3+V3ADC
5UlauHTZwh/BKbMjBc4wohU6/3bNCKoplSOSvCEJbzr6KfJO6dPg3bWID8OIwetT
mn5WpBOr2+lDB/U/HINOUEEuvAgSP2Jv2Tj01MUpGhK7tnqIGNhXLP24op0PnEWH
9ulY+yavuA9LX4aO8B8XUqNiYKBfyfYgU1rPcgkvXv8g7mq/R+9wLJV9y9jM4tLK
UyBma5EHBGi4ODuRWQlMqlb3GDRhtbd7MJCFYUFEz6nyHsIJAebgkV7JbXx2f7Xo
A/7tXHobFXGS+9RMtt/bl0mW/hjzoX5lbjFJeIpZxUIfAy8mifKaYMu3ilWdQqVm
BmVTN6yCapCDqbEIqfU0aWdiqJDolyPLsNWjTji62FF3Ms+DtHLkbgTOTwvzwQTG
ilu0NmRKTEPpqcbhN2ketQdddyI/ZVhOLyVez5hP9G/wubuVUi2lvEycgXlT4vnd
v0VvQnQ94eFjB9AA4LBps0qM3gYSvL05eBJA5IFK44Nm9TBjYif/o1sPZV1R65X2
BHSihQnXoT7Asosa750m5j3u4UA9yQKPwxyeaEDeSFiLpswzCEqJDRQif4eQgiez
KoDzKPYdY9u/faUlmraUKIxUESlgyuH/iFHL11TimvmFhFKb5qKUHeRj7y5PHsqm
iNVFtXZCrzGjUwI2nUuItiU2V2ohP9z4DUnmhqDAGjvnBn6ZHr+CUWJbZ52SY0+e
dUEboC+i5P5XQ3tr7gW5gqVwdmlaP4iFmG+yXKfNuSRfsC2eFpe2uQ6wU7hIj8Z8
QRCxn5efrFQd1r8OLE+p31wHhXhZYtBWxoCas1PDnmMcshIKK2pWCjmBOkaBiVtn
S6MRhW8QmzEk8UKKRxsf80eAoWCe1hjDGB10wxT9A3v0FvUrJycqpmfzR1XhQTqP
n5Jxgomhpxh/Epib8ljB6wlcIQmPq5RXaZc0B41AV7cjsE2SLd0sHkvxuQIY3Woc
EvEifxyZNsYscYHo/v4FjuEE6vgKq8j6ENF3nrpZHR8ezfJT8c+IOUFBjZX1fIB2
M5mtqtWTIib8f7AbExz7CK9OD4t4TdryotA+/+2Wc7GJT1laByd9XzYjIGtSYvuh
ASxzRoYhW1Ly9PF4P4VJW+QwVkhLVQH17HkzZ9+yWjXd46zCngCV+bdxe8SpWtZ0
JZYto1TnPHw/sqE58tnPVMgSbMIClSO4yrGx84gmLNcRerJGQuIdoZEQMHYARp/+
H4WmZzkSrPLVK6PUIZA7X+qNVGxRB7zP97kXW6uh/NYg6/Am0zX6rPDHPWw6wQuD
3sStrd4W4BBlrcsPK2Kh0w+0jQKJIAgxNnbkZ5X+d8xg8LKEQC59Wvr1a+dMZGRK
ZUr6ijRTspHMOcwmZMcKaR4wjB7IPzr96fmAr87gRI7LjTufKfk8NquAILGGywjt
2EUdsQ93KGZ+Es1qprnExGxCAko01u4LcpEsin7WUE40vPhpbsAe94mdHA0ln03j
kuXLHWlOw5TxeDRCCgVwNI0krNRTOiyRr+AmvJbym5upxCmXPsvn6h9wQx7God5C
fwfk0SskbifYcM0CWdlbvtgDms7NtYuvxDH2zjUd6XiL2+XVY9/rLhTi/eeP/+yz
c3xSqisiUgRY6NBkudRkyT/tmwU4ZGExuOUs70bNbrdfSjQLuYkZWCFrVUKM85wr
vXlTdJ4BN63yJUePevWawSwg98bbSNeLpussEtUsjXR8JdGKNbSyMFQMLSurv5pf
ZiyZzPFjbiWNcI6ko0m8TFkDfK+rFJM/79VYJW8KF8kni8nGc+RDx96eGmJU058M
ER8QMLOEGcHbYkAik1fKOYJQJuy36ApTDw0OrizU1uxU9sg4rqwP43Gy1CI3SbEn
q0fU527iDlig3iJl2B4hhKnsS4VAlU12MMRgX30HBU5nXzrKdmFp+FQlcY5AVbPh
/lJ1L7RI38mlx+eRyrJ8DjWBHwUSnYI3VW+gri0SKU8PsI+7BdRGddszW+5GQ+XU
d5A4O46J770szJLDR+8KZ/gCTtg/5emHKnfvISfgPYeFt4aB/w/N2+3Ti0WPrdQv
1t8rNmjdRVFAzE5tdHeHzpXO7sDW0aLbBCwViJ8LRKwk4o5Rs7zTwq4t+KPaoLcZ
XnLIRn7+FKAg+vnLJXCkQ+FhcPaJs1YSFba6EfoDyL0pklaKkTwQOLJ4CxP8T64S
JouCpD6am6w967lfYaBfVhge2ARv0enXn14lXIaQAf4gu06L9XCJJoTdYB7YmXOS
Bmx40ambvyfx6z4yX1edfcA6rCWZ91REySR0xEzCui7Mis+H7b2PSTkIwclyszsA
DeCDx6kgldclHZ44l8muxrS4sIHaQhdlfq14DXo1zim/+uEsqRh6+cAVTT74mzNd
CKDZ8ntevDrLx4bIRscZnziQ1asqGLu4FLzSe0fGIlQQaYfPT2oyDBjIDGPP6bRp
5dGUj3twmHPoDjZFy877M8051O2eXIQugwtihWOI3LXWOwR80Dc4+q/qHklpkJun
fR9FGoLThXVlUwkoBa3iisoa9J+SWHtcZyZomyJcQfX+0lSR3pH/Ux3UmGGzGH0O
boWDR+V1KNP6J+fMKX5ZHpk+BFfljY9PPukfyisQqpvPynUI9Dn4REhfn2Tr2n35
Vgjhri9rCDDnMkNGsSKb/qnYZLVXaJa9J/N+O1jjZM9vVDYssOiGXXlzz+YvdnS7
KU58v9scFa0QlrhcD622Vwe1aZH9SpvnlM7vVw481XsfpWOMaXuXnVIJtoeJ9MrM
i+QFQInCmgZBLPS14DdAo+qktUkbNjr8HbJkqHpQeCHPR1lPtayT8QNKjedNXVln
77nXMk5VlDB4pgNlKhkseMq4JokthG9/PHo8WVxE7uVKNDR7xYjmMfSzPr7T1yrQ
xkZImtadpHWnzqY72kzRjs7FeCRPC+Rb0SzCElxfb1J/zhLLD3XBpba55+wXY8Zu
g/FTcNaVwQLJXSP63RmlPBJqdo/sGskB1Re9JVxGQyQIyfrc/RyNKg9dcqquce1L
g2Q2WB8vsqMvc+3DMs2rNxMWyBPEsFiGS37iOBJGCZNVI3Z37CJlUWR5z4hOvt78
xI1GzpV5zQA8gTWfWuqVl4Eb1L1F+oyRtJCw+DJpvXY1dGzJd4nKPnEa0x2FXB4F
BizoMaVY+tP9OrGCMFXqOHZvC+OOhIyqxaWGsZ9B8dr4VNfzcXAa0OEHXV7xD+kD
E7LD4yiW6Fm2lJi03jBPUkkwvx+Ry5XQkFM4JzkpWaooLLpIVf+ZontAP11QGf6X
KUa7cZ8krfs4ERhS9wPetZ14NmstCTEMDGF75j/b3s2tNI/hwgrkWxIBq8DQnvkG
C/aX8mCgOu7N4TBJAOXeDLP7vYcDVgYSbmZ9R2zpUmrm3PTeNlcx2GxodK5PVore
h23JyDEJNGd5PracOwPwIXhfc3VeUTbXXOiic1sT4smJaYhxdpZLbPnXz3Dnt8ge
MWSTJFplUct/bwTM6V5cLuLlxdKHPWm7UXXerj8kqVe7egDWLF4tkUzaHA6uFtDl
DYKIge/wvmn3DE6q6Nr7lu7gWX4TH/3psUqhcaU9K+pHZxAOFk1LwBNJbxu7lTj3
gVTEa6ut+auBtiKPhBSvMBGDr+EeW1Bqiu/d1kMVO+sv7OyQs9GINB7R1noOd9bm
5Q0pmwslNfHPT3UpCVKjI6GjKBuJKv5qUbmSy43RfU5pK/1xuGgRbw2jCXR7fk8Z
zsGplvmktQTUudXdrA8/FELNFRbBwxQjwwyqj53Pr9brGyEY+x6WkSK0U6GHMJnB
edMUttJHnzsmo7rEk8ESd7ws9Y4w8tW6YPp8D27YAA2MiUCkPdridqsqdboksWa/
cyuSNbv47KnNyWpBSFlsM9jNk0tnzx2Xn7u+KcSSm+gOteVmNMJwzVNSKMFApgEC
ygHa5DaIGENICZP/wRVx/UbHd2BCEa8bdphwE+yCMLayQZrJDSY4PAneVM0uWj0S
SkAPpIdL0//N8/1LuKqTTnAfUBD8D7Q2zdv7HJJQcpNoy2mPmisYq9FBmUxeanZw
m98p/IZia4wV8FWDB8ekdRoq6vlkoyx3cGug0TGKodC8eVxLQLjVMsjoKI9m+Kzo
fPINFaWS1A37+qmJSVVeqAzo4QtBRSkDRiIleHpTiYySpBUT5ma1GWx707LYrKrJ
DoKyeI880/l7oDoAsTPOpLygeVx4CDp2Ahr6Ms5hfNIWObWHUDKGo0UBC+n7qhiZ
NqnG/zrECh9guA99ZNJge0AqFO5Vg+08mMlzg6Iul4t7Bk4CnGzNN16KHi56+NOr
5wlA9fEXc5lWJO31Wo5WD+cRBkugyNqp9kLHqXDpdkPk7tOhxiIj15EdIxDVu8K2
TFMJSmvoCYKBR2qAie+Lo8q6WT5NCtlMKEeM9NbtylRS6IKExvex+Tbu8cWev14S
GPvVldSfwKljWsU3b3TRrafhlHiPvqF+Z+8kBuYiS8j62g3cgdo/mNRPYMm/4Vxw
8S8SwaxQfSlDJ6itB/hYvNSgCGqB0M8s3mxDEvse7xieEOMAbkaNjX4Fij6tEL96
r9fVfm+M0wiFDkn0Cf/eG8QYpnSaFWJR9wHWQb6ubTE+w8ql/qP9lHepEKyKGM1i
mGug0n7W/BZ+ADLAdxzv0IKm9NiWJBgNDaroL84dYuQhgUBP/sZ1bp24JddkG1ab
A4gSyIMU5ludfMJhuw3fdX1ckum9Y9dAIKObDe98+rugnPq04HHxbtu769iOZ9OD
fDtt8l9UifHuIru8Sl9B5d03oW7JtxMo0I8TuX5XRPlMqcRMQR5JG/pyj6uUopmo
6L578qCsbpJHZF6vAjN+ZnvLMlOm8zMkboqQt58KjpmzxZrKKY28v9nx/ys2lYzt
Qq8ww5S9nVgRBg2eBh84o8d1Ng6ptAYP+kKjKsWguulqJv1DCzX9S3+sH4NoaVcT
NrKONy5urq6PaygoIMED0nVR6UlaehjxnSi3unL885wa2e40SC+oCe/JTqLOA5dI
ccBXjMaz50aeF0bFokbgOHBLd2s2HGAXK3oFTilnRHM1cYG1qycAaV5dbKcGE8ib
67hLY5OcI0OUdunPl/TMlgZreMSOq/q48ab6pncRrvlbm/vxMVDL/aSVNcOPGlEk
kiUormHPwgaWwvWSTJ1uY9wWvoDcfvnDC2wW/X4oNoMR358GeOtWgVpuxB3UrQRS
Xr6RvHa8DAdO7dsrHMalBton4Rwmv0lzUpWMnkvnZgC1RllD2MZ0AbwVD3TwEUJ+
203QyAsEwGPoLXuIWAeIkyJepVGExQr/UnjwmlbfM2q4hj3nBbpvsRA58r285P7o
Fih7oQ7JQ9ZNfJtrvC43qP6Y1a5qOMesWVLEBwpZ93i/k0Yg4a4vakiHr27jdmH3
+Qkxy6CrhddOSSOkDkm4pmW20+o1e20jKCP0U28Zsmi/9TL8tDU/eI81C90mbEp2
Yb3zkkqW4GoE7cBj2gl+zris+XXQibZVhF06FHvbSfzz9Y/+2TYeAIenAgqOYul9
E+C//0wO+M1COSDKt9RVQCoic5pfe1iQSWXmYxQdbdU46XGPwwmIoaoCe5GhIelI
43NrX4074gryl1k0ujMYjmk54bfnUmrd/u9N3Xa3km2tdUEx14rSLQ/oozjA8pzh
0G4vHmzW2egY169fTARvTO/pKA0vGPu9kkqbFf4E0ZOZO/qZGu1Bblj7xuYdhEk3
noRQ+0wF2UCuXizXcEq+5wrAQ9nG3z2f1mRKIdGweaEUwPySLANEX4TK1bwvpT7p
TXdXxJKhbrjDM9+SDAt7Z/QtAXcBs8DaFRlqBZD6MfBO5E2I4+Xm1RQEMRDTR9D4
+eeB9ADzKu5kx52g+GVsqKhrxegVHqlCQS85JneqBE3SnhNwLDaAKt8LNWKv4NDf
H90JzUptOXpsunxPWrIwywpa/0X1HrpwIBtj/ElEYm3MOsYCtbLQWVPLV6ZxPCAH
wdBxUt+VfWzdshftITF/4mWvhale+m3QdSfn7VbUt3SFnBMUe4OgjcErg4VzZdpp
q/pvendQoY+o8FEz8z2vQfsuBvUxA7mRgEQioi7XkbGwhPnVxFyCcTgLG8q+1pkz
EAwcgnI+70LLG/ynCgulvArQCnBZe5tzeugrjQaFLyUR0VUDqrONSdR7uMjky1Iz
/Xzm/UJ1GuPs0IHzMSrSVSNZC6Sr5hORNTZJJInxGcgNwYO+5PwIntI+AB1sLM6Q
BQMEDfIJ+PlwKlkGFXzu0I7oxmSZUAqCwOD7mh6oy0YHLmvyvGQx3FfgEqg/ydZi
2dDSWOj5MZSWLIc8d/YAci6ho9WwKJ1koPAaKV9uPJx6xpmw0ctrF5fx/yL23RkC
WsaplppXS6ub6w2BQZ5YpGdu3fl+s3xSP0Su7HV69otOTGDQ8jrrZPjH4uhxRumI
MdfqqdfphEGpFzPl+cMkc7x+OaWY5+Y6XAHgMJ4yl/G7aBydpK7pi6zFS5Mh+icV
uP3BDhmIL7RU6d4TiFUq5qCt9gk+Fe8/on811r5ncLBLgUlVdBhLmGhGHcOHb0XH
9J6kA1gHrbgBHzmNo2kSwdBg0A8DN7uO2rA3N/06mkEGU2xNnqunq4QY+B6bxcm2
rKkjQr+iS9Y4LKq38fAhKUWfgFND3+mq8SlsBPayb+erk5l0tRG7AAdrjjJ0OL/f
0eqps3rYzv0aEbIDIYCIdNUI2wcYRpxULnSLjJOIm/YsRon750rPAXpfO9znxSPH
tCjK9+MsodbRMN81vVJIt0df3LEJkYJ2ZtwtJvQfFfB4hem07Ovsk6wJjb/T7+5b
VL19zLBFsGflYwhx4JbmBLkQtTeI60ItBI5YOadltvv9fhq9hgPUS/w76Tvg86Aw
3NHzaul0G0+/7e6zPv2Lzvt2PnTzdbyOIcFByIdNo8CzuupIPO42qnddC0EIwnFM
ctLvh23tNY8HtGtTX38L7gjBvX/lV4B9iYS2NblAFlOIWuOCV6CYCXtQIzEhrN1Q
tJDl+VoHKANok6MYHBOiyb0AKx42sft1ESDXqJFc/ZtRaIZIKpm/Q4ieSWRh+gP+
NN7eznCD4ayhXoHqPCbX7faiWz13mxJi0o2Ni2Y7oMHzO1Y/Evr6+3ZDlTSwh91A
2zp/sSDMYmVFmsuBeI2D+cc/ThDh3dZTF1/Ymu/q1zHVUnISFrHJOBimvUyDe7Zz
jcWiMcx14hvUl9kirXzjpDHy4zdJyCPzVzK1+zlRUA14eJoD6PB4xYvlw8KZR2T4
MNPa/EF4C28vc8+RlnAdA6m/U1lureKD51QYYRdrA5e3vUVzLgDXWaOX5IbNihUd
/EVlWKa/6mjXqUN9WJnkK3FY17UTi5tjEYLNrd4BraUlAmUcFigVH8F4+ZBurfRg
SPSfuufl+YsDmdYpcLAGWqv3XVsP5S+/7wh7i5yKf69oJ30X31vNJwXTKIq/o1E+
6LOGvOr4wDxVh3PpjtbU9kx4rEehfLKABHJxRma/MaNYT+AVD1nj0k1ZsuN9U67W
jsfzOqIcs3R+h557WUeKBmYnZLhlpzLpVD69Ut6kZIGY93UJoB1vLeBjBsSiHi+M
Nuj5Mll3rNnbvGa2dJecWTgX1XCEEgdBoCimtCxBbh1iunjHU6lH2fctvue06vjI
B1/Z08MeWUaTqzwMl6SJKWwhV1Hmb6lGX8Kl4Y2MYdKwo8D3ABe9mcZqa3oKh7uN
uRlA4RoqyG4QCnpKzit+reEP0MS1a2Y8x9ihjMBjPhINP5ZauIMuX/HmdMdfcTCY
51eq259Dcn5Cztn7wNDp0jf3/DBkui8kq/VLsl7bIZUPRtmrNtdvHkPwXmzu2KNL
BNwpu8sTmPl0klqVcCvAQrnvezoryhLfzvycl/HggUJ9wA1NhE2LUihxCeBXGLpN
2oqfBYXknn0wEaNaZKeMbgebsB5+aerzAe5QNEIKCAHK5JHonFEBQsUShk02KHvF
4ysIJNanWgQ8IcviUlg9KCRw83v8hKAFcHO0DkrRQmM3Fzbq+dobW8K/V7psDR09
pNnDyNfvzMyxxCVgT+iaFmhpegB8uflBl4/0Ky3ZK4MbjeJ3sGImqf+N6NQIXQwI
KMv4SKVmyZDjmRpcCjf6lPz5R0ouvRyit6g/pJW3uZ9k7aNl+F8knwSUTgUotGd6
mK4ENHPDPqVQeocDBwKKDwXuYR1KbkrpCjPUG3urdRjbnF6MSB9kWy9oCz4UR4KI
+HiVwDoN9Ajbvj85njkJYn/OSF1verxdBXfG9bvp+tiovppgMjs3Vq4zaq5IjvT9
rXOh/9VG1/zx+eGHbt+rQqxrRgZN2P4fqseb9mcWVgEI/jWPeaWKv1BxbIXT9Pgg
anjU/sevZVJPyqYhsnw80MKXxe3ZqZ1FNof0dZVw2aMHgVvjkfqGv+6oZowptyEN
RlVUAkA51g7Kyc0F5xLKJK4QBqKiXq7+SuBAF1kr7xdfJDY3FB/wqTHD9Rii9Q9f
lbIvjIP7gWlc0BswoIngxCuY0LNAghf6WEn+7uPMwXjtMjWe0H3tj8qGBFhX0Q2F
3k61a7WgK8H37c8nXoAtFIJI+sMZvcr75M+a6oPQynVm4i3BJNYusUwRo4dlewIF
gpCPxPslD5gt5rPjL+3BL0Y4R1UQc/w52ldoCcAeKo4inBsuKraGubvUp19AlodP
uGTjn9vKkRuCrP9clcVO2Q2Ne8OqH25IQ/6CunNjCjmkGgZnHx1NAGT7EFg+s9WE
KKo+1PWcNuyDywQ4y31xU2I4V+tDF94P/paHdVUf9ehQK5KgKMGJf+inYKKQRsWH
VVEuCKL9dHUDB5OrS4hHnvAlq/BzwS2RPLqygcdvRF5b9yq3qTZR41Wj/tx5gYOI
R6w2eg9uJoJTmxj8bQOKCFgFoNmJACd37GKw9DfGbrao0nDDaV2+448x5crmCus0
lOFlepz/Jl2FSaaALipmW47BpkPxeF3nTy0MMEI8c3yNGp9mN/tJWDrHE4X+66LQ
AZ0v9lZCkpdhXJt1vslnj4NEhkvt1zpTZa7Mgh6RAanSVRWwCD42J006NW9dpd9U
lI3RQN4Oe2CdsABPSIhWAhpudUq28JzJMMvNDjrcaK2omIqGjUR57rFR1Js2kHX3
r49zi1+oZRkzLPJnFzgeOPtXA4KTddEhTjOUq82Yztoe10e2o19fhdGSivM5J1ja
J7AqeqIJhX7f9ChvqedUL8m/6PNz93hH3xb4fMYHeOLfaowkDqwiXf5B1EraW91E
LoLKpvIAF00Hhpwev6X/dovRIIqqw0x9B/pQWMHpkl+UwOd1ovYLp2uaia97nWJl
AmxQ1jsVNXDD9UZNSenINDVaZksp/rah0+deaYFl3gFdDsMvnncWr8eeBG+nmKEB
RMvQ9xgc/YZ/pldSemWKjZB5SjfsFEipIKw80XIGvmSIXNbbz5kgO0G/PF4JVWUc
+RC1gBJ9OxydklpvZ3uEO0wDJXD9PGQWEzb2BU3zBn9HzOTgWcPmNS6x1vGi0EM9
+Q1eHEXMJ5+5bI9lVlcn6MuRoyLyFAAlwZB/ao5PPWxK1dTyC62Y+1njeACfZh/a
WTcok5TrO3nh8rSE9XjuGk/cVP//u/8l1f+SfNnEW4z+mMnxOhd7Up54W+axzlYG
JsMV8Pi/qDEmivRKv9h+PztVLDqtlhsHD8o/7Lttt/utW1UGbmGv+5HHTOkbrzKI
KX3pfbRFtmjP8katwiIFkVZN5l/uzarWGZ1/a3P5fTQ3yhZ7mb3AlRghXsMVo+Qf
7hukJazGLjA1DX3NBuJPCJDdCOhe7JBiN1nalxqG4+3pgoEMg5ZfFaqxxRSMkZx/
jz+6jD6pQZuAwNPj887R0qpifilAVAMCi9VIBGQWu09EyRTblr91QrRCWhMldv/Z
szRaFJ7HR4upIrPy2W0l9hBVE+qhFcxMUNRiDaUGJhTnThjg0OkZkcMgfMEHCwDK
beEDrH1sYaWOHrImWxTay3IhIpUIECgW5mBRueS1qIepvWZ6CBLB7/iaoiM7HtyR
49asXNx3v18pzXcQP3TakWEaWtiLZrp9MbHhakhnigXTyHVCpEoMPNZ5IQO1zydF
CMxUKDUAQBqcfSBm2VRtY2RgjPv7L0J2wMlKS+2iMASbG1WyPepHKe25/4h2kVhA
dVo7nHTkraxaq96j/1EC7aHDK+CjnQ7ybAwMxQub6GQpGBDOY5TAD9QDXY2rF37I
O17Ey4PtI9MoeurOC/tMnUSLs/ioBZIr98aPjv1C+KiJPcSFO6hRxCdFNC1Kk5T6
Avx8I9jfPpmPrDOxrZ4/Jt1rJFar4I4vKFanzkuOFGanlLK0k1dHZgIPcutdU9RE
GwNt1SphBSAG4QaMIIDvwi4+4acmdff3WQXwCFUDIhUHyy5AJ3Js8si/uprR3mov
bJmw3s0taGEJUCKUJlQO+AF/GInuJVYBpeqgkE+nb+g5uK3h8da6Awkv1hSMsa7x
tizCTxom0E7X0OIwEgeUZkzEmPOdNGpfmhI+Dmm1STQVeKj1qIibPcQRYR3w2JE1
P9P63aLXEm9a3F0K22hnvSUo9Me1XTFi9GE9qpCTLqNK0mKIwSn4L1dq+KaAeo2F
6plQIceLXX/4PPalLhlWhLsIzkT7Tbi8ZtmbikTZujRZr0cOPmNUxciJp1jDbnSJ
SG3fkqn7pTuQkvZ8fXHpvWO8ms5wWpDkRHm1az7v2M6L/2rjWcKUVQH8IX8ruoxI
GJOVPN9acjYDxIfFpcr60jk+l+Nq4iW0MTNnnWwqzHRB+hsGwuoiilJRpmHryLWB
Po3xAj1GrUeH1DAf3km/N6THFHzxqZRSzEfGtmQIFFScQxidSTdmp0WRIh6paAJw
T9Z+e9MbxoxXTi8W3kzEyQzb24mBprtJwEtNWdiiVvj+TTaUteQBxCUbbcAkd9Th
foWxo0taRh2Sc3DXGBpdv3Rl7sYW3HNgCm+Cw6iuiPAPQUZJcFdEriq7zF9SakFD
kIgGC5kdGb7Ien4bg/e6/u/+kuFM2ykbKZIeHTz5Ho2+Pkj/P3fPy1fwSuCs8GNi
HhjOqykIwaDAsY+4hT+zxW2SI8wkdJqLTC+8ITzzc4STUhs0w7MolppaO5ftmMZA
6+wOQhw4VBj6+d+w5h5AFBzU7XtvQG/f476S7TutQhEQHxg9DtZSJfc7JWGiHIMl
MH7Z5u2FDlF+lb0hetD5E45YsaWK1cc+lLWInP6wkO6NRiQxvBjnZLNDJ70Xx4uT
UO7QEVJSsRr1G4AQuIffyfHnYbHSfuk4yEkE/sbPYhquJGYZd8kfttN5DW9i3Juw
8ufLNf6bMgw43VX0EUIQ+knPvMOOyV7IpWkfLIZVKglJojWaJ9P45KySpQ3EVMJU
EUGNtvF9esJ7fVTqaT9KlD4FvgCmMvTtXHi8VvzlopkH5E2aGoxzb82Fyt+1YAy9
s3dY9coZ/R02tjZ5P30kdWyAPAfS7vTETOCI5bsSlK5eR3xEZATereMQMdPaywWp
p1U6yHz+ceinfGjOl6XzwF4mKwvBFpZGQvFZtVcafMpKJ9BrY/zvZBwAbIqoxjf8
T7ihhuvS4Pm0Vzx+JXI72mpm8B316940xiKBflhz1oy3d0a8/rNof7KxhgU3B+9u
HILzrCFx+Ja/DPi5+453AZj9ZQQQV4/BQFpVVneKNOQeRuZw79FYUHVMnCRHYDWu
p7P6KzBR3G2toJclfKCCh1zt8sELppgMylCtaL9EwT1rpN4in97/qI6tktLmgPI8
2283Tphucw35RvF8x7gUYqXlkzu71F4DcR3dggDXncWUngbjLummfVKWaFzM5e+r
3mby/L8/4/TSVFpG+93lQkq8f0nrKCj3ewXzloo/alGpx7IA50R6Om1l51jFQmR0
kOUGURZY+//Fz5OgWArH3924SMqfYUldnJhpJSeqh+Q64QH6ZfuUC4bAd8sl1Imz
k0kvqP5LW5yFQr3Zn6cqAWj9B8wJP2/HLe1bLl0n6UMawHuhnq5gEwV374JOUQIW
nKao3guUggt8FgaTKFuH5SuQA7yc9AseTg87fcSLx7CzeT4m1n8ntH45mZJtr4lc
IFtGX/P+fC/dy4ZSphHlNSL4IMsl+Jsd7myd84DtzAwaD5+0cvJg9UjCQVVvdbEZ
QOkqMHlXmWBKkrHlu2QO3O0TrP1P2KxYumGbkpL50wgpDc/VoF6pMs9p9/4mOu8m
Iwc69xptn3u0VYfHjjXfJu+sAjkKQRysMkd0EvLlXCgbKCMireayytJ7Og1e/HiD
hD44xWa9meuXf4q69Zhv+MtL1EdlEBVa5WWmZBFW+pxEbybDXjca85xpBXFdFwEz
xND1hQS8H2NPU+9RnD3RfIHiq5ORSGwlExwI7Xq6q4a55TeqEAUvDNBUDROVa2Wb
PAsoiPYmCY9jQDuiOzQNLitUJ9Si5Km/yuCtshaiU+0MU6Ok0GvAjGBV1WNI8GBu
LUtQaJCpgaQrymO0rsrnAIsmMNI3eTS6OccjVNUKQ4mby5A3RDP+R/6DLwy5isvg
KBvnKtVyMiE1oOTLAnTJpNObQqon2ZMZzwr3rbNeM5q7/NIGWPJnzCzX2rQdezfC
O4Xpd61GRkKh/cU5mwN4sTEzfpk9G94IdTMmHTtDyEygwVhqotJ5+c6f+tKHPsbO
BZ3Cg0RtVufLOn9NIJkjfxHj6iBnb5yomPJJsMDsrp9xKbiKXhsKY9Yik6La0DVA
GnwlZeMnX7qbieXlKt5xjhTLdI9071OS0h27jVcjKZWr885HPcQ9Zg8ZA1rqIBya
hWXhz+AarfgAldEfRNZ9bUwfsTW8+lPBIYX2gV7n+Fzf0smBLrK4FF+U83j4dEIH
NH+7GS/Xk5oToC2xqMF2xhYi4/9r1oGYFjYGwrwv7b5uL+1jaSH7ZkDSFH2UTrsn
/eBafLr3iXLUbh1f1ibYS7wAHgC5naXfn4ZQtv/JkTXdH0IEV2FxEQa1K7VK/XdZ
PjcNyz/RUxX4NQsA2V/ikaULO+APsqKwVeIp04VGxeNsT/lX0MR1rqW44wThY+Xc
rfsY3/g/7cpFz/nLvZQ9Ej320v1XwxhBdBPiF9/RJdIZnLGBkDoO0dyxiXkmW0hB
MrgCBJOf3idD/IPHqiUWvxPCluWgRGUyD2OmwStVV/fRoiumjQRiFPtxeOIbDMg8
fAd7jezgIHFyGqbe7QKHlaUxszOYji2tH8BIpoceYDT/tApJBAYfFevUi6LhETfU
/HA82ht6X3+y8o9oCYXJGbqyoXwin6a4ytRjxdA4q7pGJu2pipM4ji4PwmLhr6sH
+eZwFlbzs12IdTuiA9dbHs0oxxXN8yqwZxynCZxC/x7vey2jRzBD5g0Bt+BUj3WL
HyarLzqQCMflTb7aMjXeuvvlD/RYHC4y6TnCka8guLNfjBpJ9EKMY+xp0x8KvqM2
ta92NgUIaNTacHg7GskZBX4UD6FiIq0H/YNb/B7n3HNkFLdbYTK13dxdEZ7uxCPw
ZqWKVu6SEh9h14ljMpiBCiXxJg4+knVp33wLWNPH6b4cpkt53hzpPrXxxgKtyCrv
6Y3a5JNXaNdBiXqgiHAW6G5zRCMXfjNSTOnBE3qkdHVf1s/W64x05LLVHSGU766e
gKyAWCJYsj38v+r5CVTNdM2p6w9Rci1y27NWQ7HySNcMdmk9aIUx0OGLMEeb5kT6
cYs7h52e9AoAvYuCBiwhilFYTJ1ukWkcHdevYzXDcYuw7PAw5sLCAzWhABgB5TQS
hWTJFHYNroU6tz8X+sDN/FADZnOAkYFwJPh/mB21FdwKEgIExMQgMzBpbRU+Lwou
2fwQjyzt/NN1NfFTyBiJMwgMn8x9ZeI+nf9vCPig3UeLRQtYtHFik1kimrDsvSad
M3BY0gklO578r+wCLVQJSwDmaNVV5KDPD5v0njwOx4zGVIh1UjZ0kneqennHk3CT
h94yk+3pzv9J+kzXjnOefHHtDbnqtIEf/KF4Z48rWhupZyUH4vmUagF9a9Wjmiii
i3L7yq5v9XZw86oXrGlY9YkZ+FFRhwWems07BzAoyRPSgkrJ53N26srdGDd0KIQ4
3dL2Vs2ruz99DylpjULHW02AGu15f+Bb5Bnb9MjbcuACtg+7lNsNCKOMJpBo9kKl
mX5ULeXpbAb8sH8NMSfQHhL5B283Qr3kt0wtTTLKbbdIAOaAIY1Iy9010NTO3jQj
1dydEEiBWbY8xqGt5Y0Wg0nwFGmYD1tlPN/lA/2/Cw2VNzliTK85MXtydYBgU7tm
AbQfrXkPDWapcZpjJPY7+FsLI/vJlyba3I4EDwOFfU3MM9Ch6VuYP9mdfM3Jle2R
jAI+QQCPdIcfWP0jJyqZsWMTvUV3qAP9zcrGXssx5JU9xjCuC9jGjikMJ4qvmIGs
wgYL576ZqZxvQezp87roKbUPrVqOP1VbzNEQCysg/qoqufk+jIE8AzR4EAPZ/Prn
LpG5qqKr1V1/0715Lds2N8ESRjVOWzwjXchsks3bse4WuiqenNpRlCWQXwcN7Uiy
yOaCk+3Xt9VBBJS5viyq5+Az/XN/yepextx5+BJOCpEf2VqN6N+x8dUzl+CEFY/O
uHoVpzFIK4FRqHVPpmRAdgRylzJCjDrCNjH8fI9VY3CW5zdRG+vYwwZzfEJzeppS
my8qJsy1qR0N77NAv29bLbesSAl/dLWMqVSOIstLjc89ZLdjAnTgwQ5e3hOYXZPD
HZAEwWNwcKQba0O2W/UXO6F7BOhA8E1WoUZ21xdhF7Q/DFv6IM+GdsJPObaPPMbL
s1N4rPiaoWbWhI6ZlB/flHxL7topQyQzu2wvLs5irCHgwsthTREFie4mPSyB6ipa
h0WWZIfu9ZZW+BpsG2gL2ETFGl5n2prtyiTC3S6gnfVrz7BvKVjKE3xtihRLtZeU
fsOx4l2oxDGee6r2OE8OLKXlyyEnKtxcq360QZz8VHs1l+swe3OjHOzEtn2j4Njo
yOiEoxgdyD60EhvGjmVxD/HVM1sI/zD3N1vmzPtAp5GU68THsUnjJPyYeVsnsfqD
K9eKWjYUUTeqG4s16MgCRZn622hHRp/+ifRxIHC6uq7oXW6pvwHrartpo7+dd8C2
hOM3nPMGyUC8qD0MWJ9ZdlPt89WNmIUJ3W0tjE61C6H4/Jesy5RTR5gvKBuNdbG+
jHFAKhyhH4SpjHq1cE9tOQbVAxV05CIPcs7O9EsH6xVNjUolbSQM3v6QQ2NW6z0o
qehkP77DjX0x4GaFhpACTVOxrc+Uqa7F+wQ3ZUxyEdlH06XYchCohnCHpbZ+l4oF
Hd6oLR8w5aqDogB+qCk14A6wuglNcgqSas8WnIsnk8sMVlEufKqUfqK+sVxdeUeI
U4HGHniqCHH6GFC7AZwwdLw5GcHR8yP/JBIRXsyDoVx3L+c2LR5i2bJti7Ly/4QL
r4B0dkaDzs7YjwL2ETJC6dJxi7GMiakW8Sxg1ekrqYJgJpd8koaPkyTaOJqgvLpu
3FDut8ynAzet4T99ghZ0ckSG9oCofW2YIvrVEKfc560dvM/wMeZhDn8fHpyJm6St
lxNMe+h4mlCNQuU/ntzbu3SdJCQ8lPAg9lRPzKAcWLWevtxMvgoLAoRytUnGhy7G
GAYkkaV3psS04wpbqw2KwUPpz+BW474GmlqigT/5Gl7yI+kPQk6f9bIWplrP7HeC
xK8w/mh3qfBo0u4TzhyjWHA839d7x5RZOkIBR7eqNOUxmZdsCUZyYl7cs5dfbXZI
00YcTyJ8kJucxk12+pQZN0o2GS4gB413mtzXcgjXAT90EDwzsaMFMuwdza6S9Ayg
P6CP4L5Ui5TlzoO0v56ZPOwCt+Ts26B4928AWGiet/m6dS/18HIuHg56MxjtEHlF
cvYNd7g+VFwskobbZIb++SG0aiyiMOHOgaE2pMPfettB7IfmNO7sKc/Ed1cIBbfC
96enz0PRPk6ka8PzHSodaWwcdvX8X/BhwtlRavSR1nO9u8M835mp1Wi/uwIzEPCQ
+QzKcrGeCPlnnc7el+0ltRurz369dd85tAGeLXxljIcrasPWQpU1KrYbA4PXhTN2
+dx1NpEucWO2jTcT7Th8bl+J8V8iTbbIe5IpIP+wJTbwIwPwKZYCQtFm47gZscPX
LEvTM02pD6emvskMMHfElYd2VADdmswEov5cCszU9yCSpFvuPTgMDQGWpO5wWWxI
CJM1cXgoofKHdwRMHTTdP+LjA3c/YFRwRs/WQtzWwvhpG49FpDc1wzfpoaCI9ANM
9dOGcJJ4ryLk13NWmPFtZWIDz83WAFNotumGlEMjCQjoPUTgvsRwinQVEraRu2Mg
aUpWWhNesRbZvZWS87AkFkRbsedrxLC4lC+LYt+2aE0HVRJCUYCA/RzpTaw5NlYN
4vHN65S73iI3eNAhmFaPT0YrLvFgjCbpcb+ibR8WXhepASUt1bmJaPwzuSVHufnX
RThSTHHK51SX0V6aX6QpE+vPWgj7n4DoEFRLXgLXABK0uDbm1ibHFSdEujv81vOO
3tq+UNFMkY66uJJQBah9giaOpY610T7cR8AHvg3wcM3xPZMXaF/VUFjuTJvRQAAD
b8Pr8g+L8A43zDNEaOBNf0k4qWHxAnU6MOxhmOfRAa5rt16J4VRAYIZDw4wK84gc
VHWJ2x5L7wU50Rn53S547HPRca0bPIrF75Ro4/6yGvA8Thdeagali3T6eLEsslr/
6neHz5NUMZarhJ1xW1V7moz5w3f0gMGBMYDKabB8GvwX8my3plw6unIbkp10Ot5B
mcZtL7BqH14XBsMgxwanmnmtORZCHcEwcFAA7GmARW1QYCwDvfvbtOSqLLyLPQKQ
i1wxjdnviYYTToXWfxTKsjzbVzrWi+rhAjkjmEQEcS7MPwHplTXKSjZzGRa+wbFN
UO0tg7y5DjOybIN6/Uh3F9y9MvnyCPmFtpveQ6YY1yFA1QhxMfPCSXIMFAEY8D85
PVv+3ejKyMqaGOltOuxJVWzASecq6CqpJBOuDbqRsOFs+BAFLpx2Gg9MK2tzNF9K
SW9VRGPdnXM4s5jvKUb7/g5U2s6/X6jyl13s1V2f5nzF2p6x0vD2QL3UmQ8jL+1n
9mZRpNm8psJf47jj4RXsV7fDB6wNPQyd7x2u1ddo5FfCaPG8jFtIFYigNv9YCNsi
U7kjBNq3UE5Zw8hdoMn7RKPPwGAjQo01wrAGkZ4pNiRxN2g7h6IbwQKeYK9pSgxv
399EodQvMGZ7eYIllZaq2ejse28/DnhZemJMAjm+uF/spr4D25I1Fp9fwaN20j0o
BvvvqzNA6GjjEplbJPzaHTOxDvhLHEWPtIif4UjyKG3i7pjmKOZVhwAACZBaf79C
Rz9esznAyNj2YB7pPPaP0HCXHGbldS40OwFqRvL54ZkqM4pEmsruc6BC11fo45cv
Czj62N8hPX6c+6loDT0yh0880qBvypJpSpcfLdnBlj2LecUXa4g6dVLpNh9UNdZm
PaoieHEXmudsOEXaMI0v7fEtYuRzb4dUmo8ZrEP655VKFKt7AclQiax6IQQkjKbs
gTuFSpLMR+O9apQqpXeOe+hUkR/hjfz6MwWTGqleRJ+TeuxNIZYnf0x9le50dLID
id9d1Ch9kyjQqLI5O5I+BwNoi5+4dl9n9mulfqJ6QZMneLSiN/0+0G4PhnYFsTRH
nYUQWt9NGH9GccK/kkO52SL1w4OlxqtgxH4qDj1RFm4BkhAdlo5Ou1pukGC0Vv1R
nUcfCXHBBIklCr/Ti8HD7rvGV+u/tkgGufusNq8twGLVz4irJK287qP2zv6/pcYs
ntd+/5CoRqoGRTVRRjbAbq25dMPhS6ZcIfAojIAuFN6XpXHK/NGomnM4lQcFgWzd
JL0UVQNHx2PWaMg1ZCQpLXDxQc+d8ssH5dGMDUNn4ipwcUtYBpA7TLACPUf+zyOG
m42rByTF1Uq/cST9fhNcKobaBu2iTzxXFhvGvocV8r5p3d7HGR786yc0G5cxev+p
eBba4hzQ66iZvN8bsakFFoFkJCTmpfMwPRaN1EnU0VJT34A1RepuwW96s75LoWZB
IxW/2gK4o1L2zkyol7rOu2WeB8+tU6YtTQMDDwQLreF1U0mFyDiBqGpsz/wP5ivR
HUwJiCaOBxSDiX5S30vB1cTuE/0lFdt9wGwDjqbCxtIhJNr7inoKBALk0riAkCfR
TKVsM+lbqkKmT2EsXf6769UD1mizqbh7nZbRUiqLcql9rhFsHZk7KDI4va7sD+0d
f05LadY2HX7NyrdYIynfvHhAUe8AFhdtVoKFUYtJxmV6n2bwE5KokJPmDJLLksPN
oDTxy9oaj1HwDAgN0y86iaGrsqYNaU6uUsCyUe++2X/VJa+BcpEWZUjxtNk3TH99
dcPXmfuLcoQG78RMLA62oms/9MnKkZze96CnrPbgtqUBn1w6seVoMqcXVgVoJ9hg
6aGz3ukOncFL+hGoSCrIPFdydG0FJBygO1ovpDDBzFmhlYvJg72MbvA6CsCBKsrT
at0YQ6PY7cYpWJotySCPgu3ySfGCldLXQZfp8ywJbU4LJWzsjMRbbz9cG7dci28t
I48QfBWw84Vv3WRyQxgQxHb8cvlE3/cyeWr61T5/+pwbIih2qSevH3KKSZRfBwFq
FFrILEaL+tay2ZS4MN/deKMUzqYFFJm2ClkQs2VYXQ79JAyBVnEK69UoLRKla4pN
mHFEZnoB1HsIc5KaTE9InNBgmKSh5YBBljHy6y7dyWLxxCCi/mpDV16yPi9pQfHu
TPohzooDfZ1LSkIgsHfKUnupptARf8GrZoOYBf408CX/QAy9f9B42tDB7Bc5ZJtp
s/xisGnLq66FBSbE8TZQexeay5NZ/b4ijsOAiMLck923DHX+3qXE/4veQIJExGo+
9lD0V/mE8nsd4CNec48WfiQ+21N+jtSUK1b6wxcWLEat9bRtLocca5JZEkDjI6+i
jMK4L0AYwAZtJqascof7/ymXyxfsqIppEg3Iy7hsTfDW0tLY6ZUkHlPe+MkfFWeM
StA00bOC5o07316cl3nRv/r3PNzOo/zotu7c2cmeA8k8nmybzrg0M8xBYsl5Y09X
CDHHI6ELR55BzI6kTUtHhVK6QeuwBZEA3fiP8pJ00sk8/Ph5LaHu3IUU3KVfZgH6
BuQJ8/y9spA09LPxcNzXzlXIt4JuaAg9xWcCvnfW6Ucjvs/3Ghjbgcoo3oHbEIz9
1IfmETUXAIytW4SY0i0t+PbQ8FZquYEW/WFn6fVNrLtxYxZ59MBOsAu0d0/yUGHs
TyXNi3Tsxr4qCLZkq3DAPRSBAecfPMEtMEhrxPaUQNzJgD026YzljwHuP4kPAp2n
QAOKTB6n53ookkicURkEmLjGCsxy32pEBErTvTLg/RBpSEbYxNjxozUy6QvfSyht
zyXk2XW007lE28UsvNA48WJEPRFBxop3Tgv/DhpD/i1L3WFWltWcheRqvIadHRzd
3BugOr8WWfFgTBgwNXBZmcv7RUKzvOL3hP2Qu3r86/Melzmx4gZpKbUE/bR0Rh5A
7vJG/GU9ACloigTgRGODOSvMESLeW18x6v1pA/zxjK5IMuSUHtDvSPyb6KZosTlY
PxnZ7K11ywUqJ7+l30aponIfqsjWtKTFb7Xxqx3WBSE0lSTqLy3R41QJ34NLWVAj
EmgcIq3x5+bJ5fEcEY0Rf98jbXxeqzjEtAiMds1b+PpX9HgM0oUHUtUfr7cFCBNa
Nm6qWi8YdYENuA+dTUaCuMZd/J8pp2m6uOxnXMoPVn8Xk26mLrmjUJAqvqmAxFIy
BeCsJpOm1u17+3pVUwQnOJeTWgYLRR+RiCCk5SEpsKMR90jfysKDIPpUogH23slI
mjlGmkjfoOJqM6O78NfTAyhlzujLXkkvm8UBGOa1esIewV0N5HxoIjcCymUNJ6E1
MwLJ88vhKlo38AHtc0a544PZ2JMpk0XwY4wr8K+6Q2saG042txndP3i55wCY1uuQ
j7P1QLJdOI7s8wwnMEBuXjkllf1xPPY9IAakAHzC4bEsJzuS+bYI+sZs32tgCKOF
ayAH4klcO0gVdD8BlD8XI4C3mrUJIx+mQ89jRZuJ6NZXzWcU4K3Hnq8o6hFU9qIv
8afJoFDtlYAk+iR89DKSP3Mbfz2SiJYHxGoQDius0YOk9aCvluRLO8tskgdb3mmN
6nyzSEKrR9BFwUHzUJamvBsq/E0w2oX5RIXa6zQU3rjAodw6PVtIVxO7Q+NTc/mc
3zs5g6FAG956GDnSSl3+UwNczndn2B0eKcxLhhTWnPKjbp9t5COP/sWWxn0chZWb
g4+S7X9nh/ZyLHjzwnE6wCFUddjSNFXFfpdYTrFD9M6gm11PB5CORYs9I1s/8urh
CD6C0ltZeN6r8WwHqlHFdkbmaJuOgMTXld2fsJiLzuTFGaKO+0VuqLtnRUffb4Ee
oNCZ1U9VpSG96jcXtsqcJcnt2Tw4OQr467S0FjL3Rrl3+o6L/2gpUPjXRSJVfBWv
AuksXHOat5B0kjD/9xg2zhMVM/Mw09T2nXwbvfkSaZQ7qm6yoizG4O78KPL6HmPD
VO8uFGgHNDpHKvdN2UJ7yEz9IJAMh8pOPXtCWiqmRzrO5mIyGVwQXpYDRweN9UaU
0BZ7Lpc/kntxWl7pzSN0sABKTMCbhxEPwjOOwkydZdLYwEVPhKwdeTZPVTKur/bD
Lb78BPDajqd2Rpp7fMWr1I5R+YzIOz//zGqsirmxffTtyCVmqsZanGHlK2O5xgAy
ZdkqutcEXXDiepaR94qvzYr10IETuRAIzT80IrmVGtQMN9s8NQ+TDVNlsHuKIzCe
+0mmcgj8Vg8OUfpzig/nRZcKf7v0SCUOfRzuKEOlA413NvGQWAoFWLg9/lJBjv8M
Twooqhs3BT3pj1bkcyUZ6H0G3i8RI3FYIjNOXZgjnf2Cjmt2NtTn9T753dyXCOs1
rzNh+1tGpghKtvsuhvcwB6959OPCa6h15pnEG5sqWXPtOvcaP9qUDYJ9WOOAlK59
sb3Qnt4p6SitxeLVHjTqDT87/WgADxNXS8XBLckPRc9NJyDxxAdGN5mfg2EjvF9T
A+50lPBDAvQWNjH8EESML3LG3cTGHvnntTZGEdsZGX2GoA/j5exbKOLP91jhFHBa
Fcx2Jh87vvjzMPGToK4rZnkm5jfQ7je10zPB1RuFnCEAF7tWwbAPwDYep2+HqqX3
NZLztpszWwDSioGvvhtNvKGDVY2nu3JpwOzuSdYc3MYtWsw5buJO/JacF5VsEmMD
Tb7zRCsJV2NBpmExRkC9EPQ0YdK0Gba1xxtQ6Se3g5kz8PFd+6e6UW9LqOzc5Jrc
o5KM4n9Z4/DsNWoleeCfGAqcr/dfUStB4fPFMywl1P+Jw7pZy9d3d4HWeS5C5Hef
8msbz1udcysi9kQXvjI6YUKuZ+anZjVmbM9yySQ6/sRsHsLcai8qyvU20FrXEVZ+
uQjGw+bBbU5uEL2d4vm1MvFlbxIAvv/qIkSduN/CwUoTpIslT53jkPGeVPnLroaF
bVQ/wMB67/99pxIyjC5YDew9eYGVE+OJ5hG2BECGexb8ouVCb+spkRaPeahqq3lh
LIvE+/FvDXnbRleuL3H3iZ8p8FC3Na6uYJ6/Q0b5cqsDnaARFpO7uzpIThwm9nbX
a1FniTyagNQ1uKLTeZv8Ap/lLNI0EtVZTWJk8Y3a2KKtYlKLzhOJln1obBpd04Zv
qJfm1cW2y1Y/rCJGG5/gKx3Pt4vtqZR3yDy+vL7ng0EZlmHmcecsjttZZtRNgyv1
oO79j9Ww94UQ8n6B+sxXAmbysVWpW6HDukMrn7rwTCezwJULNnX9E+0Gh9Fpg6tY
hyrElHixKCGDvzIvGfS84QQRH3J7vAeQE2LN9v0WpkGvISLZCGbq9ePddau9GLPF
QnT6XOnTOKkTnigNP9empRgtVryeaj8/5hBfeio95W6QNYmHUisRbeCfOrqgJsne
hoTUMrGERVEoY2KK7L0mCsZ0cnUjoN8bELO4WOYz922D88OcCn4ARAdWBxPvLB3w
B0uebitQNRUAXh/9/MWq36xRLS7gZmCjUgnUu1mWz7vSZegBJsEKcRtRlCo4fGeu
uVETyVZMvUZNeLM1NaSQKYx9Ue8roYc/PSLTpK+njqWsReBQnH/vDdrZMndwhfld
I9BCe0P3QXSt0usErDt1P5zNZKKrsYwcjQiUxuz4LwfnGRbf/jwZVEweNWFjSme6
jaX1PLJ9IQuTJRPQGLhvK/0Kj0MxOQLvtkQnvX5T/O/scwyv2yckQ4m8mH72omoI
z1vbxtiVib6SEdt93xhuKh3vHRdi/NX+jTPjaUDmpX/ArmtmItyyRVzx3QcPkwsh
mKn3rnls0Zt/KTEJs1Y3YFeHisbSAp1l5MC2NsI6MbEgVpFnrnV6lomanWvCua7y
ez1mYqC4I3oGp5GdQRTUa7zJ3QJz5l2BdIhj5wvtwEuxwNiCPRUMcEnjxPUNGg/Q
HvFlx1ILz4GPBmxwr1rJwAo3NfRHOxUg7/fR4XDS0PCC6XJq0G5kBK1FYkgtW8DT
OfJjONkPgy4gviBSs1ur/u3qsFmU2nFIilhR3GqunNilq4LaP+DHzVUuPv4C3Ds4
yll+7PmLuo+3NL+tar9a5ZPAjHRSKvG+HdXisFAYLIoMx9EiGlHyhsHkxLcGNCkc
J2wsGu6ri1REVmWKX8IJtrB5rDTjgb94DOVUJQq2FRcQ4zOfQrSM5HGRhWK4UqcB
VoyMFW2knJFcXxIRjvPukXMWtXVvOuuYqSDchnfG4HyCeAQhZEpU30xH3Y76Ol/R
Bkt1uJkN04pf8Xa2Hoeth9RwAAwjbTmdXf9ddEz6gozmRtsOUqZKrRwjWkYI4U0V
rNMJB9r+QDFZL4ZoAR/M5Akk/sqEsXgixzaj2O9yhmDkyBd1jq9ti7A0tFJ6Zbh0
14bCrpN/XCqkFVhoRtc1tWJ6SioKiB3kEVADTr5922t2G1W79TwKln3BSwmuSQQS
fUI60B3LzFCZsF4zADpDNoe84uQ7pUnuxhPAB+aSIWTE7ECxugo4ImUn4054Pb4K
B4PhOay8k5Mk/FHGRWb83/vmAQB1x99hkDEFYJR2bvbAM0dBhdXsf5zOmvVEToKN
mowuWvATacGvsnw9RrneofV/mQ2Ck/TcFIhspt/voUjXjyl7/fs1VRMlZdHPqA/w
ro/5L80FI6+XwQYUm27Ser7+dWZWYWDosnNm1m9naigUWuwNqQN+vSceF2Mhcr1I
K6p3hGUyr4KbI+8Lf0lbdxC4OpILvzCEQQlNs+JxM3CvDRC6A8Z6aC9lS9hAQKAW
vItL6F/IwvewCq19XTRGxy+L0X5RFK+SgVBbzgzwuMEEatLn9+hZmtZsa2PKhMcG
QICi0UeOTTpurYialaSLg4Cm8yQLxnMlQM2+QVZrC7GAKLebo/WgW6GgBcX/VhgC
e8zcc9h8UUjoYK3UfSMAq0KNA4r3goU5vaIfcWqUBl5bfXyfad7EEfrXCLmx7jGJ
+tFV5iFIUQcghDX3ID9awKKmCHjNnoUAV2zvLJtyL/xOZCz7Ef37yc0eyozDILgB
QW0KauK5ouRE2Ku9er7K90mwVJzF3kdfA3ZavNFa6gKtGgKvEdQf1znWBij0SQ0/
//7ennN586qHCDNLGhLjPWTc7AncnBnWCExgTP1HqqVzWQ4RiuBSwsfXqqCYxmn1
wzbcFmAYaF0UQCB93kf9+SqU9FGaX/gvj+n8o7wgvI4LdB9py8ySziWXgeMpBZfQ
5bWXHrsYQsoyfBk6bE5no6HutoMzcX9vwun1k2tOzyXSj2t54v68V402MBJ1lL9k
A3kteeEqttX4rlkgsDRgN2ORt7w28nBwpHEJHW8xsIh7Rwwm+SodhHn3oBMGANkm
QoQJ0xssXutEvnXmlzMVVJOvGahZ5xqzIWgC9Xwt0MhgbpiWop1V/U2Z4jq0xLV1
R+SU+VUkFIS1+nxA+oaZoGsA/p+ukVTyq0CUOR7xDphs0botGuZzpSdTBYPhbESc
rABI5FqeKg43sUf5atizbal4Y9W2Ct2CRcNNbp7PJgtNsSpzs0vhIvuVAmVymbuO
RANkLui0MA+wW3wQOb3muxvaaJ9NfN3tH87PmSzWBS5hs5tD+FAfEIkvjLG0Bg2Z
hQa7YgdCqhf3zyeChXUMHr+CJ/+ANeKT4SJhjtjgwFIMOz/4ZvEnZx7yN+AIJNj2
KPmm/D1iMpzZctjiTBZm8ZM1MWOU9cSPcyYHf5xrvHv/x+G6mANZQj9PTFNY0D7R
pVNyv1gSwbDHAoeaM8gNXtTH9LXVK7deGNrM0TKQXK9pohmBttujQlB0AtbgQMkB
oG6Ntl9hyano2vos5/33DY3glATKkTX7+faf0xs0WN37igjlO136JUMVrY4qFLkt
2zr4H47zZ6YpGbT/CjuixjjAvgEF5bU1WqduaJaM586TlToDCFxJK69BeDEhdRch
QQ6/NKGDi+dGaqZeVQPMxAj1lXd/63mmDyXG9Pt73tzZ2b+QqK9GkAhh5MFmPGo+
5/P0AyE0la50hTETYDyjA76lpnXPN93gW8bHknaIdoKmbot1AQujsF1ibTvd2+eN
OxLkJ+1hcj6NPWVRqAhJucZYcb35MlpWNuD6nqp/DMf1E/Qxvt6cWQP90B4iU4dI
fwpjpfXa9fNrWPS0noTu1nPJAlwSbrhZpwG0dYBUS61XO0oLp3L7ZiYQoiHvqryG
xidpLQXa8VJGtK0VmvyboLf2V36o6su17JB8m9MpbDyJAIYkfjDNSgS+Yy/H7Vei
L+VVj+c4z5gccKhcJci8rDLVITDoLyg0BUd659LLxl4AG76IHduGsFTJCnu6SQYQ
xUYDcKFvC013QI71cXkxRrhdPdFGckcUaWgYLPUj6VaznWVww32+lz2snIrfDAg8
oiImyZ8Y0jaVYQnJoycFQRR+KDq5CZZADc8JUuuziJb1eljml52SlTO59zkTybuu
FQOI8h8k/UEf93Py5/mZySQzOIUFCSG7NWlpZl8uuJmJaW6U5zM7fNrZ1yETJzQ5
dvyn/WYxFIO9uTY7azdhipBuhixWdLoIAiZUm5qyqsx7io17PChRdrCy2wt969AQ
mg4XZG2njbjLOEPZ1Zx6VEF+wW1Mi8FnPHqHA9TCTp719iJsZoNXh7mDkKVLmbK6
mSTJsMOK//YNy123BAHR1Udg8ItEDChr9Vtc9RfKuEbzp1DsXf16GYwZRKv7040S
nxg1IYwKMhoAeK5tAIDDKsCN6qNrxTHeSDo7ob7keMvJBGP0o0e9w1yEaGCewUQN
m26GBbJeLDczsKaP3Y1mqTun05XKujuIhdcWHc52gwbjeSxomaO4x22PhEjjW5rX
v0qef/azNuP7X2gs07LpLn6SdrVHJ4+hfuthVoxjsKdnszfZlQ41/YMtUEdsiWSF
KDFjN7Ap6f3hymefDV58DNW15YW1eFYWbHfWzB/g0+B3KkXC0PM1qYdUjO8WAK8b
Jx5hqq0FgE7xHEcEUv1noW5clK+LKen6f9P9Vi/B5gkKJqI1emL1VLEmpw9eSf2i
9MGrSiCZIqtIPkSrmjRYORnNnROV3bcIlJWoVJYst+BSEv5x0y2fda+4RHOLNwb7
T57+PDh3of9mlY+DOKbnrSMDhz7dD1xAc+ObqOa11br2uXYVsqypqD2AeqLzIncT
2V91Dm9x0Iy3AHD5yMaTSKOvqOZlxil1AJdlbnKiG+qBIiVLuZlOFsf/ro6ZGunc
7qrJ9SMloA+MrhmG66KyDVoBPA1VUT0jLq8Sd1Zxoc63vK/inChoQ79lsrzIBkwD
9E95sw+OafI+O8xRrI0VKCjrMlblPLhWjWYo+OQhu/Cf5TXDSNzL9FCu+16Eges6
ZDAkzRjNjYMdeCj6hSirygVfJvJ9N9jqV4KGDBUPrrO1LR5yGrVAbjuF7j4TRxLF
4fCLalVbdDyJD08IgqGKW9koA1tWrjLVj8tiXXeqPtW8/74kHgsdv5etwF0k9y6W
eleq7EjwCK5mNVjSOBWncbrDvgZBZNnLvi+M28mFGB+t2fsdgjFIUO4raT1I3gPW
D10/kVvUx3yDBt/FHhW197xT7c/yyOW+EDFX5CyJjn2CYKkMv/H0/RgHTCqEA1/s
KvNPL2K1bwkqgVI62YLCywdEOmYZjuQf8y6uGZyl2NcHRXSdg42hD5KZighfL0yj
uI0InVrCE8ULZve914QcVKMs3tyT1lmBgz8zzOyEg7JDTx9DSAr1/CqGUNULrzB9
F/n+qvnJNMLmBIts+YCrEFjk09Vkt0QmCWBKxXKnLnvBMAou7JZYHWNjrD82fObP
ieYtK5n990KZ7W2Xtl/1KJhRtdidpU4vzRENM+WIH2W9+RfN+jjYEGaTnF5selEv
E8UnjYvAQVqrRXpROMFBgM4eFBFgrahtxLMFryO/rI+s+CmHXjZQ4/8R+Ro9c4ay
oysXfA2tWedfaRePDpwOfUqIhZb8iRGXxay0Xw2dOscMiOgspyT2o8ep+SNV6bly
Tb3UW+cKUTmmqfmlk5T8LHEGVN3ZIOUcbCsaWMaP0mpXZZMZlfnQ/FhtnsrdrcgT
0iqhTsp9efWkfDQQXjYHl/iUHsW3orxdKb5YjheZ8gQSu5xycHwkWDhtpHtBuVFE
6KY0bGsFXJwb8cafYHifC4Xj4sxfh/dGkqQ/IlOeiqlrOwojmjpLdrtbxCA1hmAw
JfEy9Hz4NgbGrNjxo6rcERHYQ7d241eA7lMsNnd9HwnamZzzG2ZZpRtlGamysSnT
p/Qr5HLEAJRhNdAkGy12R/AXZsTmG8X0Ge4v3XjTP/eZhcm1kxTVOTUgFvFXlkF3
AWSaRbWh8vVjKKEHmxXdOoEruuNgg8g6iBb9dSsnbGqJdXvhIRcg7f//9X26ipux
c7hhwdfGnDlKxB+rVh5Avstmmi8JzUmYnCp/nUfX8Pzq7jzGOGSS/4qAF0xAgPsQ
pUH1JLK7YGSH6h0inEz+pLZimjagrboP519ligIczFRdzFzWC9shbS3jXPgzaRVk
wZRO3w5uKXGFm8TZXhhsZa/x4XfC1zwNOTRoEBrl1ulOP14YrT1wZz2znL1CF0Ef
0+YqF0u/Uo5AkyYHzsreI4mh6g6TDKfRUhGFbIwtdmtqfOu46uh2rB5agso0PBNH
rwWod9x/Xqhmt32uvIDrTJUrsXJUyoP9RTS4oXQIoZRXGPniH7Ux2X8zKDVgseqW
UEraHEz0MQvnfegY2049CftZ3q9YmIWQa8RXtR2KpmnDy4474Kk4Kp4qWGdZl8qL
WX+hvotZk2LUXs++xBJFHNLl3v24LQR+ckjafxBjUU3BA/pi+KDr9ByvnrgD8CtF
FaM8FO9awcEG8W/7p1WdS+j0rfHlwLMC81tfExGtIMZAqPX88KUKiwIJfSiahfOj
YwI7UdWjlLOuXPS0Xpt5qHvu9V1sVQ50Uvicw7Z2QdPcw7yfOap+3oySe1ZeqxrV
uYxjf+LVwJMhzRsKSNQK/Z80auYqEm8MrOYNsXXjWXXwfxcHFQntz/kCFgNarR/1
FH+VVT0HY4SGzPF6lMzgiCbvEinlZq7oFbDv7bRu1d8mqg8uwYyRmr4UTN9Y0bmV
KbQrnBtkOoKEek9L+vU2dKTFu9Y15RUH4CSSGL7aXJHfQiH1eUZfHCQmrk3dNs8E
pJqAGgfRNcPdp5gtJTvn3H54X+ac5L77EKuRkL6cjku4mRlCCmC7o8EJMRJ6OYJX
CV2Z0IBL4gVkxBIpjUyAYxREDmlu4U30InMEAgpD61VqzhOQYfmQd5lYufDEHlb5
0J94a+E32dsvBDnQxYSOeJ7NdAKaFUq5b5XmDgdc/HMw5FqX4yVwotyDsM7auZHs
xPuVG5WSGi2pvtOwQwt0XM7wBKcH4dLsSnVAAIU54+1OwEToGl347YuUGGbHquN5
Frl1/j2NDkxs0e+fDG0tzzPjnQ8MeOjdzGH+foQrR4r77xr7e2Fq22a3wDrUWIkN
R83otO/YrAw5okaAZfG4ZqUxZFw4W+zlB+CbCBloYrh/J6QuZWhdcFF6pPUqlFGt
XkHDIbvN1wwd3paR1W45KcJvxYO7PqfoWVbAsEIYlX7M5C47LwO+bXVWpIUb+APl
QCMJa1n96tQP4EQeavRlRI7lmQJUaOmx6xxvMdlomdQAoFMmQdDgxvdB3t2GHSbB
48nQI+xxsYE0tFgiQ1uC0/8LwR/AX4njrquBb/UZGnjP+ecTiczZjj/QtWQrkQUn
99STQmzKZtrFLeztPEgTUy2lZcaZiIcIGs0YhDkGNcSgA2186PnTxRPLKdvNoIB/
yFdfBqYr1LxFH3qmNay4Qwl4Tb/NjnV6AxXkPKKKvXLtGvGJF2qbVROylUhnpPqv
IBW4DbCN8GNmi5syNIlzM/UyCVECtAP4wDkqimt02Pwf2XXBBDIe7gZjHZlm+eEX
tw4xL5rH88UQvvrgUncxgMurG9LUI6uqqjXuLtL6MIFUZoShzPc96vEaPhZb950C
poMZmifyil0Y/dFUgdSId2/Q1of6LsRQ94bjXQsSfmBNUypx+SRAjFyB2jPsOjfB
Auia4s4BfPyquRME45hs5B3FMptEidyfrOHHRyC36N+JwzLtBCdNqnQu0rox8zep
uYkOZEVG6FwAC8u2Figeo8CqJ9VBCt+DBZQUeyIxl3GtlV2N1cajccq02mEi2yjw
OIwXRrwlPrTiX9/JOGiwJ38gkLEUGyTum6MYT6lJYxfs7UITmFyEXgBLGY51zAm3
+XkgQCQqT0eaRH0ILbN6KDsJbbln60uRgNN2vydzwNMdvExZ9LqsiAFa4/1I/nx6
2KRL1WsJOMlAPMiij7TYIdT7LoUb1DikXwDFkHZhBd9piOituOenYSv2TBy+wvqR
U2H6FvzH99Vw0w0/VbUhDUKoPu/X9u+34l3chtS1s1geToh13HsDeaAOmZMoG4E3
FVvKj5OY7x4sHzmoZvZrjMNo6q1c1WaJG7ZoQu6iDgohR/0EjzAOaVoLj2vKE5gB
K3muLEksvJfzHJ9rzUkHKSebsRMzEEIGOGvohlQkiwda78VXApaxCZOfNH/FhLgG
RlDQ6v9UsuuCxfB/tPUK8nDoNXEtZQqfcDvNdrYFQnEP/bYI/AEEtQ1HSD39tVPT
b4vEX8Qm0hq7Ptvf+LFxoWWq/lyPhgO4Km22GTPcc7/Aat1UqdkjwPgZChX+oNsq
+uH1oAGC1xfuq0Kyiz9HLVHlgLVeJMxofg43Qn/3PBRQlT9PDaDiQW5JPgAfGUuI
BqOFQJIyVcxaIt5/Q9eOxUll6irA2aGRlkra86+ADmuzZzKGpNWGSXee3r3yjW5l
HtTF6sZFC4G+sZGHFRWZhLm1u1TALUHACh50CRVyT6wMZ5g4gTVWXWZrT1RDCmK5
ZR16Xu41HRzCW83YMfMlD2xLSY/zQS9ooj7DrOsH8rxzd6XVV5uLktsHUE+F8Fa3
CrLQOe6C3/kCJPHcEq6uVPPpHqt+cH3FmLg7/YMkHVKB8YYJImUj4Bsw+s20ybEV
eIn1qAy8xZu1956gF4yVZbP+lPfHUMMNkSzYig4HtEIp0HwSC/Egi8v4DYJtqgKz
gU4ZAPhObaItvpoLV+ISUv5o9h9pG07/m9PvcKTfPyBTneqAUmzt3irNSz8J0cV+
hwunvh7114Sy9tQGu+cM+vB/dSKk9plEfhT/sBu84+M/qy3Cxl/vnFJ6zSc3SREO
ivrAOemEXWsFcDCvtlo+l6SQ9hshQnJTeNzKIl69lcllMxxsAYIB4ih1wUwju4g+
5/L3J8TiPwrHru6nuTdtXK8+Qyyeot57Z5j6Jv5a+pQiPOC1aYaLryVjk6fvuKHy
HY0eM3vzR0SELWhd/8gRl6Uu3iKe8y+pSmXtwemSSNMaUKVQlv4i88zFLmpj3zSw
ns04A4i5V8WJMtIG4AwOwBbMtsS/vddPfVCJUAnW0NVUMyfI5fU6sqh9W4a4XvHv
XNHanViX4gbS+Ikq/VjpSMJC3pvlkdCn/icoTuS+NsR3uKKG2hme0L5vlcfkXEY9
MQX42AFS4uHc29u+60n7Ot/KKPzanEWc6F5pTDfPA7UFbnqDtBjVEZ67gxMeFj4x
8nyxYCuut6zFQ29X0TIDuqGW85zd6JpoWQUZRAv4UAPzuqSlvK4zldkExzlSVbDe
O0SRFTEUhjz4Mj0RaPB61iONUOPQKOQWqXCjBaM1VWQptY5kFJFPgj6J1vZQu/JF
iZl/nR5z0DKRVeSQpaWc/sAIm4k/qb0mInzefe+mGKe3DmPq487GigMjso8MOksw
NPdtQ0kqcH+brmRYb2CTF6qbE8r0VlmgwUELgJ8R2iD6WTI4FL5Mu/lU7tokg9dJ
OGVL4z+QEHJIzUNNM5O0BwmMofpLh/2R9jAnUs578+W1qNnLk8cV0DEtTDxell//
uULjHEnAfSe+9f8Fq2nGjA3tk855w8iRrUUVWa60pIrAjU5vOiEbuqXK3h/k2tMC
ua27NiLToHpchxVoKGrr++gFZ3x5u3SCF3BcGbTu6AK3upsvU1BGxg3BNeQ+Zdzv
Az3iXvtRrrywRltcctYGumogy6Q0RAP/7G281SIvL9bKWvr3qM3X30ZSS6Kfilhp
O8X/TK1sYTFoHardTqg30MptWQoTxBJP0EiM0z1JvVy0PFXQdK8nlqTFbuwFnFrQ
fcwG1jCdPTe0yJbkQFbWnHyv5djUho2fh8TxgmCVhiUuNuM5syh9Tr+RnBbK9fGM
8INrcQaHiXsA/vsdBhbnH0JgzEOTxkyhAjy+7a3u6khUmlziAPF/VpXvaTh7ETn6
XhRazERRyzBu6RUoyxDuq+ZXvpdxs6X67JJnqwLVuToceEZAuZG7TgsiihMVyOeG
M+CVL/9dWy4zBxOKXIfQwH/wh0LpDEmkm+PA955MV9wES0Y5C5dERf701BwwMJGW
mgxqVJssHrKJmc/TRWo3MMh0jHsseqhy5bd0Ef+N9Z3Td3tExvMm/nMIreBGQOJ2
Kt7dgzJQ4skIofTNrgjMlE7WKTXaswcqDh6f+1LA8hL6NM9zbLQeetWlj80BTKbB
d737H9dxCSb9jSnc3+bkEobVVuNqqWs9Eing1oudsKaP7+51CZHOL76NJIA0yOl4
FgqfrAmsVNBQxfev7+WT9raiORmiMyV5LKUA74z/9f4w52uV2RQdw20NlT61Y65Z
Tn2CmYgFPre+a8yHTKkSgWANJxBmy+eWXDfWeZIFcYC0iX0sMyPu+gpLYNkh+V0V
LfEg7gjBONzdpTJN/Mvve1Z4q8VAIh/Epc5v8YHAE7VrtW3TIs11XeNqtCY0mFGb
/I08S2NJz4JoFdVrk0YPYqoZhuMbfK78aBnxIPOgJJ6vz34HTMQHGHII3zYfI40R
X1aqDx7/t8A2W1BAds7zQQoPer7fOXYOBI7yt2rjtTRVQIJe9fdeKOIh+ATWlAJx
K8xeVkz+f9WWPEBH1U5BxixDegLUpgz28rX5qUeCqIMR3tz2rEO2hBLlFAZYGaGO
gaIuCJQSeHPhfToafksx85VylCZhmscmGX+I9khXuI6TispZT50/l/xjaosRKD+T
Wqna0mATpdTVqhjzioiuCTaaqhsTWdUhE0DG1JOp6aqYW1yMskCZZvq3vEuK6NnZ
O/DWV+45XS5p0w9ZLWDOAbaz50ChfpW8VinspjIG9Qkdn98m+cBt1AEcUOOnzDbk
aMBbLEk8/Cam1jcg1TWGxgDFNd2Y2Ve6GW9C/KF5fziPQL7X2azyo2E7Mz+B3PSW
TTecAQuIY+6lwKezNozwXLqw0x66ngjmnO2ML38oF67UNr1earJzzSMoxNoh648a
6Tz3vkPr36d9Eg+QCRv0uRoWxv7MFw6Hxz+InAMm0RzIZR/YS5L4NlRWVeacS8kO
0PdZ9fZr0+OT+rH1MLxppHXRLFuf2ZlpU5zufZjZMyZV2cozTwBWi7Zea3rrPKTk
HN47asvEGiadm1lQE0TDZaQuI6wbNcTav0/JElXAJFS7rPxXfcX24DBkwl+hBVyi
z883IURI6MUeZhak9kGa3abZefcb2u8WosBD4Dye4gZ4IyCkUXseGOhi8EQYTpNl
cuB34AWsS0NWfG8tfNRZsWOlKIIjnXJrS8ArGJvQTlC52/Hz/Lxvs/kuC7+M2Gwi
6AJwDY8GW+HinztEs1QRLObEiNHEBpopKE6fBMF6eTltw88gTCKpYx3ZQyZQEgre
7Lsq+ouYgvH/dXJnu9fAik9fTHVOGSV3+awS054y9qlxG6+JMc7A9O+679k2qWcx
rDvpv9/j2qmO7kMmrkRt6u5lIiMmf0eYP+vRKNWuO0VWx3L3gDcM7yW3Sdlmu33o
411mSUkQYup4OSGxA3gmks6FtscJqHnwpqeMf5vpisNITf+zBXalkekz+IEVUiTl
R86MKB0mz7lE2EZiRZOswn8LlE1l0wwRMBlpRZhY6b9m0BgZg2Z5T88mNj2bq+HY
CniDsFbu+oI33gfPfloyw6uV1xHQMfI47tl/7yoWM+NfgY61/QZJBttDevtEIjwj
O22nj27fF4v8EEsuXoesQbSamdThkwW6HuCe/hwZy4/1eHtBu4FW+twBVBLrxkh4
EEXIKvt4slLXYxDj4ZUh6AacMs094r718Vgo0ew6YimmQM/AW5yqjHRH6mTmBZ3e
W+EE1B3hTPlwDZMHePYZyRj/5XGc0GblkReiKtRFt6L5So07DAwzDywUQY/YQ4Gx
1TAjiceKefBAhnyxuKg6mz+RF27AGRMo5Ri3bBw3WcKO10iSd0rxelkPsxp8LAgs
ZZdDndDvc7pqpZDlk+17OM2ssdjsObajkqrSCbAfc1Hs7/limghT8mldapU5O2hA
s9PyXAsSb0+Njr8gM7E0xgJQzRl6k+95PMmH0kcJG7nJZ0NmzsQnrF8U/GVJUOYU
k6n9s8EdCQB3rULb2MeUjg6UgzuiOP1GMHrPPbhlAVfwfT1AUEP4jjIzh1PtA8YO
V4iML7qtULK26qTufi+5xvLaBGyeVTZW4bLXBCebMq8rMLrljD0zLWQxsLQNES/t
pc0XmVfpEeMHVx1BR1SMbYAi4QTrrJmBloq3+cpk96dsFR++N1osO820MoKqhIvG
mIPxsd0G7kJ/nYI4Esx8+Y5ZiMaxpH9YIRBoRnAD/qTgnZ3nJGmJWyg6+euNk78z
reI/QiKUO0qP52EOa+sQEleTt74TfdE8GDQVgIjqR+8CAXCkX+EYaasVpyUiHXBe
z26fr7YiqQeYdFuLZwcFziPqWUC4JmKl1tsC9q0duCDuCOIIVkaKbpypSvW5+ONJ
r/k+yiLmHbOy3rMMcvQeJY4rzTGgpYL64seqdrIQHLO4kWOvhv6jmKDai4+QYiCK
quc4wvIYViZ8Ntui2vvLPNNcfQoAZ9ey20DZuxjVqAKLkrVgxKYktZidZiZykukP
/5SOJegvLC6xZVviCrByZ/bq28qj802gWfTcCSR3hU+fRs3WBiwo7LIdMueau237
fWFqHzjsuxyjBcwiXUsHoBpRCC980MLAhivFaXkwbaxs7sqfEW7Zw4q2N/wpy9Sm
fOnTqhkyMnl1AX6X8IuHcBVNM7ZMWnHxDjC4Ay2UtXjA9FSVEZ25+yrerx8/5UJM
N2BAjS15XTmzWiREhJf9MjqfQ2cEXUSO7qNDnksMm85yLWGGlYx1tVL0M2gciKt+
bRn6YTeCS3e6kDtt7grnyQY4aEHCPT4iMkUJXJ83YH+WoXCcZ6rY1KI/1Sx3icn7
v++Yx478hM4XmBFcOYBkK0er8iRwBtal8zywlqgw1fmZ1p6pPOYSDIM6CzSuY/E5
kqDOK3eKR9Vur0GUbeyqPQuTeBPpSV98XOe/maW805BL8Heue7DSi0qO/u3Lcs5G
CAyFQGhw7sMpXeDLSl+zNCJ9T2rbGdsI4mjJa4/lJ55mi/uTchiPSZGfSazLzJLr
UsyLTK53bvp5StyoouJQuq+C1kmIaf1E+NaiD6/wdXVkGe/KH9+ee7yB/NcImeGY
mwNkQrnazFOld3xPkyLsN6s7MxOViD4vqNGCrg+CgVNpDx+KYVxGZWSpq4eo9ZPf
fxgA/kLVDKq9xvZ2h1QemiJLoVK+y3uZhvBq9JXDyXkflqUvCkmJOcdBSZGfOs5i
iHgo2qZsI1Vr5YNPbNnvBLAc8A5HKuOEVFn7d3WhlWUNwp5QpamUok9mq3KyTx49
E+EWlVewSK2kn7550ZdwvuCPUCXNNzWeId3S9V2cj0GLYJBOcuw3fxnon/FUXvF7
X4Ow7DIhvPcgKKEUZntanBE4CYI0BoH0S+gL9ssuYkuhJkG03/ge5AMX2u+3EigP
h0n42pdmbdqqmbFMTyq58wFSRiCel8QQfGab1chDQCEafmBk46TRrCMSCnipjrmK
i+SNtenykzIaD5FB9QMmCuumd8OaqjGy/dEix1412DjZsAIAJ/ibjCGKgrIqKnQU
JZ4vIvKdhmrcipF7lZZMuLV+dhbt5bZHqJC+K+avBRGlXB4IKyyDoBEHEEf8fXyr
VBRF2db9QV7qkm6oyip0Mh579YZX2eAs/IYKJVhLki3FAOXd3k6WcA93KVjpd9yD
mz/epo0TWojb7xGZN186P/8fb/w21MR8hE5rLqp8TviIZnhH6ImJHRGERtNAa82k
gTnuGv4FwUWqpLepZgya8DNMp3ir1r/zHPLBZ8GidNzG2NxYnh77oQqQQKZVY/M+
t7tbO2DUUxphiCc5lbzcUtL2SXm4J1yDP5gTSlNluoJnDuE6hzUmj6cut0OyWSIJ
qy8Zz6IMUSk1bxsvRrN2AhC0iNXnnlK9gUR3j31fo9DX4rZHzPRkUyNPclhYA6JV
LuTnSX+vS+D20I6I3GSDQo/gnUDHWWEsQjmGOScOHADuhPWNbzSmYok4zW9fAM1i
nIfBjDNRPG41pfZzHS85hiueZoxrjjMOxET2YRJRd61mKLqk6Mtn2zFRW9RVaKDf
7BD5+G92dUucYs9QHzarlRqLwpRSyJXNE9ZEAee6S2GndHibl1hc62zzMnWd4w5T
wxo/IgzM3RKYx/k9Bgk3UrfQ8T6q5eRqsmotITAQ/U6xfte8BhEo2xc7ii5hs1P1
7v/NstXrORrizR3Q+Hiq+IdqVDnvvAKJMgJlm25xPrYp2Z7J6G+ywJhipk55vPDl
Beebjqccaa0NPME5d2D/CO7VVf6pkYUb7CU+bUSP4B1cDqimX1+jxCR06gcEexHJ
k/T77omGDGt37XCLHfSbMrpZ1dRkxEreGUBSIzpB4RtLMsfpPTBQbi+oUgP1/m9B
PL1VG2U7lcR3Ic8meTMiE44WNqxI+ySQKwTwo+tq0UbVFYLEV6dPqFkc/vM5XTb+
xZxoZ+HrJisDifYOIpsOZNBMSZODKvNmNlMR0+lSuk1AqIOHsqOMzp7dxAx0oJzW
n3HTc9MOsh8npGBFhSBsfiKtlqcIUocRCmWoT8/Zc7l9DG8RBqdylXvFytINz21T
hn3FfBlwOxZfVagLeVs66FWvGB4XhkKJMVc7hRg4CuBwtcCERjWGuDIk+HC9itMj
+pZVSr5VnJIQVn/NJD9kdilv9YIAYh8frkys/Uw0I4BYekbUeo8tXktQAXn/Xytq
8/+8De0rEYsa/pFhekav9Icc+CQrQKCV/3PDJaaz3fJgS7bukSt3KDxz8X54fPvh
iwSQlfjR2G5JHHvFRIfSQRTjmewefislv6iS9fn0wJdTwqMCszcXeZ76IcPh/As2
a1CLnfykAJ4MU+L+vGoo8pB1+SQpCTjF9i/lYu1gCdSHXcEBnhblktVJkm1xCXi2
p+jtm7xjf4jP66M4dtsU13S7msT4c7/fnTrI+B/jhWMs0GXC45Xd3FaDdnO9bXvJ
/kgriORVhb4NDhs4TSPAqrshoSLITGC/4JSu6M9D57uIp4c97dL4p3k6fEY1tHju
t0HOAgE6F9KA429sEqPsOELCEwndmsqyYXOJW02jALW/7Ey8gonYMLgJi9q0jgCF
1DlMzRowkJvlRC5LpnmzJ/RjfaPNq52ndudi367bhblnBZe/+XWUGFM5fHMWeYxY
DHH0hJgi/5DukTt7bHVOnFgoKK6kYnRtQVrsYWqXZUVWXUoCBW5BsLerzOKcS0lH
gKVoqDWXBDuCnJPvsPne4zxg8IZSpafX9o9r0WOiXtNm4nuAymp0JMFoDOqf1fzQ
0/SYKNbt8/PadSABS1xSJi4pBuC2o2RHTnN0gLAOFJ7pbvRzi8vuwNdjncnOMGXx
cNy7ZaLgopqjPgUvroKDjpaGok23hjAHgDteByrcHixsUIRLBpYZaKpVxsJrCKmh
rjpKZCs8peIPxZkuok+rx/5+ZiXsZ5sPetC21I4vNR4f3KLFCKrsR0aFDXrpYZ4F
WKz37TD39UokpPg+VkATPdu0+THCF39L6mPS3cBgACHgXCrfjEfD9f/V9qzKSua+
p516ucG/h1c92K5+c9tONI0SJWpjy+JhJyp867xwkria4QF/238UX0XVDFz053QY
N6mlGMSX2Ad6Y1k3ZXrFIDHpH6ZyrtseJXpfE1t4GLE8jP4vmxAhkOLe8oTrw96F
vvfQuCZJhLdJ/0Z0yjUB5Q8UrAPgdvtSHz8foRLGFulvQuGgBAqzYyWh7vAoq7qI
C0krWAO3hwsMxsiw61laQwduBwrgfs/m2Gk9oaJGpo8hLB8hooIyz72th969xPBw
Hbv/0nmP5eS7WIiUwJhSwy58bdtbDwyv2hnvjYOREW0f1JHZVBPfbNPrnA764SRZ
5YXQro1FHZo1Lohs8uaMqPVEbRPs5ZNasyWsq4TPdRQIWvLH4H1jEkE2qns4KM8O
4QOV2c9w4pTj6L8qCCZo6MCmbhTm/HbgdM9MOlCfvBspd4E79DOPN9XEsZq3vUar
2FZFCCqBq34kFbWNFYS6KI79bvYvJJP+ZyOn7EpCZjHWBl532VBD2kE18qQzlg1+
drYCG05cAVrFhB/TKW3Se1wf3JXGID1YrwChfxluwDLhwDW8+KU3V30fdjxfcicm
enbc4l2HpELjN8+P6oNTOOnAwtPWM3GGEVNHP7X9RYUJvZAr5eok8oBWJjc1KN31
e5EBQ1/EMFba7d6WOfT2h4fPnO0S79Cmal2xoLSnokpJMLq0Fhzir7lDYGqPXGE6
aO0neoAMnI9fPi2QuZ4J7dItrOySg2GvB8NYNEyrdeKRiKdK/V5HT8VjYym6Dvdn
sNAaw2oXbuIO6vLnxct6YZuK1m3fLGL8SccNFU5aaMWAy4dg6nEEMF8YGMPGXk00
tEGw2dzAOhZsvtkDcmgGuC90vysLEtiN1ji7vZgDwUeGrFgO1qg9ofXVdX+DZCAx
NCHdBfRjWzY/PQdBmxjbrzcyn6hMcicnnRhlgAPzogKdjduFvGTV3MIVHPKsf1ah
ktEuQnl66qL5yVgqZPKWbzGE/cGstiA7kHeQhYPDYSZ3d+CkJrWFLAmeKn8CIqWS
umtn3I1JTt4BZopVu+Uayo6/zPJcP4xYX205v+pUBYzyOTxYc6bCZSsC6LtsVnt0
KwVDL1wmVhbMIt03gpSYoDsULU2QEp+k+s9tM6KFYTDW2LdjmDEnj8ZkNYI6fCY0
iFrsUcpXB8+Zmxiinz0Udqf02BaTsJmPZR7BpqTV4lQfxg7GqAXe6yYgpCbH0XqI
QjpXsUqFLdx8q3iBgWrSoBuwMYEZr2D634LryShi/jfVWzsaPtjm7MceDEBfSLfv
Iiph/U5zRdm4o9OekiautDK8Gs9b0GTScM35yeuUQwTOoGRuIt11Vkkpdcx7bGcg
d1D9DhQzmsPyQUfTEnrB5WH7otmCRDHRO1soMqhr97evQCOPj7T/ODJoaAJ4PiDi
OGQHK35+vF0IFXUujpT4wl5EwGXPS2+cqBgNrhJXGU+O17Ov74B7JNo3MEy1s8xu
7B6arwX9ga5Qcd84AIgA5uYANTyXr/iqMvJQ6zDiFYUjyv/Htegx5U3PeYGQrr+P
iKCQTTbEYHnDVPtc7g5tCidgF8Rjj6eRrGvZu/03GOSNxvmT4QGayA6EzCwbPUDx
jN8Z3OJmP/lLbPSq2J/zAmiHxJmBOFnoR+R0tCDYaXV9ZSobBT4tRvOK9bjJc8jE
G93DP9uL0emcCNh/IbELzKohgUT5K1GhWnMV4z97hNgRXfcZGERws7Wlz1BNebPB
fY7EYFTJyutkI9p8TLfDxPTjlqra1C9JXXTtAO+HhNrSKG6jNk8vyU0GpIGgMRn5
NoPSSURgjAW6DrVxmns0NmQT+gLVsEDEa01nEsGN0VoaPxk82302p+yns6XWYqxK
8MZDicDgEKXjlRmXzk6eK7EfKxZ5vJiE7dQB1Udrop/Wk9RsvW1p9MCZG3l/Ul39
+qS+sq2ZU+OBJcW9wh/mxDBAfy355WPCeNgOhYbAxaa+cvLNQGoWhxukuLcbz85H
7y8bIoCp7JmlZsH3HsIvabLzNGPZxg1xLmhhNrO9gPgwyQdKLEpfa9yw/K0pXiUX
BZ/7whsMq2xUF1g5hMohgOjXV4nrRqBZSzlIWaxq84oaEp2p0CACsKNHVbZFX/jZ
xSIgJmrhCFDLDSj6mmxS0kxpJIQywcWlcErKBBU/gi93HV2yJpMNC32t+p/jrd9k
jP0WXuW7f3F9q3fpLO0x2+IhY8pfCvepuGy/md8ET3zyZWJVsnQsQH2KI6tPjchP
7eRdRXoVszZrGp6wcRD1NnvBn0xe+2O93ZrAdop2RqhDUpKGdhdOw2Uz07VFjyQj
Mr1psi5Y3VEibGTZBqbI5SeTQtdECssic10Rc5r+fynUtLoUCuWgDVUWBwwkWWlb
jKo71+CFl7TVfanZuTZB12V/YtUt4uUUlmd++tYi0n7UC2TedpNee8kQn24PuxGK
2M3pQhUYvtdbzIfgGBy59U4LFA1ikNL0BIVuirXCmcAONfn2WtS6CGjcr9O0KvBD
agQegGpD+AYc5HSbpKKVoFJ3QobueK0VOV5BSpmp5gpbWyqtUqAqaadCg+9NvqT6
Tals/22LYzPk3ZyWiqNviJ61dWtO+DtT92Z0k9lfmaz+I1vXQeKnBojjiLQp2Rvu
ygnzNXLvFQmmuoZ5qptDBVhT3LJkbvHjriV4Vhs5psVXvSNXFblIxYdF6ClifHGR
UAA0xTTJCZpByPW9RaRFwCj0Os2b8Vw1qySEXoOU6HX3VPe6fJcpXt5JSKhPv35N
ep1gEYFuP3lZK00udF8Man4givQ2VyKHT6g7CfFRAz8QeKPP6UC5vuNAIzkc6OPx
fXx4vzIK+gAzzrEV6vJrorG2V3H2Q00Pp0CAwlWqdnM4BWckYtUwLp+5jZaLQhm0
wC0kq7HTG4BlZkkN2VkO8+3DMFv354Vb0QGPu3aDmy/NruCH6BbX8SJ+i4yLl0eY
LDdzvklP1PiAMxWf5aXsqNPXER/9qNqMzO3dK6bgMyedS1fS3qvLe5kP8JaLymFQ
al7rDzIlgMFMbSGkAhlZnmyLh1EBE5sH0KLuuBVJ/2N+xawx/S5otH0pqNcZjlGY
EsE1yTO7pPL74MZsFzobIbqcxJ1YxN8aos+9hLVUqoiLV8MuWL6m7eY2/RTgjSn7
uuQXXoRaJME41a7j0UZog9oYDqIWMMKKtOHilbrwSpqgfq5yKg4CyJ9mmxZkY3/r
po9diBD9OzfExP+vRLo1J6DN1Ii7Rk76BjCe4JPncD81UgudrOOm3NGH/ZaLqx1q
iZoaTDs+rQGlp4FNGOn61FwUplpfJyMabWDLsqNMDrJcqNy/AMekwHOkNJzEZrEm
R5Vw+HVvUKR/KwxjEE3D2sJMwzOJjeaCmvWlRt/ioH6U8ki12KWb+pSmQ8ReT+6O
3o5R6S1jEs25yVv2gtDfxqleQrUdOpxVGZgCB6oLNBBX0it190ULRUM35fXWCItJ
beAK6IZn4JAKu7fAX1Lc8aLsEtxlBPdiYOsF15kuFbCEh6mo1Sxm09u8oWYASUkF
j4eVjkTL+DOa4PEC+UEPHphjxADyaYxJK/Ct9HglmiEEKNcpQsRcZx8szNn2WZHS
DgL8mFqB0OipSIlpGnX+GWTt+lU6cR7VSVs9dCt9785r4p2Kx1xnGh6BtzJ4v2NB
0kTYnjVeBmyS+DF8iKbkrYM2xC5R4vBynSaybT6CC9H6JeMyax0/WFoKSM07ojdM
TqhoviPNVQdTsw4wHSwQgd/NeWkR5XdBrmZlafrcN6DKtKU/dJRdkmCTnZwv54BC
uTkH+9k5UlFsukax9JdqUZ53cLxFW6uF6eni1nyM08EHfG4pLBk/DUMjsvbwuHsk
inwjzB/87DgWU21TIY09G1WdymaktfCgyo/xPERMQz3YdUUjUREsoObFayWLK2hF
EisilGXEYx9s8IU4Ayrt/oGP8/GmVpNQfJWDPhCFfXEEITJLY2DZSNTYwKtb+51V
de8oTvywwOwPJI/4L0TblFXDDcr+5BS45OxExv4tSc2EGq2QpkGVgJVDsEufXqx7
BAde6B/S8D173BUFKnRi4WiW9y5DEjEaGQrfA5K5Qgeuylo7ousBa+PmJM7QBua7
dj2DR/pC//xea9QM3L/kYAtTTZeVfFZQBLT0mvbcedMRfjvMxHB4OJT//CqsLcw7
yWxb9V8ajGmPZ32p8lV7BPInHrVJoWD9/Ar74HCTWorHmOFZILOTRlwtevwCBiHf
YnM2AivxsWh8BdFOZB9BmYWwM514IsUz+TTh962Gk3vS4ZM5gPMjw/1QSjtpwduI
hs6BGUSJmMZ8bRNFDvlOqnQgBbS2+j3diIpLcXyzCai2Pe9JRVGZZV2915i28KXv
J/6fi7juHYRI/1MfqcyVaa9IVox8feAu9Y4tis3LHEqkloAjUC9lUAjkzYiy3kF0
MlunzIR3/7PXi1Ahc2vlr5UM6sK8gLePjh01Uw5LysrXk6yZiCLgjvpG9dil1AqP
J19ZWS5SrUSDtV66X8wGMKjfGReObMhzE6le+M28+Hz6WYNGGpIJBFn9NWsRem2d
AWwH7Uyat/JhyxjFSo0GrbBEbrmB7mXrNIPKym3uhnphDymAcCSDfsqpXS6KAlK5
F4hIQd8he+LAQPPnrTfxLSMlLpyrrwITzZillAxm6kRR2dBJ1oPIkfNHD1msZyWh
INXjpdx2xOaIpWscrZ7mi2s+CSkgy0SZSfh8FegU3dYy1+sxxkpIUnCRgFfsvHUq
gksteokGZXeID1XnsqhclbJ+j+lhRJYEe4YI/a7x3hmV7JVHteem9EqqVaSgkg4H
Wsz1TTUI2sVbxe1K/OBqjIR0/VEuPfB/NegVcYE4LiOxvrobnrEj3rViTvO3+7/K
NwEluKnUno5/zH8nyDnm3y8g2FFEkL31fYt2ieO92Ca/HWIydE4ltl9WyfekfEIi
wA4aMyplxGBmUz0wr7ToT0ovfl8tzyNbAEY2GNL8EbQknLROdpl18eIpH5O6hOe+
1YVMToD7i9sRXaw3uJDxOVvT5EfafZnyRvWbeXxIa0Yypi5Iow4tADDibTPMIWl6
Y3AxiiBqmWvBhb1H9EieNvTBD0vhI+jU0EW2REl+8OqIiT3TgmJYwXrO0jsKlbiw
OoXYu6m+WjVcOjMRKS9ygRgCmpbOOS7vzFekS6AUUX8i+Po4dCU4rvuBA9XUj8no
zqZoj0ofKAR8HSYCY3YIcGqlR3a5nQqZivEnopzUaBHvbJqY6Bd80j5SpiyuuHeF
TUXaz9kvbfzb2qM4P4GqlB2QFiV+JlDFPnJb3e3WtoTevCW9qzP5yN9oSfyJrGJ3
e6k6sMgFEf2ADy6H99btTvgWXzLtZvgmWVAaDBr7mlMYHcIQWrESqn46nk5ERRnq
5koIi+/K5dV5XBrqajoD3hpSk9QVr2TroajTec+A3z8hkMZMO9O0iFAZhS30aIYG
kuqEidtkaIsbMfe4DW3ZvEvDhSRMCFw24ODNGGf5ZuJFPcOJNUnfY1UYUSDuJOtB
yazNeUI9xnxbnlPtFRkec6GERkcOAmT3bTxzCciq8BlNFleNO+BFSrPmOGjBwvEn
xsBDxOWWV6pX9pBSqxrlMacJlcopAiYq4/jWr8Y3bz5Y1/2uSpwenEi8WmfMVuAL
VxMBRiOqz65Br53qvMm1vZ0+bhpRn0N7K2THsZmXkD6k+aDH4Rj+BJ/ITY2i/43u
nBIF2XYInlnmstV0pkOqFp+R26zBvY/pbD0BIxn8Ilo4vu52KIr42NcqLQJzq5Eg
4xXLWfqAQovUhRPpg4eSxFV2PdpD9AevgKpFMRQ1OEY1cidAw29wIN6vrb/3CA0k
ONFiD5+HgMz4LzpKev5urYRygKRZvPsPy4iqDnv6xe5jt5G1ZNbCybUdBc8Y0v2e
pnED4tHy4CyicPe4ta0ldgrA81CxvDFsdtOH1etn+sJMxpWkkCrdgeEg8JCxi1sW
q5sNSehtga2mcE2Eyst5zrkpT/x1ZGj5V8mmrVSaX6HD0GBiUCUv41xbP6kZdHr/
ghAoc6HF/PeI5yRE1iLYKP0g57F3FQPOkILPGrEsS2SbIEPdCWXu1guC9k4A59U3
UDsiCEt6dBvTr7jHooDoIKAr87JBq3ye5udLTu8MiftEHHnLcbDLDN+0MWBj1rUn
tuJtqWzSMzs03C/byRu99a5kDTd10VA4qM/c02VW9VM8klVAuw1LWUvzhQVBou9c
uyC0vTA7qFgVg4k2bshyA8eqlVeZl3vb2cpdLxevxZNG6Vkt4YEL2tPTKMlxuIao
tNwbHc2qMWsSGjQT+nij5YcFUroh1jFHuOAJSzGoR6gikNDRHnPLDz8F+5wCBBPU
a9CVCmqjessk6a//wrCg6NaoDopyKN/ARglFZ10JD2Rh0SnKDgWQ3oV3H3L8FI5q
ysvbsnf7QOBBfD8JKNBpvXDeYSOns9LIS3dSWZmiemgfvICWX1KFPC7VR76PejNP
3X8mzceiF8w8eR2qBk13Awsz82myM/Q84NzNqTSVpkYPOXqO+74YfIIRNZs3Rfgo
cZ8OhwXnM9je/4jV5imGSRRJQzKuHe6e086t5ToQM/cfa21JuicCBifY6iIjr6Ej
dWD2v+Am6sFcQI7YGboK4IVJEIgIpVDHqnUtKhv0LzLRLqAE5pwvw0R0Mp+vPrBZ
aYxbThIZKf4RuVhk1DtZYXamdtomyOBjdSQnecpgSmVp3JxY3YSNHbPSKRe+Bitr
Zh9vDWr1C2VbZnPEhZDvqOm6wH6Og6XPlt7R+1Cw8+dlhXRRdBUwBg9zpMejmDRU
RYQaXZrbuSk9kjMaliSqyLsX6aj5FDuzELvObjZ7de1GdBQJdCQdz2XvkUja9ivN
ukLYxjMfQWL7JHMhhOwiByFI7epw7mXnINzxFMSXPWq6ZZ8npP5nelZLqLdLTFS4
PE0Twl0J3mEdz32KdcKUy08kfdLxQ2CNwdVG9sCEyX6IdU91NZd0rBDefIX9Lc+L
CUxXSvEi2LK4KHQPuPuGb4a9rFROnTt7aLxmXFkWru2C9G2UdYjStx4Eu67BAugV
4A1yjX4vJqEdZU56tnuFoYNQpoxyZHbKNCnuArRahAv/xGr8gpFqbljeTf7O701P
wmZLy61E0h/udnh8t7i2mB3f+HVmUuR3hkRyIzP7+BqYAvrVmsT5mkMbKl+VXmOq
yEmzLNf58tnoNfXj6O8z5Hyy1Ygz+o4qbyeY84KiPyKg2vQBxfcuU9XV5bNmcuoT
Z7WJAKXvT87v/ABvoPIIq5nYHj2zPHq30mvqo3d0L1cvIGit9twYLbPVIWqkgnm8
nNEnUcV940FkJzha/p6n6t9sKIzkmnBIc3CWMSRvOOO5dZzwiuA57RRanrFdM6k9
Hbooc8EHu20CVIOeJhE6Y+RS8Kr/TCqPb3R7Qma6mwO2C5bNvsVM4rL/s0yWx+Ak
e9aiKxJlrv6H4wtnbwvextjuEVuIG1SxejEokUM0F8lZA92QZCXPCINgNdcDskjy
ARxpTvyJ/kFSCgr0bfZyW72KqY4LmBkIQQzjM9usO+m5/VnsSSfMmO1cGdK5j+Vn
w1xTJT5k6dISM0Y5/Jiu75JxdssY1OXEN128NoiIZwW9DtTmkarEkEsTCOMi00b6
IbS44iIsycl8JrYgkF71CcYEk+nQJ3+62T2ZxfwqC0WAE0s00MaqEgdrOsi/pJc9
S4Wvm9N2JwuJde6ivdUq/JjSUk+M78aBiejvzvv66EYWDGPsIONKEgigOWEuBJri
aKfsUz1+Ndo/nuodF3rxfT2AXJQcLP/nf8+EUih0lNTICC4w4WjloZBt87fnynaN
k+ATfuzIIn8n3Qsj8Jr7bz0B4x4o3QGLQkZBSBzzu5ayyo00M6A43u6u0l7auCQR
0K4sButyWbTx/EpTwPya9V4U5DneFbk6FvXBklS8ytjONBEDmILGFa25NclibQvk
HmboJouqKp7g6S5UvYi8uZtAuGskRzahKpX3AcG//5vxtHcdzZ2nqfAfCBysfz6D
fkVXHfZtdw8D1RoffY7cMans+cR/2DaduitR+UPjtnfPPo9XpLBEUdTnY84XHTVL
HWr3uhl6VO8MV83vUrGcUwctIMO8DBI5l1BTIHXLdKnXJg9F4Lj5g2LgbGm1q8ec
fmOv1fSPCn+FU5qxkrV+OmcycAzSmJFCBbh46eABqEqOwQsomIOv0e///TQKLYmm
uDWyU73pPpoyicjJ/rZbd7MrLEMn6Kbjwdi9S0eqDImUz8y+WYEfBCdH2tS4PEAq
3YC2eiWKfvGra8VK+bq+qIiMrjmfDuK058Il7SbxPab5UIaQdYqnY5V1TNIW0VBK
xPoG3CHcBolXgFwvzvO5rN7Q3H6XljGMj2E7gwi2evrxW/c81rYFtd9MkFjmz5wY
6J2+PJgmKrTkUu7C/GR/Os/IsxwY5K3wAhWQPvZwtDN5zAg02WOhjfflNfAiwHnR
8TDBYv7VrvRAez8yeam9IKK1Hc8LgmjxgaEs3CYnnsGAavDr1+X9OE4oCczKirFC
xRNvB0jamO/I2F0o/gH8ENT0C/4liaH7kLCLARyKryhTHBAFDVsGt7aHQebANYJG
w6pE/avB2mMzrxd+7SsL+dL5AbHBZhijRYesy4nItXbtKJsel4EHsqr/F5Yu1D4K
JEzqH5ARRW5lKSpNybcOBcYvev6MJqRdpjfliFJlv9mn1ctVB+oVnZGgBZRiEIdT
OhYf2kbtHoZOU7fXAorI0NTiuIKEcK3A4W5HPTbxvO6xgudkFgiQxlMFSogfbVwT
v8XoN08VZAFJ/K3VZusI4vOsDCjRa+LXCCjW6EcwVkXAqlrl3JydhwV3cGzm/j9A
i7Cbwad9E5mVlgb4htlZHtF6WH5ZijGD/5L0ht0EWuSbyMt0dfWO/aW79HWqmFjo
AmfrruThNGg/+Lom4O09JU/SiAc1+EORBuHCA5qi1E4zmom5izu3NwwMJcqaDhCX
Mc6KDDtv4J7s3UiYyIs4qg7eeHEGB7allw+J5H15L0Dgy+G7RCakkSCFxMRL+FWc
QJlwxW6DJWWn2WfhK7qUsPfdMdk21dyzBhOz8Dc6BzsomT0Z13cfQ/nUEM1EeRx1
aMcVvDoBVIZSCn+xEcmuNozRB6i4R00pM4d18IRH+i8DJBPe1HPjYykFkb+38iEW
Js1iZs7BvjbbVKfakCeIuY2eXP/KNThuUArX4o/9FM6N7O6KSuxkSUSD6S1LgTZ7
S/08AG/I8p1sncTX5n/JLq2wDWsNNZM19jpiEPKEn6CANbkMV3LJ5gKaSynWaWaC
0FNtTwmMgFPc4gArv9J8NnKa+O6RNxilHRUL+wZsVtp7MhV53OFE7bmTncdsXeT8
+tKnq13RQaWgleRbq+rQSU42QYHc5hVJ7N4jInDp1BDieWLlTDgjUdbms+VeO+4E
OMSlc0BOY9nnkKhY29DLPUCURrxy7QnxTUY+BiyWr8walYv6aY+q5gSJ9OqVUNJy
LH5cF5rmhVKeHkRIC8yYH9KgwjSzM9l9U6UF+nFfaXxwsmO6X/K1E/ucA8aPrWUp
AhQdOfwPChqCQmIH2bUf3qun9IsNZ0mLaYImD/1qliinfaXXkAiIXQoTreO5A8+q
YM3i+1OZAC23VLB2XpcWXTbBrAR4ceOfibqxDVoNXGf+gfI9F0iaJFfKiKn0UZ1E
TAz1Dji57ggjtJ65miB99SpX8bIeif4HMgcRfG4L/ejHTIXyZUNIbKkVntevw8uA
5ynlA5LCn8BzyjshPcaLWo5ZpXnLL8f0CEKEWOxFWnoGe9zVnNOI27C4QP1aX4Zo
9BO0/KGdFIWa8Yx8HqZTZsdevFnt9Evr2eZfJ0ilnfgUhdT1iB5qXgrY8LqAyEa5
8oP+tUNHfNCbW9rJMc6S91V+AIvZp2//X6ncu1pdA6ThUU5D3KYF1K+5UmorQcR0
sgcVzQDn3r37uzzDIBDs6pCbtNfL/ZzbURJ0oIVqYu1JKa9OpCbT+8ngUlIcSOKk
/Yj8d7xiKE3z1Fm1D2za/+p7fPsgptfmGMxSoooHOtT802SziGphKmpNgeu2P3s6
A9HL67ef3syg9xRf+fkg8aHj54WHo86TV5gV8uNSSvwGAN0oBHkSRbXJAB0h3Iue
q5+JjnpONR0qKV3uOU32rmZzz00WLQ86/2E75Jre/u9pjKLNT70KBQ4nqRc+RVp5
3muEZur/sj6oqTKqFMerz0YLIEK4sNNdtzk1z95olWbBAbD7En8sRkb+a5fAcS/P
ITIN0uWV3xaLSqbHS0re8hTfHs+wgdpDFR0KCWp0KddlVdthsQ4bApC7YUlhiKOH
9V2Eusg3879B5QcfPY+rMKBb7tRkhgFM9KBcWFRolmnbCfFyIkxGG1Q1cLlifZ7f
QiQP84FoOAbPusAVVRj75IUAuHZOLSIRpNLPF0uiR/Ku+qoUEIzohdO5JAWRXupW
RE9eCFeKa8PACuIC/a3LeSEkXQVnudR9cbwJXtNrzhCoEPFoJ/AihH4isLAGMBkJ
xs9h4h7NszKZ8Fzqe0IhMho0+WRj6uIeQiukeuD6CVP/GCeCGH29wpaKH5QG5if1
8cwEqrN7gxS9kF97j/nwAVtXVnXs4Ii1QjP7JPaHVQVoqoKEo8Lv753iYTzzWxSk
KD61Fr8/fg7CQyBF3jdSLFAQvvXrfFknjsqmQ53p/iVLHsta3JvYuEoMCtHD80ZS
8ZgVLhotFcMKe4gc25x7glTz0D+EMdCy6FG8Jwj2odL4WJy5Fy8VYpkd1NNfNnoo
iV8WlD0w/GzFjmuvHM/4QOUNaVq0Zg7UBIPH03K/To5WYZgGN2VUjUScuR8aWuq4
FYUBBxAUf5mHF+Ta3SpUaSLU5thcIUi4WQB4VBH67rmOzXS/A7NC+rLN2+KSJzoi
cyer+hmndJuEiijXXVeDpw/Vv9MkdQfsh4dNVkq4/lIkelRTezSUH27iMF8et0gn
i4iOQFY+iR9Q68VROYk0R+NzIeC2imLxDoJQagdxSbBX/uMx9rbVJATkvfB9KCgw
ymq9WK+rkCQ7e1WxqMdR4QA7fx565Cl8W8d8q95L+NREDMMD2cw0qr5JAhhzbT9T
jgzp1naZSFBWTC36ANOiLk8IUdMR4NYc8GqzS5YYVe7lIu1tZEplQPpUQ9VBUHlQ
KpQlIOsX7pXlu77IQJEHP8l45StuYvXNdimVl9zCn8hyuIruJtHFeBpCHJTok8R1
NpbJQXCeEESfT4vY6QxsbNbcJFzN9VzygXTC398KlL9uNwGm1nKq+C/2fqN544gT
XTmxJZ+rfxm0LRWSEmAvZongUNJrnxXnBBgnA4h0rfzCchDaswqUysk1EJhK1T7H
rD9ixsMtVfDv3RThn4ISii9ahmsLHjzkIgJvfOYkGsSQz1N1P30Q6oeSSl4BGazo
kkrOjaLl3m+tYRLg1DlvwuSNYTlEuC09/ugVxMUhu//FrLF0v7YFzHG78gntu3F0
5KzLd1BYGEZ89TFJ6i0a14gthEb44el9/zDZhKml1ghaw7bxsvk0+TQjCfehV0TG
VPxYv9xChjEIeJ+4hM09jGRBreoef1CJBScRio71Pun8J3dFSW6I1zfLjG2yPCeT
cxtlvlu1DORKubDQXxVNTuHeM1wszz4NCphZMz+IbL1dzM3SKj/XO8VB2zPlUnLE
cXj8/Y4/8i2zedU/AfFmh5nomuFsvl8PG2bQjDyQDHNWVLGqoPIxDZVlKlnoeTD9
VODMouGkCpw7bCxaadxoEzMY7+Nwujcxx3Oxcc5nAeKfRq4ElTEc5ZdW96EfXyK8
BEdfXmUhSYc0FJbNtg/Pcdm2rzQI5XA3B8enNYQ/k6R/24euFCjjusbQlj9KGlcA
rs1x7yTzpUa334piJLtUS64kmpfyDNRMw6OfuiyxR6SScBCbNFCccY1oh+J1Bo6C
TJ8k5pSDzuF7uwm+q3NRVXQPYLRhMMSux19kKJ7vsDJfLDrBWHfKsEk8cDCgkPQ8
19TMeWQLQTFMG8cHL1hlviy9b49f90KKJZvBXirBG00KLsX5LqsKdbqaoDKnXXus
MXCrUtcpXktINLBK2bvgaiP0TyEmrohQibiWpvm7nUN+e2bFmcj+wcVM9jZl+43u
TXtz81FO/+/N9AGS++RKCtBFxFLX7V7ukwwpZZytZkpIQ0rO0lru+6RLYuDpQ2DQ
z4lBafO6BqJYBWpcnaWrJ2duy55NWAxQAdkT+1Kc7I6lN34M72I+4KRi3TtZCC/t
rJF+386SUpMq3HqNVbFCZJZycO4baCgVoGuBuOqoAbvIa5Yk2WC30XPphtoKwVJG
9OG7uAoUNZgcaoDQPlzLyrlhjabEMuf2k50vUe0AbIXanKHn6DGt6pLMCMXc1O4+
z2xXQE0gYI2PJmWaELfXT7yClH3xA5txxfoeqJaDOsoxxtU6ZcRBwhpnxGEe1lZo
3t61SNNKFAwaOJRGvk6Dkd4eVKTXKvtrHuMvdtbErho7VkGzjnFzhA86Ccf+uVgI
5YnYfiybgVipBpBsu6Pc8VrqMsxqKliE0XqZTOS6+roj6gfdXuyEtm11P1XR0Bpj
zDvK5e9uB1TpW09Ju6vt9VFwgqmYz12LCReLkgvBO21gr/mjTgot9+o9YoCQ8cJZ
cRlH1ybeome6IknTSCZBtRPDI7Nzk3zKcurRC+XQP3MsCv/DcmB43SXcSCSKAvoG
9RoyFYmRXI+wbNx1+hsDBRgm2/zWvZ+eKFb0nLRkoX2cqcPVaGT8Ld890mcly9op
TwZSoyA/yXoPx/ENg2m8UBsMJurrS3wxeg2VCZlseTfCRNQk6+oeUfyEyjmG468X
5jlnc6dxR+xsC9ZNk+YudPJOPZP/rDuebMrXw6VlCfIwmBXXBeQ8MEN2SFTnjANt
1spZxxon3R1aqQMIxeEglmWt91UOs9vKAD7liulcVynE36WH2LihiXCNEJjk1Yb8
cU1TU8DcaeZoi9Vb2zTqbBzgDM+9s5ElFSWH2Ht4LwXf0klxByA3mn8+3WRCcIih
nBSaf6MCP4tfmGGHEMxBIjRFe/i/SKqc+apI9LjDRw3OtqUFZRw3avqjrGaFXgeM
1VWasFGtwqWC0sNN+Kd+qNtmtzu79SldASNpL4hpmKBdYzLf5zjczwhNwtt8Uk2s
40uVzsQP93roK9bkVl85rBhAttF0aedQ+7SalB2kFq37bZom9VgYv/5mizI8LxrF
5GIfk5KqCfi6liBjLIeJb0z70t2Kzl+nJEiCLMr/RrRQlcqDhFmG2/RH3ZiOfJyE
YlTzJRakzrzEu+STkoqMzRPe/OqrvmXvKgiB0CMOHDyhRTb8ez0jrJpoX4Diduzo
PEuvTWPtK1Yz06T96I0kWo5F/PL1kC07VtVTYeJ3hYw3U11a7pkRJyqp/9NubuxL
YG5NIVp0bSsDzjBH0zN3xZBhEi1fLGh0dj0WrXta9O+QV55VBbpW6/Q/3QTYpbqv
SCONOtYJdQspkA6bo4dhcqCtA9JvhvHoo495BSfwyetlUBl7e1iMbsSDE9sr9/Ot
c77Qjqd7t40MIi5GkkDRJCLHWEq4QRWjAaZhTn9j8GrS6ss3IdqbRW+M1r1FZzfg
SwuuSWrUTQtBBxuA1FaWf/EWp0WZ+AXXMr6BtQZd/4dxv4AO7wRMQQpwEN/Ik0Nt
WiLaGMJdHKzSd0LdARum06SQjIKg6rRhLQUXj29B7RE3I6b/+PlH2e8xzJNkRi/s
iLEPKGfAjkc4PMhs4zomY/uhUnLXvAXRY9c1uKZb+db4YU0/HSgPuOT9IhiWsygU
oUdAWuc1xoOf/0L/Q3EdIU/0Yac/hBcx5APrnHR3LFfgqBfaHR4nlE5GYqIo+Fdy
QXdy9JVbNz74Imnns9esCLnkSxCxXfY4uEdx/6/UGxeLkNXQBWSKLakjkZzNcyVy
DLYIEcFPPOkJXJ6zUnHnsZFrDKhUoYKRRD3CiXOJWM6CJuYWlrKgMsIVSSG8049N
8a72Ba8tt6hGGHSIAlfdxqB0woxOz72DutpycgxvnOHg1U5DzwXotsWomjDcK2ha
dL6KSa6+o0OcEs2XEUnSrNB9RugzKliO7ZzvIstpVj2ys3iSDuZt6E+wk5ahgblV
w+kt8VKbq2e84Ku//Ucd1HSsBRFC0aJlJ9MysJph1tJr+NGMkNUU6X2DMM3s6418
pscTriGTV0/Hn6zqnfE08IHzFGEwXj6+shXMzsPMyl/6b6cOVsknmiw6yBScc9bb
oqV91f6Ufn2AG+6L0RWNy3jYTY/TxP4UtyrTUmNAv41zHB8PkHJt2wTNO35ejmfy
btpEgUFC8Q1SqN5dIEODOGay6vpwLNarkAoLiazk+p1OmnneiW0y2ONUIoWEwaZ+
NXHiwFBpFEk6PV437xThYdjO7MSQ1E1mvhmt99rFPMv8IFB8a8PezPnYaGAUOGrF
GkZixU7sIf6he9U4wfjBzmN50BMwc/orlzH7LGNLqswck34aBRkk4Vt8Lj5FFNTT
j3ZQ2CHpkRPcHrpKLH54OI6vdziQ4pjkTGD6q/0kNQBlZoiapHBw7rr5gJyJPug6
IiQAI8RN2ve3eF3w5MMvQLDb8evGrEsspYmcDBhEgzGdXrcWUeweAYluT8rPLdZA
xUI8ypDL4Yrtrrra60p9lDx63IJCNGNIjNJJWU4WdvBCBTeUoutjpycJLzr92Q4v
mp2JwaxWeH83A8Ix4d7xl/xQPyBPD+KqDWcS5/XrZagNyRl9uz1yXo1kHgeWWNWb
xaKQHMFgaeyNeAhUlDW5Ou7kWC6AQUw4EisTgSa5EaeuHjysdEwwck6og6maT3Qa
XiXLIMpglak3WveIiAhjB284iuM3Jh5Z6yY7ONLKZPqXMp9CVVsiH1PO/gfXEOw3
H6mQJRrdwk7sZ/ZenAF73eK5MOc7kACGShbag0eE2dsnkZsIFjfYSl+BDwKaSbEZ
k95lbVGWCCzRSy6WTKDy+fV3Z0hcuLJVd+tPO3DhpZCWknHURH726PDymomeE2ad
/kGqMkMvQb1HSIvLYNoBSGZs1OdMtuCCHUC/qIisRx+laK2pv4bAc+jwsR5t++Hx
9xlaECNrsaMmUWvzx860lERHlebDRrm3ENvFnRbRgt0dqQ0m/xduPWqKjLE4ruL7
aFnQKvMC8FtygPKSniQMlYDYBkRSYebrt4YUqtHSE94R2Y8ifBujfp6KvBVn/l5z
RlloLYzdWmM5hoMaG8dEmoPWCcblinYdjqX7CBoPwGSCnUF1d/CiTktIAZmxkuAc
MHQ08EwbNqPzF+xX2ZiN4shHNuBwghBZTryusDfGhVtV5tdKXGE/QbtsmbOYcgXl
C8WmygjezB+n/kiyPXAsbFU+k0XYBsvzfWrP1DoF5T8j9r0Axa7jd82jwSpygcFD
BbGisy+tw3H99x4zMe3SR3HLKBY4Cr5/2/pagr60Peh1CCnP/j5Qzzs5ODO5mTt3
oMYcyr0INhqAlPlcNhVG8oO0LVFzQWGKfKSH1A34Z+VZu/S0YnELjb9DkKypgAnh
+eRQ+Y9CmkENfiqG41VZtnz0xMUEcmZ/nqaOf5zJg8SsXJZypQSHdXe999VTtCp1
xT2wAjDRykfBrxu5j/d7QrFNABvZNIHz7c4M3ERGl9F9vYfMl5DnP5ZVvyFAnzMQ
SUtnEBk4urA3a2J6bUql/25ozpfdFEY2bctpSD6oFURQV+BbjMcdPOaD/BzeZXIr
WHbeYg4Ny6YUVvI02YtNKkBMLPAKx25fMJX7+lDUihZsrbC4k39SIZWag0M9AYOF
l8/fp7BMtRyEgGtVw4W2XdE7pyKp7aRq/4Muxt2iPG06Fp5byLVXNdZvRVldmE/A
X/OpTvpoBIDHHbZx+TykZRZyPpkrReorcdBfiQ4G3T3Hlgtpjn2EXmzged4TskTj
Mi9k9StKcPNcuZP6Q6ZteCm4Q3xcg9WYzkf0T0C46BusXWkmuycaF3dU53p08qh3
MSUuIvGmvVyiGkwRnIRud24Xjsw9KvcYR5niepa9IMURmO4kNgXqOetn/C67XF/R
NL+EMAYP41OqyGXB0U5sT2Bzyl45Tm/B9ARerkMJ1OdEvPZxG4HQCu56wgs3QVLn
RSMnQpXOFGipR3iyIRn2X1BaryhgjYeQW2Cs737DC/r8PeeZFpy6XoA4rMKzTjeI
MUlY/4cJ9b0WHiSmJJqrsuW8UJBo1y1Wykp5UhB4NRIFRLbwWZXRTJDSqyFHn1k+
bLqYY+dAT5fQ50ISEju/huFhy4rONLZcwiAm+FAf+WF1eseTQZ+idLu54xElUPL7
j0FB4hvJ7SgSjDd7xhv9lAkRknFdYLJOeYCKnk2XYJnuS2oYzRdHNg210gLj/cZ5
7yB6lJltUQyaM7cw2TSM2DQKp1M+QlYdVMp8pGLAI00BP9U0zN8TwCrXOZrjLKA9
QiZdlwqizqH/46UstNXHb7q0ORV/6UtgiRDfWP0Nw6W5re9gKj1kbCGe+QJ8Lzfw
EA58lpsh2Gbxl3Fn7GKpweK7UPqvyEBD18pHBRByPMKxugMoMJOhd+Jnzj4flt1J
UbJ05Dh2O6WZIkcV8/FkoOu46aMNLiofTUSuixyRb66cwIWelWf64uZefk6h4Tmt
lXC9TDUgeVOjP8dHqGG4kzhiUnN/3G2sMCDxQhaNG7kaANrFswsx/pexrNOjw2vk
iyRxiRfdKlfckm9Czo3xZg0uwMkbDIB4ESdQiwI7ZU77YS6bBeeV2sE2mW0+Dydq
zmT60b1yI5c73Qpndd3GQ/RpjBNh2zhr+sSpi0z5M7o5OsRI2vjsDM50/67PNBVW
A+o/EZTomOg9MjDrT8eKSciZf5KggaRRNbjF4/DAuy+FBq+/19KjF/R2Y9mx+o+e
9XDbkBW/Geod7smQYxE2aWHpT2EC4UzZbO/0U1kpFrVznF7CkHOAmKojfcS5jfXN
utwe2R13SROwsefoSLOznkoUaS3xTaI0vdUWz7RUceR70djGNIzK/cCyXMwyGYPr
qsJa95mDLbOB5qTG2U0zdkUs8M60Dg6/m7bxe8vnZfaRTOqMOj6WvdO6JH99T7/Z
08UUiwY9APgSdBKpivMkWqavYI/q3HsaKnEoW2JwEorJCoxBCjnny8DZGhzYqKkC
9NI0DPbixGNPb09o1CmDhfipwEL/86uwMGxkk+O2nwUACsCYFFf29MBZoBQ6Ldqm
cTN1mQhh8iZjGiWaXlGEJmX6zHwi/n5BvARwfI/M1TcI2Oc5YOy8nW27l1JrOsc9
SUrpiauL/NSjnSnO3hOsmpmNQR5ft+836SFRFERrnW2xerq68uRo4K86PwXpvlu2
1S22bv1qMUCIFJsTepnvL/or+HBY2Ko9d3pFEOHzn6eKQyh49hnNcT1KSNuz6Imk
h5UBbmiL/0yXgcP3wqEY+xhXn4mX88u7sB9ZCVN2N2XDvtNDAqrsP8AZf6Ps5gn3
Eiv81k5799KVEXxEKudQ2yV1Uf1+ScK3QNRXHafbRcEZEb8r96P5z4NBL6OJFzOK
KFgOrXGLaNKTw6FPy6pdebmzbxYhqAXBQ+kvaK+yZFc91HSxz3m0vVEPethxLDzV
DDETBjAcTqtNva813loctUvmw9ERMBslO/oDv8wyijJRhX1NXjSIemUU/ntJP1A0
wEnzUfLcJ0HbkIAraVsFMDEAFoBg5bweVJpL/U+CowKK05UwsUo5eal0FuFapC7f
PnXNblyg1fclBDJr0uQz3ib+dBOBip2xJKWG9x62Xd99vrTRu+Xa+Pgpc2kRnPr9
GDyKfMGhW6pZT2EaDQSDsGHmv+o6g5NZ58olXgPtY0Mf+9o9BOdW/H7JFU3DEsQc
sEUBc60jEjQChLlEN3P+FJ5ubzfnOv6X3CipAUeR676i2LXgCt4Csg8CM7Mxbarr
T1vkRdwrrT4PJgxaDeFo+SInsC5PUD+rbdOqDJTd0HBD7UPO3qM2hEavwf8QXUu0
qh5M4LbTbk7hzXG8xu3dT2Ak62CWB8yJd2d55Fs0/VNpNW1V/o4ATfI0DGhNzzJE
9mVpZZj/TbOP+tTvvAb7khCJAAYOZ9vM/du925/aDZASTSYdayNA8GuKd4sqIUi1
9TPQE50lFAsarLLTOm7Dqj1bYZLy9EHS6+NIMzZ2d93ZvkeqKn8/zyv/YqByTuBd
tBSZ/jmgIybosDMOdTidnfByDgGrF+jhgT1dyV8WzBtsoCRmx5A4rDaKBK8mUC5v
a5oPVcZCXL6lNhH6LkSZ2ROupR1HefbdoPeez+RbTO88FInlpLH8WBMZ8BzXJt7g
nkrhmPp/c1qkW9qKd+ulAkAJ6UNTZMTO0MxMLD9lUDF/EQt0BJPjA9dIRSjrsjJo
bif6SKekmATennTmhie/aj2cMZlnaPYz9u77wYykBN55VKkBa0wzKTKhNWHcMjrG
gnNmIwWOkoaJ999d9gGD79F5sFg5JZ1xe1rK7xDodwRBExYedUMrh5hVam+494SB
KkO0Uqt+T9nH/JWKvq8aknlv8ZWRvHY2evCsgptAxi28Zj5OCc3Z/nPeqFSobopc
8AxdRxhBSCYPi9pfa/xL+0YTIvLFOJNKRApFayY7/Tw+SRWptvl4T9DUTGbXywe0
mq+BrfrDDxO0T8qqxfJIP0P11YdyDHt2x7CmH3Mi0X+MnzK7Dr731SV/1QqQbiIV
StDMGobhx0zdj7fqPI3ePDpN+U+gwEIG+y6vmNSL3JPXTtuomioII3hnnNTp1WeE
XihTyEkw4l6eCN6exA3k6m1q7EzZo32NYxprsU6R98kGe1UK/qb/MpYyTYZhK+OJ
hgiPfxGqDdea5tw4ymyevhBpqJorIqeNKC2ptfY1YGKQAwx/9SG/zyQCbTbS8o8Q
erJdzvX7fazyWIEbgvLzVm875iF9thW9ACFt1EbWgqsbYA1BIQvju/50W+hPUyyx
sYpTXD7JdrAP1Cf2d6bPJ4h9gUxVShpVjhdqAC8H+lO1NTlgrzn6xrKZOb+vcUqi
B9V6E+v0Bicby88/OIAPS0o3uilZCbvqSHgY54n349OaUa6DCxKd3gcozJLoZUzF
PA04466JePhHlVWkpSWbTvJanrwu2HR88o9XhRQsjuhjjW+96rbQ20UsT3/Y0Ddh
CiwMrG3vbfVjRMvLgKFmrMLF+2Z5NfjXaWJ0hmsmWJ8EPUhxsIIBm+f+ry7LZobH
wiDOnOQ5X8MLkskYWkdslj3j1HcnkHT+vdk8W8cIJYFbRPLlNmo2LhISOR33wuPu
SYGdo5qqinUQ9UoP71cLthE9tAoAKAZmX+XT+jCeMvTk3hRhqa13Ym7XZLPBIVFH
W9bOBKHf0iYVcYK1AbYK1x2LGahahgJajyRqboL4bIVub2IqwJ9qDtl4NsMIYnNU
it3Klcw+aYDeLsalpwaNfqVIoJyxiY/n63ZTJWVjtNAeM59zxKHN3M9XuYjgVRgt
GLnhRmu0x3rm0Humsw3FzvEaWkexLWKymA6QRzhyF40hXrPkz6VDnXEHATLQ0dnK
CYHzGqTnPWXywKOQtmoSTX1COMHwOcnrtdXKLyPbRcMn/5itlGnqfeD7KmvqupTt
hrac4nM0sKRry/F01Lep6vNCJXzf6s8ef+adTStE7ks99VFlLXM1NB1chP1GpbZU
3Hw3CoZ5NcihOj/6AGkd3uoO9VkrqobOTYU6zdSXqXvyl8gHBVwckyxAkKNK7JDF
9NhOHN3nq/oLx796deRUhibEb0kXnf98bg7acfy/8BK3GtLDB8Hd3MeGleLMYNW6
mR8zpi2zj9bGwaq/48DOIpO8H+H3/CfgwBDwJbQsu75DJSgtWXZ/TKEZNSJtCwe2
kWd9mYJjY7AqkbCUxeQh7kQlwkGc5qw15Kguw52jNQ6chviFcPdv18EiponyBGbS
HU8Ysk19ywORjdh9+QXINsmtjKubGBLcSIf7S+xa/mw+vY9D2dO63uD0QRjL1PXB
saPgBwjlEJjg7b+yOCLsFNHwtGgClChTIDtmgPcf89nLg9TK9/Q4rLd6tCmA4LGG
hzGhz2vYf5k6GWAzUESjJ9qVmytZMpL8OpKfXVW6paM6MS2+29mU1sf922M3QFgC
zluNF6Rs3u67kqONbYXzoGuOK8hQQcJ1L2tVUoeqnzIMI0e4ORZMqmqlH5BSMNqi
XOK9Gb7pVHsDbHRYaH6QcjgXyHx98jbAU+0SGnpzoC9VV0mVWPhSLDqd15pdZ7qK
KD6d2OamSw2GU10iS8G/ichUD18EAr5hPv3n2i1/K532q91aSO6aibcE1+KZ6jdn
FWJcwWvR2rismbLLAgnyNZ841fUYmIsjPqim4vR4QPRoipEaLqWRETgF1lXGo5Rs
tftXwHjDb7EofvqL8Hpc3H9WtTX3+S7hU+NHfMYiwCEtBOCoKzz9AmkZS2+eIEdC
JRk6i+hxY1UAT8+CLm33cvfXBEYqO22uLlttaoBUaKh9QreDM6O/lenUuX5EjC2v
X+evcgiiDcVrYjkTkYI6fizoEoMRLzJH7KV+1rRXt1HJug9S8eEI2r3N4Z5XCuzK
O/+mjkVu1QE4TgeondvzsxFHY+045aCfsMgGeVNVZFHcsmK7Zcb2p82BLXSZRg/Q
wKG71fZgT+AYY3RBOPGlozLphmFTb//xA0q8vNBJPq3o2UCAzZ7PUKX/Ebw+qTBO
wpKnkxlnBaFNYNIgpDkOvgS+B81Uy/EDL06w5zFOBVVQxGy25zQeZKZZzts3l5ep
KkqSSph02ZC9b8fLhdJDJ9hbLXHU/LpV4pWRC1H44xP7vq9sd1IM5A/5PmLG9o/b
P7kWQTHXjFF5sxhichq2wdQvBHvdjgadP20ulODK/rSGmu2cnK6Mni3b/0CBwM0r
udY4d6tvsfNxPJAKKdPZZemQ0rbIrtxhv8Q0B540IlmMLTgIyoYK/0Gmk964qMhq
0s32NRobP2JLTap2o+T17EOnnY/bplbv1a/LsEOQKCg3/ghhujpYa1zS4gXRc7Ak
acbJKeAUVw9dw+K1yaB34gGkw4MFfj+tTmndjIPVbOC+HIkmIWv5o4WXlvOkGR+S
CTSUtPhXGeB9VMGKDIlwv/pDMWSiEoikJ04Bs7TIIAbDmmNm2Zqpk1CVutCZgWT7
vuWT96UGgtiFFRHIkU+fumOEV7kvBQQmpdCKyyPgmX5dkzUxOhM3IR9sq15IVpjm
LEMiFHvc0T102f0QsgGJuDGfk6mq94vgenyqScNYzN/s3c8tVrubD6RV+F7wSNga
gqMhxMyD3svYFVNJ56+lqJJyAT/fnnI8rwAp0FI0e0NLZjaEMQ8uUme51L56BPFf
RdBkX10rUaaseJw78bm8YCaOox+MI0Gqha8Mmyh1hkf81uGQ4bOi2x9hgVMpCA41
s5tL08SM5o69MrB0g/SBaCyxbCFYrgo4n490IBNn7WNJD9sAB1ZrvNYncvCp/FF/
dwf0TvCLxhEy4ivZSXq0lB6L0kIURaoUuC+Zb/cx4Rq0KrQPtmiqfPFT7cAmHAuH
0lOtb7UnT5P/sOCjsljYcE7/i2r7sDGYRJTJSf7j+DNNubvnYiPym1ykfniCM8Qo
s0kExrD89JJO+08qQRs0yiEV4sXUzIsXiZen781eWW3xzoyfmKud6u1KjAz5zfZB
gMOreS9SRBzCYKJvU+RnQssq2MWCiDCVWyFDiXI4PpTMEe9yah7QWEdQAiSb7pTv
X5sSYrgofas9EszItST2xDo+BJTHhB1tmj0CR75VRQtB89Juvv+KJT6UXEFFftzN
geARbqXe+xZyfNiBZNsHrdBkZefbjEHGkEV5xo04V0o4eJG287+mWxLCBFYOWvD8
uVq2MeSzNxMHdrBQt/r4jgvdsFEi/kowllqnrqs6XdGdkhjKaslFo0Fb7Gu4pFHe
28W4uu5Mct6Qs0Cc+qEToPTaqkw6sPtRfQfzCfvLeoXbyuLNgjWuEzUKzb6WUYMP
YJyd6ZQc14YWUldRHGM954+opajbBMGpCfvVJj69Z+QW4roJgeMwbtuBrNatMCRf
bGy3il+hwhWHVke2eDdShFCpq9W2JseB+3Gf7rZoP/QwSTlnyprK7+E7vAWxva58
FmZVXABe6o81nGzsPbwpe8h1AhixNNT7asEyJysKxpmjvzhCOOpRNeS261mfn+bN
ezSCpReDEZYzpP4obgSn1b+HLK0Yfjr2m8NY+yJyy/OqaaWNTICIO2uxVfTxBEwk
i3n1sVF8qUSvg3Ubr/qBlAuWqFdzx/BKDxpm7G0VDxUtuKvMdXBfxl/p/v1oyZ0+
vqTDFb0k04IHXRglc0WnQW1OkizvHssgYMiaEAaJMe0/vHRR5JKPDwc/4KlK545R
0/tiebFv+0yZhP/k0RuHuT/YfR+5M1sQ084fk5m4xssvSTzeBx5WuWX+v2T2ll4/
3/sY7M9rVL6Fze+d787akkEljDb+MTDaFdw4pUeujuwD3j1iWH7qD/87uoK+AKXH
ZmiFCp7MWdL8cPlDB8XN/GBr7rYqCvVNBWplImEe/rCypXgXSn0ITN8fn75/lU+K
2hfU8/yeLhKUU5Rafkt5ecwRM/TDnfs3aI0kpsQq0il2DeSOWZyfgENS7PAxxKcm
4MImnrnD5bJhcJAJcZwl7kypioXRt39/hV1+1diHeoUVl7rw5yJcI74SDvWIo87O
hlqjKGLlV/wqqx+CNGDnI8ZDO6w/4c+f8xk93lo62iFtRdjoMZULp9fw/UBm2QiW
hYr0f5TEUPL6L2Pg2fs5ANopai1oHLVexDX0scAk6oPh+E05pMB0zZfQ30Gl191W
wht/wqro0/oxVeidjMIb042kCLbsKkqmhRwRyn+GL3WUD3b4g2n15kak9yZdN081
/d7NdMSMIPgf9Rw6jfhUh5OZBieaejrP9eirJnE9Znvwhl4wi5vULDAkhQewC2IN
gLOWx4Cl8U7LTDJfKL3bvNcYN58/yeou3FYM1ykDrlSzrPam627lGKljbvYPdPQ2
LsAMXOGC3QJA19dXdaushh+rktV2pExm2DgvauAw+cn01yNs8f9FNmZajG8+adgf
YU4ysTpi7iwovVyBK5wCQbuWSK7a5NbCLFHVuQXcfv8eQlILi5YrvPdkiHVJl2+B
ZejvldGpha0bXO8oVGXwF2X6vbnI+ZYazF2qKnGngMzcIsHQeGeW51dff5xuKBXX
96Kp/ujBfCGZLUcGOf2nY2tDTO63K00gEiHWkG17Tzqp0sBAgQez+G8CF9tC+WJc
a9/ujTlddRwyAZKjzkgHCQ6VJRGaY0chEgxd/0mQFNUkZCAtBfnQ/0yiSeUsfEmY
6RrwUNJxBaQgflpiYJJ2JIxGGlCiOsjMCwQw3X11dgC+hySZFTmG811Kr+JWbb7N
27OHl23afqh6wR2HHwAahD/kSgOj0fthlmQ69Hw8BDS9ml/Chq+FhuRfec3yAlqB
tFXYxNzzKu9VzWuyPbi0BV9QbcCcD1DvITe/q0XN/+yvHX3XHPa2Zsy7CGoTTFgE
iYF1OTDR3gy45tOyZB5sHrZsXDCUIToCvsW9pUoeRyX6PJQh/a8kjq3pfDTOcQv7
z/62uqbyK5JnQ547X1WWTc4l1VaYriuIJVPDo80MABuB118t8RvGQzuunvYfVAGq
txRIMU1KDyAOCza3tL4wWv/uBCtvH3TM5tfhDwocYiuR5W50UCP3J85VmYmorEDF
pWnLSYXRx11m0xXyF1oP7G9hdRSK9dwTob20oI86+gVB5nyVoKIE8lw+uO5I9sPO
IuJPtDIzxFMrnfgyPURDZ3MbgRDfTtnLfpSiZWxmPo24WWQa95LnBMU2swKYWtoe
HELwf2zyQ4bT37nOFcRk1dJAbzynQr5S/q6+ry6d1cIVvJwZgSpQZSPua9poTHTJ
auba/pn9I91/8hOsyr6R9AW2dw4XKrMU1xs1p4lpo3jTaZcsdNl0t0Os1K2zjhrK
bqrr6fVlEl1ETvsiI+hAQySCPohTRV4J0Pf7gLzSv4NIEa6yM6j2s02xBmnxeswI
RUBc1gQAqN4KJjMfVFQDPe+fyrq1QPHZ3sOcn0Kl70FV38I3hDUvoWwJ83QaeHVf
54dZOIAU6iEwlUx2lfh4+iu2vNTMdc3Q6k5z9EO7auxfyM49cHqY+THRXg64GduA
VlJTPxPP5iaI/LvfoU2wCHewiWF3Oxps59dwCZDr6ruEdECTryIZNGEaKKw9K7ks
PdRXOxhrr41kJFnCziAsPNhp/SwKLVAGIh34Gj4Vp5Xm/Q6whOkpM4bGm8WlsGr/
hsHudwVRy478AU/MEXjJCNKqxLfb/dLyfVDxXMlgMGqY2HcdODl7t9SSi5mBvOfA
cRqPc+OkXV2YEXsQIQWjAwoF+KRLY/xjf3mkzSu+/Ms/yvilUHdRRNVjxJb2NZwP
ZRaRlwt5Yp+I6PsERM1ggKcNRQ3VVtei1hwZRb6unWvSLqG3BP54nKKOH2Dz3kOn
1vY7sz4p0t14uoLUrqY9i281zhIz9cSOUc+wQAv4Z3Vzzf0hIegdOR0UjUnuXegG
gGLqFgK87XyERvQt4FiUIz5EId6EUa5yaNjIT32+PiduHvX9cUIEN4zBoJF0iHz2
AgWdl6vTf3KlVUt6TX0eGg4xvA4qWV9O6UeHCexEB1pontwSYnUBR1FiyUM1XcaZ
2x30z2VLu+xh/28rqEZhzuGji1zsiwq7es8zBmdi3GUQKqSvxMLf0FVrv8OncW2W
LMPIJGR4REAZ+MV+swVwz0r4mwfzDFo4Ns4oXtseB+/jW7uLQvG3YP8+31mFqdt0
jq+SBTyzqFrefFu7a8r+pHsBMAkBDwj4aOjCk6J1Vueqzz7AdX8wlOzYH37WfYvx
mqHd2omUpLVNUPqtX3/hudT41dtuRuYf3AW4MtX7dk9jdKkKWbfGAMsn84SyrYy0
Q4CNFbBQ6AGVnXtYr/t5ADCD1hlgkoEb1h/me/Re66ZRJe+sfWAqLK/h3ItHS1X8
DkVEhMYev/wxBsJzvUqk1pR3lWcVp3UTmpnHDq0L6Dl1QPwtpJuAWlC8iGH3recR
IDjLwSb1CmWjfN9CvJhCXXYvGLvL+Thl4ooDn2riw/hRVOuQq8Dy+XRDJp0ETBRL
m9rN48ZuxoDsgsH3AfpvmbM9iSm/NbAyA00AgPuhOfodhiswrPKXyJS/f8NpdmfD
T2Ea5EKAYPQYHWqzF7nXO82pwfPW8jRHarQv4yl/s6uhnl3r1+8MSoghDZtzGyGY
8g1sebR3gOCLoTXWBxQVcrG1Wm50SNssxKWS6VXvTPp4oCpstaLKqRI9JR4OvjHw
v1G9U2DycFJr1NMVeLSVGyktEcXu7nXFYBFhvO1zIqvkJRbBB+gX4vVArlKgl1OA
A5hD/UctmY+Qfm9AC66lJL+ST8tuh5l0aNgmG3bGSVEpWznl7eXDdjIW84eASWt2
hrYqlA/4O/CG5LHKpgvP7NwXV2e2AZsqyXqKKGHuGDEixHmB1Grv7epUDZTrAyue
IA2BqcIa1BZmpfRVmjQi9dZDh6X6+cyiCUj2tIyM2KmrfYQpnoRK6NFvys6YoPrc
sZhIDXE/VE1rRWd5t57TEDwWGJ7TVPjdi7SNN4/43pW5dQdaEmxVeCLzgTj77ygL
O4GCCQTDhOHvlBFpxV3ln9SoQ0umkI+pWJujIdd8/l4Xe49hFsfp1R09+9tapk8+
NOYk3tP+9iizbaLLZVTeK6zcxlgSQUHBye6z8+ZNXbaDJGsA1Bdq5C5ALz9FQRhr
xyijRynUDrxX6fzpA8zFlfPMHIYV/ONMI4mTHkF/g+JMuGyx9QkK3CEHbH9tf/tV
FcRBWToAE41AJo9lnmNAFsGmw1wAW1tSqJnCJYRkZBRwpMsC8PrT3mKedLkUj3ZO
VuMtcm863XOUgyBImW6wIJvDzTzkDj7MrhpdvFNb37EwCTGhy+WkJEuF5u7KHW/X
R5+SPS48pK0fkADOo9LoU1785O9a8i2aNrFlybZtQZl4fXLupwNJttXD8x20AA0G
mTlDAOiNDfq1Hof2hZgWT+LzueeJ/yZnMBw0nqL+AlEI28DVOyO4XeI69684832K
LTT/lCISHgyZwFPtu0aOABZkYGbcuP5/YJsvODEPp2qK3VdedGr59+Nxo0a4BEjl
Y+sWRFCVxDeE5YhYUyBNXaI5JAWcmWZuc1+sf+gJEViSuD7UvRbc2kPanka3g9Wf
/83qyxXjLHReQGUUphDpXmiL+J5pJQkZc9XYc1+AgF/Vew82fVAuf8exOb/mzDa8
s/p0pLa/3u8053yLxOgnkhNZCHlgEO3N+zUFnt5yO7LK6GgtyLfxFTfUAQd44xUn
4HprkGbdFAOQOQeoEtCo77NpjUJSJdN6wHyNiScNrCTg2YcEXKw/BoG8E1+MiDvW
d1jSQfJlZ4jSAW6tEIrR9H2Xci00zwuLDbGS9njwQoMnFq5thOea1Kbg7Muto/lx
6GzkPIcyIcowWwm7WKxqEk4RsOZWd4xi4fDL9qEo32yfamk0QtzpXE5u3QFquO77
QhzO9nFco5kYhTvr1Udmx2UWkuI8CErB/ecLcdu39vy0mhudboZ8FdEF49zRqeI+
OQ+mCk29ofEYhWIBpodm6FWqr7eHT1X76gjN0nmZhCvJ6tc72hxb6bDiqkjgbA5E
Xgv8NxmGULcNHzvrDbZV5Ox7mooQ8muZw8nR+RWWvwyaMXvDVgzbpE+fh0kmhuMc
RB0RhTFha0zlULONgX/cH1pNLQcLw8sb+8LjRPT01klW7DgKmvBEiCWM/m40HvqA
DgGpmFo3Rs2YUWWnTni0MCqnSurvpS30awOugA27bh+VkWC9+er5n9iEN5oTU4iG
oDwZQXRmqJHneQ7i+icarh1WeBC/bRL4UZmjckxPiYCkLth8vuMsVYKeA+UXjyg7
CDO8QaxvTXOU0OrLv8HEo+biJqbO9enq15owC4kd0AmuPD/crSxNLJk3bX8tKttC
8YRF+t7xyihbpyS3P3aKpLFSEW26+otX+8t6ajK78mmBxDQBiRxTMbILQdxK5SjX
XUbf+fmFvmf7ke5NMXkobFvI313awwRQloqbkgA4FUPuDJ7C5F7FaFAHywdMFgIH
eRA86R7ioud4A9dvZHlASVIgR0xVr/WtbBwFMybIvd2rlDeewz4jp4zZwPsX/Lxm
ghhALV1N21eWVWFHhnz/5dqi2xnea7yCyLnV/S8LbAO3oEwMDtEjPnXx0tFAoUrk
fFseWXzUSBKAh40jY9zA7oug717i5VN4XjMHxfKfxbK8kRCcYpfSMcwULu8rrxJx
kHpgZSZxij0xQ8lkBAucpfhrvfaxdplnUtD3dZVN79PSXm35GpD1S/OQzj2E/rYI
`pragma protect end_protected
